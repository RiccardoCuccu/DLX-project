
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (OP_SLL, OP_SRL, OP_SRA, OP_ADD, OP_ADDU, OP_SUB, OP_SUBU, 
   OP_AND, OP_OR, OP_XOR, OP_SEQ, OP_SNE, OP_SLT, OP_SGT, OP_SLE, OP_SGE, 
   OP_MOVI2S, OP_MOVS2I, OP_MOVF, OP_MOVD, OP_MOVFP2I, OP_MOVI2FP, OP_MOVI2T, 
   OP_MOVT2I, OP_SLTU, OP_SGTU, OP_SLEU, OP_SGEU, OP_ADDF, OP_SUBF, OP_MULTF, 
   OP_DIVF, OP_ADDD, OP_SUBD, OP_MULTD, OP_DIVD, OP_CVTF2D, OP_CVTF2I, 
   OP_CVTD2F, OP_CVTD2I, OP_CVTI2F, OP_CVTI2D, OP_MULT, OP_DIV, OP_EQF, OP_NEF,
   OP_LTF, OP_GTF, OP_LEF, OP_GEF, OP_MULTU, OP_DIVU, OP_EQD, OP_NED, OP_LTD, 
   OP_GTD, OP_LED, OP_GED, OP_BEQZ, OP_BNEZ, OP_BFPT, OP_BFPF, OP_ADDI, 
   OP_ADDUI, OP_SUBI, OP_SUBUI, OP_ANDI, OP_ORI, OP_XORI, OP_LHI, OP_RFE, 
   OP_TRAP, OP_JR, OP_JALR, OP_SLLI, OP_SRLI, OP_SRAI, OP_SEQI, OP_SNEI, 
   OP_SLTI, OP_SGTI, OP_SLEI, OP_SGEI, OP_LB, OP_LH, OP_LW, OP_LBU, OP_LHU, 
   OP_LF, OP_LD, OP_SB, OP_SH, OP_SW, OP_SF, OP_SD, OP_ITLB, OP_SLTUI, 
   OP_SGTUI, OP_SLEUI, OP_SGEUI, OP_J, OP_JAL, OP_NOP);
attribute ENUM_ENCODING of aluOp : type is 
   "0000000 0000001 0000010 0000011 0000100 0000101 0000110 0000111 0001000 0001001 0001010 0001011 0001100 0001101 0001110 0001111 0010000 0010001 0010010 0010011 0010100 0010101 0010110 0010111 0011000 0011001 0011010 0011011 0011100 0011101 0011110 0011111 0100000 0100001 0100010 0100011 0100100 0100101 0100110 0100111 0101000 0101001 0101010 0101011 0101100 0101101 0101110 0101111 0110000 0110001 0110010 0110011 0110100 0110101 0110110 0110111 0111000 0111001 0111010 0111011 0111100 0111101 0111110 0111111 1000000 1000001 1000010 1000011 1000100 1000101 1000110 1000111 1001000 1001001 1001010 1001011 1001100 1001101 1001110 1001111 1010000 1010001 1010010 1010011 1010100 1010101 1010110 1010111 1011000 1011001 1011010 1011011 1011100 1011101 1011110 1011111 1100000 1100001 1100010 1100011 1100100 1100101 1100110";
   
   -- Declarations for conversion functions.
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when OP_SLL => return "0000000";
         when OP_SRL => return "0000001";
         when OP_SRA => return "0000010";
         when OP_ADD => return "0000011";
         when OP_ADDU => return "0000100";
         when OP_SUB => return "0000101";
         when OP_SUBU => return "0000110";
         when OP_AND => return "0000111";
         when OP_OR => return "0001000";
         when OP_XOR => return "0001001";
         when OP_SEQ => return "0001010";
         when OP_SNE => return "0001011";
         when OP_SLT => return "0001100";
         when OP_SGT => return "0001101";
         when OP_SLE => return "0001110";
         when OP_SGE => return "0001111";
         when OP_MOVI2S => return "0010000";
         when OP_MOVS2I => return "0010001";
         when OP_MOVF => return "0010010";
         when OP_MOVD => return "0010011";
         when OP_MOVFP2I => return "0010100";
         when OP_MOVI2FP => return "0010101";
         when OP_MOVI2T => return "0010110";
         when OP_MOVT2I => return "0010111";
         when OP_SLTU => return "0011000";
         when OP_SGTU => return "0011001";
         when OP_SLEU => return "0011010";
         when OP_SGEU => return "0011011";
         when OP_ADDF => return "0011100";
         when OP_SUBF => return "0011101";
         when OP_MULTF => return "0011110";
         when OP_DIVF => return "0011111";
         when OP_ADDD => return "0100000";
         when OP_SUBD => return "0100001";
         when OP_MULTD => return "0100010";
         when OP_DIVD => return "0100011";
         when OP_CVTF2D => return "0100100";
         when OP_CVTF2I => return "0100101";
         when OP_CVTD2F => return "0100110";
         when OP_CVTD2I => return "0100111";
         when OP_CVTI2F => return "0101000";
         when OP_CVTI2D => return "0101001";
         when OP_MULT => return "0101010";
         when OP_DIV => return "0101011";
         when OP_EQF => return "0101100";
         when OP_NEF => return "0101101";
         when OP_LTF => return "0101110";
         when OP_GTF => return "0101111";
         when OP_LEF => return "0110000";
         when OP_GEF => return "0110001";
         when OP_MULTU => return "0110010";
         when OP_DIVU => return "0110011";
         when OP_EQD => return "0110100";
         when OP_NED => return "0110101";
         when OP_LTD => return "0110110";
         when OP_GTD => return "0110111";
         when OP_LED => return "0111000";
         when OP_GED => return "0111001";
         when OP_BEQZ => return "0111010";
         when OP_BNEZ => return "0111011";
         when OP_BFPT => return "0111100";
         when OP_BFPF => return "0111101";
         when OP_ADDI => return "0111110";
         when OP_ADDUI => return "0111111";
         when OP_SUBI => return "1000000";
         when OP_SUBUI => return "1000001";
         when OP_ANDI => return "1000010";
         when OP_ORI => return "1000011";
         when OP_XORI => return "1000100";
         when OP_LHI => return "1000101";
         when OP_RFE => return "1000110";
         when OP_TRAP => return "1000111";
         when OP_JR => return "1001000";
         when OP_JALR => return "1001001";
         when OP_SLLI => return "1001010";
         when OP_SRLI => return "1001011";
         when OP_SRAI => return "1001100";
         when OP_SEQI => return "1001101";
         when OP_SNEI => return "1001110";
         when OP_SLTI => return "1001111";
         when OP_SGTI => return "1010000";
         when OP_SLEI => return "1010001";
         when OP_SGEI => return "1010010";
         when OP_LB => return "1010011";
         when OP_LH => return "1010100";
         when OP_LW => return "1010101";
         when OP_LBU => return "1010110";
         when OP_LHU => return "1010111";
         when OP_LF => return "1011000";
         when OP_LD => return "1011001";
         when OP_SB => return "1011010";
         when OP_SH => return "1011011";
         when OP_SW => return "1011100";
         when OP_SF => return "1011101";
         when OP_SD => return "1011110";
         when OP_ITLB => return "1011111";
         when OP_SLTUI => return "1100000";
         when OP_SGTUI => return "1100001";
         when OP_SLEUI => return "1100010";
         when OP_SGEUI => return "1100011";
         when OP_J => return "1100100";
         when OP_JAL => return "1100101";
         when OP_NOP => return "1100110";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

   port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  DOUT :
         out std_logic_vector (31 downto 0));

end DLX_IRAM_RAM_DEPTH256_I_SIZE32;

architecture SYN_BEHAVIORAL of DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_DRAM_N256_NW32 is

   port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector (31 
         downto 0);  DOUT : out std_logic_vector (31 downto 0));

end DLX_DRAM_N256_NW32;

architecture SYN_BEHAVIORAL of DLX_DRAM_N256_NW32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RF_N32_NA5 is

   port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
         ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_N32_NA5;

architecture SYN_BEHAVIORAL of RF_N32_NA5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REG_0_31_port, REG_0_30_port, REG_0_29_port, REG_0_28_port, 
      REG_0_27_port, REG_0_26_port, REG_0_25_port, REG_0_24_port, REG_0_23_port
      , REG_0_22_port, REG_0_21_port, REG_0_20_port, REG_0_19_port, 
      REG_0_18_port, REG_0_17_port, REG_0_16_port, REG_0_15_port, REG_0_14_port
      , REG_0_13_port, REG_0_12_port, REG_0_11_port, REG_0_10_port, 
      REG_0_9_port, REG_0_8_port, REG_0_7_port, REG_0_6_port, REG_0_5_port, 
      REG_0_4_port, REG_0_3_port, REG_0_2_port, REG_0_1_port, REG_0_0_port, 
      REG_31_31_port, REG_31_30_port, REG_31_29_port, REG_31_28_port, 
      REG_31_27_port, REG_31_26_port, REG_31_25_port, REG_31_24_port, 
      REG_31_23_port, REG_31_22_port, REG_31_21_port, REG_31_20_port, 
      REG_31_19_port, REG_31_18_port, REG_31_17_port, REG_31_16_port, 
      REG_31_15_port, REG_31_14_port, REG_31_13_port, REG_31_12_port, 
      REG_31_11_port, REG_31_10_port, REG_31_9_port, REG_31_8_port, 
      REG_31_7_port, REG_31_6_port, REG_31_5_port, REG_31_4_port, REG_31_3_port
      , REG_31_2_port, REG_31_1_port, REG_31_0_port, N156, N157, N158, N159, 
      N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, 
      N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, 
      N184, N185, N186, N187, N219, N220, N221, N222, N223, N224, N225, N226, 
      N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, 
      N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, 
      n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50 : 
      std_logic;

begin
   
   REG_reg_0_31_inst : DLH_X1 port map( G => n10, D => N250, Q => REG_0_31_port
                           );
   REG_reg_0_30_inst : DLH_X1 port map( G => n10, D => N249, Q => REG_0_30_port
                           );
   REG_reg_0_29_inst : DLH_X1 port map( G => n10, D => N248, Q => REG_0_29_port
                           );
   REG_reg_0_28_inst : DLH_X1 port map( G => n10, D => N247, Q => REG_0_28_port
                           );
   REG_reg_0_27_inst : DLH_X1 port map( G => n10, D => N246, Q => REG_0_27_port
                           );
   REG_reg_0_26_inst : DLH_X1 port map( G => n10, D => N245, Q => REG_0_26_port
                           );
   REG_reg_0_25_inst : DLH_X1 port map( G => n10, D => N244, Q => REG_0_25_port
                           );
   REG_reg_0_24_inst : DLH_X1 port map( G => n10, D => N243, Q => REG_0_24_port
                           );
   REG_reg_0_23_inst : DLH_X1 port map( G => n11, D => N242, Q => REG_0_23_port
                           );
   REG_reg_0_22_inst : DLH_X1 port map( G => n11, D => N241, Q => REG_0_22_port
                           );
   REG_reg_0_21_inst : DLH_X1 port map( G => n11, D => N240, Q => REG_0_21_port
                           );
   REG_reg_0_20_inst : DLH_X1 port map( G => n10, D => N239, Q => REG_0_20_port
                           );
   REG_reg_0_19_inst : DLH_X1 port map( G => n11, D => N238, Q => REG_0_19_port
                           );
   REG_reg_0_18_inst : DLH_X1 port map( G => n10, D => N237, Q => REG_0_18_port
                           );
   REG_reg_0_17_inst : DLH_X1 port map( G => n10, D => N236, Q => REG_0_17_port
                           );
   REG_reg_0_16_inst : DLH_X1 port map( G => n10, D => N235, Q => REG_0_16_port
                           );
   REG_reg_0_15_inst : DLH_X1 port map( G => n10, D => N234, Q => REG_0_15_port
                           );
   REG_reg_0_14_inst : DLH_X1 port map( G => n10, D => N233, Q => REG_0_14_port
                           );
   REG_reg_0_13_inst : DLH_X1 port map( G => n10, D => N232, Q => REG_0_13_port
                           );
   REG_reg_0_12_inst : DLH_X1 port map( G => n10, D => N231, Q => REG_0_12_port
                           );
   REG_reg_0_11_inst : DLH_X1 port map( G => n11, D => N230, Q => REG_0_11_port
                           );
   REG_reg_0_10_inst : DLH_X1 port map( G => n11, D => N229, Q => REG_0_10_port
                           );
   REG_reg_0_9_inst : DLH_X1 port map( G => n10, D => N228, Q => REG_0_9_port);
   REG_reg_0_8_inst : DLH_X1 port map( G => n10, D => N227, Q => REG_0_8_port);
   REG_reg_0_7_inst : DLH_X1 port map( G => n11, D => N226, Q => REG_0_7_port);
   REG_reg_0_6_inst : DLH_X1 port map( G => n11, D => N225, Q => REG_0_6_port);
   REG_reg_0_5_inst : DLH_X1 port map( G => n11, D => N224, Q => REG_0_5_port);
   REG_reg_0_4_inst : DLH_X1 port map( G => n11, D => N223, Q => REG_0_4_port);
   REG_reg_0_3_inst : DLH_X1 port map( G => n11, D => N222, Q => REG_0_3_port);
   REG_reg_0_2_inst : DLH_X1 port map( G => n11, D => N221, Q => REG_0_2_port);
   REG_reg_0_1_inst : DLH_X1 port map( G => n11, D => N220, Q => REG_0_1_port);
   REG_reg_0_0_inst : DLH_X1 port map( G => n11, D => N219, Q => REG_0_0_port);
   REG_reg_31_31_inst : DLH_X1 port map( G => n11, D => N187, Q => 
                           REG_31_31_port);
   REG_reg_31_30_inst : DLH_X1 port map( G => n11, D => N186, Q => 
                           REG_31_30_port);
   REG_reg_31_29_inst : DLH_X1 port map( G => n11, D => N185, Q => 
                           REG_31_29_port);
   REG_reg_31_28_inst : DLH_X1 port map( G => n11, D => N184, Q => 
                           REG_31_28_port);
   REG_reg_31_27_inst : DLH_X1 port map( G => n10, D => N183, Q => 
                           REG_31_27_port);
   REG_reg_31_26_inst : DLH_X1 port map( G => n10, D => N182, Q => 
                           REG_31_26_port);
   REG_reg_31_25_inst : DLH_X1 port map( G => n10, D => N181, Q => 
                           REG_31_25_port);
   REG_reg_31_24_inst : DLH_X1 port map( G => n11, D => N180, Q => 
                           REG_31_24_port);
   REG_reg_31_23_inst : DLH_X1 port map( G => n10, D => N179, Q => 
                           REG_31_23_port);
   REG_reg_31_22_inst : DLH_X1 port map( G => n10, D => N178, Q => 
                           REG_31_22_port);
   REG_reg_31_21_inst : DLH_X1 port map( G => n11, D => N177, Q => 
                           REG_31_21_port);
   REG_reg_31_20_inst : DLH_X1 port map( G => n10, D => N176, Q => 
                           REG_31_20_port);
   REG_reg_31_19_inst : DLH_X1 port map( G => n11, D => N175, Q => 
                           REG_31_19_port);
   REG_reg_31_18_inst : DLH_X1 port map( G => n10, D => N174, Q => 
                           REG_31_18_port);
   REG_reg_31_17_inst : DLH_X1 port map( G => n11, D => N173, Q => 
                           REG_31_17_port);
   REG_reg_31_16_inst : DLH_X1 port map( G => n11, D => N172, Q => 
                           REG_31_16_port);
   REG_reg_31_15_inst : DLH_X1 port map( G => n11, D => N171, Q => 
                           REG_31_15_port);
   REG_reg_31_14_inst : DLH_X1 port map( G => n11, D => N170, Q => 
                           REG_31_14_port);
   REG_reg_31_13_inst : DLH_X1 port map( G => n10, D => N169, Q => 
                           REG_31_13_port);
   REG_reg_31_12_inst : DLH_X1 port map( G => n11, D => N168, Q => 
                           REG_31_12_port);
   REG_reg_31_11_inst : DLH_X1 port map( G => n10, D => N167, Q => 
                           REG_31_11_port);
   REG_reg_31_10_inst : DLH_X1 port map( G => n11, D => N166, Q => 
                           REG_31_10_port);
   REG_reg_31_9_inst : DLH_X1 port map( G => n10, D => N165, Q => REG_31_9_port
                           );
   REG_reg_31_8_inst : DLH_X1 port map( G => n11, D => N164, Q => REG_31_8_port
                           );
   REG_reg_31_7_inst : DLH_X1 port map( G => n10, D => N163, Q => REG_31_7_port
                           );
   REG_reg_31_6_inst : DLH_X1 port map( G => n11, D => N162, Q => REG_31_6_port
                           );
   REG_reg_31_5_inst : DLH_X1 port map( G => n10, D => N161, Q => REG_31_5_port
                           );
   REG_reg_31_4_inst : DLH_X1 port map( G => n10, D => N160, Q => REG_31_4_port
                           );
   REG_reg_31_3_inst : DLH_X1 port map( G => n10, D => N159, Q => REG_31_3_port
                           );
   REG_reg_31_2_inst : DLH_X1 port map( G => n11, D => N158, Q => REG_31_2_port
                           );
   REG_reg_31_1_inst : DLH_X1 port map( G => n11, D => N157, Q => REG_31_1_port
                           );
   REG_reg_31_0_inst : DLH_X1 port map( G => n11, D => N156, Q => REG_31_0_port
                           );
   U3 : CLKBUF_X2 port map( A => n48, Z => n7);
   U4 : CLKBUF_X2 port map( A => n50, Z => n8);
   U5 : INV_X1 port map( A => RST, ZN => n11);
   U6 : INV_X1 port map( A => RST, ZN => n10);
   U7 : OR4_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), A3 => ADD_WR(0), A4 
                           => ADD_WR(2), ZN => n12);
   U8 : NOR2_X1 port map( A1 => ADD_WR(1), A2 => n12, ZN => n35);
   U9 : CLKBUF_X1 port map( A => n35, Z => n46);
   U10 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(0), ZN => n13);
   U11 : INV_X1 port map( A => n13, ZN => N156);
   U12 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(31), ZN => n45);
   U13 : INV_X1 port map( A => n45, ZN => N187);
   U14 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(30), ZN => n44);
   U15 : INV_X1 port map( A => n44, ZN => N186);
   U16 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(29), ZN => n43);
   U17 : INV_X1 port map( A => n43, ZN => N185);
   U18 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(28), ZN => n42);
   U19 : INV_X1 port map( A => n42, ZN => N184);
   U20 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(27), ZN => n41);
   U21 : INV_X1 port map( A => n41, ZN => N183);
   U22 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(26), ZN => n40);
   U23 : INV_X1 port map( A => n40, ZN => N182);
   U24 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(25), ZN => n39);
   U25 : INV_X1 port map( A => n39, ZN => N181);
   U26 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(24), ZN => n38);
   U27 : INV_X1 port map( A => n38, ZN => N180);
   U28 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(23), ZN => n37);
   U29 : INV_X1 port map( A => n37, ZN => N179);
   U30 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(22), ZN => n36);
   U31 : INV_X1 port map( A => n36, ZN => N178);
   U32 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(21), ZN => n34);
   U33 : INV_X1 port map( A => n34, ZN => N177);
   U34 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(20), ZN => n33);
   U35 : INV_X1 port map( A => n33, ZN => N176);
   U36 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(19), ZN => n32);
   U37 : INV_X1 port map( A => n32, ZN => N175);
   U38 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(18), ZN => n31);
   U39 : INV_X1 port map( A => n31, ZN => N174);
   U40 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(17), ZN => n30);
   U41 : INV_X1 port map( A => n30, ZN => N173);
   U42 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(16), ZN => n29);
   U43 : INV_X1 port map( A => n29, ZN => N172);
   U44 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(15), ZN => n28);
   U45 : INV_X1 port map( A => n28, ZN => N171);
   U46 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(14), ZN => n27);
   U47 : INV_X1 port map( A => n27, ZN => N170);
   U48 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(13), ZN => n26);
   U49 : INV_X1 port map( A => n26, ZN => N169);
   U50 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(12), ZN => n25);
   U51 : INV_X1 port map( A => n25, ZN => N168);
   U52 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(11), ZN => n24);
   U53 : INV_X1 port map( A => n24, ZN => N167);
   U54 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(10), ZN => n23);
   U55 : INV_X1 port map( A => n23, ZN => N166);
   U56 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(9), ZN => n22);
   U57 : INV_X1 port map( A => n22, ZN => N165);
   U58 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(8), ZN => n21);
   U59 : INV_X1 port map( A => n21, ZN => N164);
   U60 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(7), ZN => n20);
   U61 : INV_X1 port map( A => n20, ZN => N163);
   U62 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(6), ZN => n19);
   U63 : INV_X1 port map( A => n19, ZN => N162);
   U64 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(5), ZN => n18);
   U65 : INV_X1 port map( A => n18, ZN => N161);
   U66 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(4), ZN => n17);
   U67 : INV_X1 port map( A => n17, ZN => N160);
   U68 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(3), ZN => n16);
   U69 : INV_X1 port map( A => n16, ZN => N159);
   U70 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(2), ZN => n15);
   U71 : INV_X1 port map( A => n15, ZN => N158);
   U72 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(1), ZN => n14);
   U73 : INV_X1 port map( A => n14, ZN => N157);
   U74 : NOR2_X1 port map( A1 => n46, A2 => n13, ZN => N219);
   U75 : NOR2_X1 port map( A1 => n46, A2 => n14, ZN => N220);
   U76 : NOR2_X1 port map( A1 => n46, A2 => n15, ZN => N221);
   U77 : NOR2_X1 port map( A1 => n46, A2 => n16, ZN => N222);
   U78 : NOR2_X1 port map( A1 => n46, A2 => n17, ZN => N223);
   U79 : NOR2_X1 port map( A1 => n46, A2 => n18, ZN => N224);
   U80 : NOR2_X1 port map( A1 => n46, A2 => n19, ZN => N225);
   U81 : NOR2_X1 port map( A1 => n46, A2 => n20, ZN => N226);
   U82 : NOR2_X1 port map( A1 => n46, A2 => n21, ZN => N227);
   U83 : NOR2_X1 port map( A1 => n46, A2 => n22, ZN => N228);
   U84 : NOR2_X1 port map( A1 => n35, A2 => n23, ZN => N229);
   U85 : NOR2_X1 port map( A1 => n46, A2 => n24, ZN => N230);
   U86 : NOR2_X1 port map( A1 => n46, A2 => n25, ZN => N231);
   U87 : NOR2_X1 port map( A1 => n35, A2 => n26, ZN => N232);
   U88 : NOR2_X1 port map( A1 => n35, A2 => n27, ZN => N233);
   U89 : NOR2_X1 port map( A1 => n35, A2 => n28, ZN => N234);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n29, ZN => N235);
   U91 : NOR2_X1 port map( A1 => n35, A2 => n30, ZN => N236);
   U92 : NOR2_X1 port map( A1 => n35, A2 => n31, ZN => N237);
   U93 : NOR2_X1 port map( A1 => n35, A2 => n32, ZN => N238);
   U94 : NOR2_X1 port map( A1 => n35, A2 => n33, ZN => N239);
   U95 : NOR2_X1 port map( A1 => n35, A2 => n34, ZN => N240);
   U96 : NOR2_X1 port map( A1 => n46, A2 => n36, ZN => N241);
   U97 : NOR2_X1 port map( A1 => n46, A2 => n37, ZN => N242);
   U98 : NOR2_X1 port map( A1 => n46, A2 => n38, ZN => N243);
   U99 : NOR2_X1 port map( A1 => n46, A2 => n39, ZN => N244);
   U100 : NOR2_X1 port map( A1 => n46, A2 => n40, ZN => N245);
   U101 : NOR2_X1 port map( A1 => n46, A2 => n41, ZN => N246);
   U102 : NOR2_X1 port map( A1 => n46, A2 => n42, ZN => N247);
   U103 : NOR2_X1 port map( A1 => n46, A2 => n43, ZN => N248);
   U104 : NOR2_X1 port map( A1 => n46, A2 => n44, ZN => N249);
   U105 : NOR2_X1 port map( A1 => n46, A2 => n45, ZN => N250);
   U106 : OR4_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => ADD_RD2(2)
                           , A4 => ADD_RD2(4), ZN => n47);
   U107 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => n47, ZN => n48);
   U108 : MUX2_X1 port map( A => REG_31_31_port, B => REG_0_31_port, S => n7, Z
                           => OUT2(31));
   U109 : MUX2_X1 port map( A => REG_31_30_port, B => REG_0_30_port, S => n7, Z
                           => OUT2(30));
   U110 : MUX2_X1 port map( A => REG_31_29_port, B => REG_0_29_port, S => n7, Z
                           => OUT2(29));
   U111 : MUX2_X1 port map( A => REG_31_28_port, B => REG_0_28_port, S => n7, Z
                           => OUT2(28));
   U112 : MUX2_X1 port map( A => REG_31_27_port, B => REG_0_27_port, S => n7, Z
                           => OUT2(27));
   U113 : MUX2_X1 port map( A => REG_31_26_port, B => REG_0_26_port, S => n7, Z
                           => OUT2(26));
   U114 : MUX2_X1 port map( A => REG_31_25_port, B => REG_0_25_port, S => n7, Z
                           => OUT2(25));
   U115 : MUX2_X1 port map( A => REG_31_24_port, B => REG_0_24_port, S => n7, Z
                           => OUT2(24));
   U116 : MUX2_X1 port map( A => REG_31_23_port, B => REG_0_23_port, S => n7, Z
                           => OUT2(23));
   U117 : MUX2_X1 port map( A => REG_31_22_port, B => REG_0_22_port, S => n7, Z
                           => OUT2(22));
   U118 : MUX2_X1 port map( A => REG_31_21_port, B => REG_0_21_port, S => n7, Z
                           => OUT2(21));
   U119 : MUX2_X1 port map( A => REG_31_20_port, B => REG_0_20_port, S => n7, Z
                           => OUT2(20));
   U120 : MUX2_X1 port map( A => REG_31_19_port, B => REG_0_19_port, S => n7, Z
                           => OUT2(19));
   U121 : MUX2_X1 port map( A => REG_31_18_port, B => REG_0_18_port, S => n48, 
                           Z => OUT2(18));
   U122 : MUX2_X1 port map( A => REG_31_17_port, B => REG_0_17_port, S => n48, 
                           Z => OUT2(17));
   U123 : MUX2_X1 port map( A => REG_31_16_port, B => REG_0_16_port, S => n48, 
                           Z => OUT2(16));
   U124 : MUX2_X1 port map( A => REG_31_15_port, B => REG_0_15_port, S => n48, 
                           Z => OUT2(15));
   U125 : MUX2_X1 port map( A => REG_31_14_port, B => REG_0_14_port, S => n48, 
                           Z => OUT2(14));
   U126 : MUX2_X1 port map( A => REG_31_13_port, B => REG_0_13_port, S => n48, 
                           Z => OUT2(13));
   U127 : MUX2_X1 port map( A => REG_31_12_port, B => REG_0_12_port, S => n48, 
                           Z => OUT2(12));
   U128 : MUX2_X1 port map( A => REG_31_11_port, B => REG_0_11_port, S => n48, 
                           Z => OUT2(11));
   U129 : MUX2_X1 port map( A => REG_31_10_port, B => REG_0_10_port, S => n48, 
                           Z => OUT2(10));
   U130 : MUX2_X1 port map( A => REG_31_9_port, B => REG_0_9_port, S => n7, Z 
                           => OUT2(9));
   U131 : MUX2_X1 port map( A => REG_31_8_port, B => REG_0_8_port, S => n7, Z 
                           => OUT2(8));
   U132 : MUX2_X1 port map( A => REG_31_7_port, B => REG_0_7_port, S => n7, Z 
                           => OUT2(7));
   U133 : MUX2_X1 port map( A => REG_31_6_port, B => REG_0_6_port, S => n7, Z 
                           => OUT2(6));
   U134 : MUX2_X1 port map( A => REG_31_5_port, B => REG_0_5_port, S => n7, Z 
                           => OUT2(5));
   U135 : MUX2_X1 port map( A => REG_31_4_port, B => REG_0_4_port, S => n7, Z 
                           => OUT2(4));
   U136 : MUX2_X1 port map( A => REG_31_3_port, B => REG_0_3_port, S => n7, Z 
                           => OUT2(3));
   U137 : MUX2_X1 port map( A => REG_31_2_port, B => REG_0_2_port, S => n7, Z 
                           => OUT2(2));
   U138 : MUX2_X1 port map( A => REG_31_1_port, B => REG_0_1_port, S => n7, Z 
                           => OUT2(1));
   U139 : MUX2_X1 port map( A => REG_31_0_port, B => REG_0_0_port, S => n7, Z 
                           => OUT2(0));
   U140 : OR4_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => ADD_RD1(2)
                           , A4 => ADD_RD1(4), ZN => n49);
   U141 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => n49, ZN => n50);
   U142 : MUX2_X1 port map( A => REG_31_31_port, B => REG_0_31_port, S => n8, Z
                           => OUT1(31));
   U143 : MUX2_X1 port map( A => REG_31_30_port, B => REG_0_30_port, S => n8, Z
                           => OUT1(30));
   U144 : MUX2_X1 port map( A => REG_31_29_port, B => REG_0_29_port, S => n8, Z
                           => OUT1(29));
   U145 : MUX2_X1 port map( A => REG_31_28_port, B => REG_0_28_port, S => n8, Z
                           => OUT1(28));
   U146 : MUX2_X1 port map( A => REG_31_27_port, B => REG_0_27_port, S => n8, Z
                           => OUT1(27));
   U147 : MUX2_X1 port map( A => REG_31_26_port, B => REG_0_26_port, S => n8, Z
                           => OUT1(26));
   U148 : MUX2_X1 port map( A => REG_31_25_port, B => REG_0_25_port, S => n8, Z
                           => OUT1(25));
   U149 : MUX2_X1 port map( A => REG_31_24_port, B => REG_0_24_port, S => n8, Z
                           => OUT1(24));
   U150 : MUX2_X1 port map( A => REG_31_23_port, B => REG_0_23_port, S => n8, Z
                           => OUT1(23));
   U151 : MUX2_X1 port map( A => REG_31_22_port, B => REG_0_22_port, S => n8, Z
                           => OUT1(22));
   U152 : MUX2_X1 port map( A => REG_31_21_port, B => REG_0_21_port, S => n8, Z
                           => OUT1(21));
   U153 : MUX2_X1 port map( A => REG_31_20_port, B => REG_0_20_port, S => n8, Z
                           => OUT1(20));
   U154 : MUX2_X1 port map( A => REG_31_19_port, B => REG_0_19_port, S => n8, Z
                           => OUT1(19));
   U155 : MUX2_X1 port map( A => REG_31_18_port, B => REG_0_18_port, S => n50, 
                           Z => OUT1(18));
   U156 : MUX2_X1 port map( A => REG_31_17_port, B => REG_0_17_port, S => n50, 
                           Z => OUT1(17));
   U157 : MUX2_X1 port map( A => REG_31_16_port, B => REG_0_16_port, S => n50, 
                           Z => OUT1(16));
   U158 : MUX2_X1 port map( A => REG_31_15_port, B => REG_0_15_port, S => n50, 
                           Z => OUT1(15));
   U159 : MUX2_X1 port map( A => REG_31_14_port, B => REG_0_14_port, S => n50, 
                           Z => OUT1(14));
   U160 : MUX2_X1 port map( A => REG_31_13_port, B => REG_0_13_port, S => n50, 
                           Z => OUT1(13));
   U161 : MUX2_X1 port map( A => REG_31_12_port, B => REG_0_12_port, S => n50, 
                           Z => OUT1(12));
   U162 : MUX2_X1 port map( A => REG_31_11_port, B => REG_0_11_port, S => n50, 
                           Z => OUT1(11));
   U163 : MUX2_X1 port map( A => REG_31_10_port, B => REG_0_10_port, S => n50, 
                           Z => OUT1(10));
   U164 : MUX2_X1 port map( A => REG_31_9_port, B => REG_0_9_port, S => n8, Z 
                           => OUT1(9));
   U165 : MUX2_X1 port map( A => REG_31_8_port, B => REG_0_8_port, S => n8, Z 
                           => OUT1(8));
   U166 : MUX2_X1 port map( A => REG_31_7_port, B => REG_0_7_port, S => n8, Z 
                           => OUT1(7));
   U167 : MUX2_X1 port map( A => REG_31_6_port, B => REG_0_6_port, S => n8, Z 
                           => OUT1(6));
   U168 : MUX2_X1 port map( A => REG_31_5_port, B => REG_0_5_port, S => n8, Z 
                           => OUT1(5));
   U169 : MUX2_X1 port map( A => REG_31_4_port, B => REG_0_4_port, S => n8, Z 
                           => OUT1(4));
   U170 : MUX2_X1 port map( A => REG_31_3_port, B => REG_0_3_port, S => n8, Z 
                           => OUT1(3));
   U171 : MUX2_X1 port map( A => REG_31_2_port, B => REG_0_2_port, S => n8, Z 
                           => OUT1(2));
   U172 : MUX2_X1 port map( A => REG_31_1_port, B => REG_0_1_port, S => n8, Z 
                           => OUT1(1));
   U173 : MUX2_X1 port map( A => REG_31_0_port, B => REG_0_0_port, S => n8, Z 
                           => OUT1(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_NB8 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
         std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);  Z
         : out std_logic);

end ALU_N32_NB8;

architecture SYN_BEHAVIORAL of ALU_N32_NB8 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X2
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal N96, OP_A_31_port, OP_A_30_port, OP_A_29_port, OP_A_28_port, 
      OP_A_27_port, OP_A_26_port, OP_A_25_port, OP_A_24_port, OP_A_23_port, 
      OP_A_22_port, OP_A_21_port, OP_A_20_port, OP_A_19_port, OP_A_18_port, 
      OP_A_17_port, OP_A_16_port, OP_A_15_port, OP_A_14_port, OP_A_13_port, 
      OP_A_12_port, OP_A_11_port, OP_A_10_port, OP_A_9_port, OP_A_8_port, 
      OP_A_7_port, OP_A_6_port, OP_A_5_port, OP_A_4_port, OP_A_3_port, 
      OP_A_2_port, OP_A_1_port, OP_A_0_port, OP_B_31_port, OP_B_30_port, 
      OP_B_29_port, OP_B_28_port, OP_B_27_port, OP_B_26_port, OP_B_25_port, 
      OP_B_24_port, OP_B_23_port, OP_B_22_port, OP_B_21_port, OP_B_20_port, 
      OP_B_19_port, OP_B_18_port, OP_B_17_port, OP_B_16_port, OP_B_15_port, 
      OP_B_14_port, OP_B_13_port, OP_B_12_port, OP_B_11_port, OP_B_10_port, 
      OP_B_9_port, OP_B_8_port, OP_B_7_port, OP_B_6_port, OP_B_5_port, 
      OP_B_4_port, OP_B_3_port, OP_B_2_port, OP_B_1_port, OP_B_0_port, OP_Ci, 
      OP_LOGIC_1_port, OP_LOGIC_0_port, OP_SHIFT, OP_COMPARE_3_port, 
      OP_COMPARE_2_port, OP_COMPARE_1_port, OP_COMPARE_0_port, N246, N247, N248
      , N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
      N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, 
      N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, 
      N285, N286, N287, N288, N289, C431_DATA4_3, C431_DATA4_4, C431_DATA4_5, 
      C431_DATA4_6, C431_DATA4_7, C431_DATA4_8, C431_DATA4_9, C431_DATA4_10, 
      C431_DATA4_11, C431_DATA4_12, C431_DATA4_13, C431_DATA4_14, C431_DATA4_15
      , C431_DATA4_16, C431_DATA4_17, C430_DATA4_5, C430_DATA4_6, C430_DATA4_7,
      C430_DATA4_8, C430_DATA4_9, C430_DATA4_10, C430_DATA4_11, C430_DATA4_12, 
      C430_DATA4_13, C430_DATA4_14, C430_DATA4_15, C430_DATA4_16, C430_DATA4_17
      , C430_DATA4_18, C430_DATA4_19, C429_DATA4_7, C429_DATA4_8, C429_DATA4_9,
      C429_DATA4_10, C429_DATA4_11, C429_DATA4_12, C429_DATA4_13, C429_DATA4_14
      , C429_DATA4_15, C429_DATA4_16, C429_DATA4_17, C429_DATA4_18, 
      C429_DATA4_19, C429_DATA4_20, C429_DATA4_21, C428_DATA4_1, C428_DATA4_2, 
      C428_DATA4_3, C428_DATA4_4, C428_DATA4_5, C428_DATA4_6, C428_DATA4_7, 
      C428_DATA4_8, C428_DATA4_9, C428_DATA4_10, C428_DATA4_11, C428_DATA4_12, 
      C428_DATA4_13, C428_DATA4_14, C428_DATA4_15, C2_DATA1_2, C2_DATA1_4, 
      C2_DATA1_6, DP_OP_440J3_122_9847_n80, DP_OP_440J3_122_9847_n79, 
      DP_OP_440J3_122_9847_n78, DP_OP_440J3_122_9847_n77, 
      DP_OP_440J3_122_9847_n76, DP_OP_440J3_122_9847_n75, 
      DP_OP_440J3_122_9847_n74, DP_OP_440J3_122_9847_n73, 
      DP_OP_440J3_122_9847_n72, DP_OP_440J3_122_9847_n71, 
      DP_OP_440J3_122_9847_n70, DP_OP_440J3_122_9847_n69, 
      DP_OP_440J3_122_9847_n68, DP_OP_440J3_122_9847_n67, 
      DP_OP_440J3_122_9847_n66, DP_OP_440J3_122_9847_n35, 
      DP_OP_440J3_122_9847_n34, DP_OP_440J3_122_9847_n33, 
      DP_OP_440J3_122_9847_n32, DP_OP_440J3_122_9847_n31, 
      DP_OP_440J3_122_9847_n30, DP_OP_440J3_122_9847_n29, 
      DP_OP_440J3_122_9847_n28, DP_OP_440J3_122_9847_n27, 
      DP_OP_440J3_122_9847_n26, DP_OP_440J3_122_9847_n25, 
      DP_OP_440J3_122_9847_n24, DP_OP_440J3_122_9847_n23, 
      DP_OP_440J3_122_9847_n22, DP_OP_440J3_122_9847_n21, 
      DP_OP_440J3_122_9847_n20, DP_OP_446J3_125_4819_n87, 
      DP_OP_446J3_125_4819_n86, DP_OP_446J3_125_4819_n85, 
      DP_OP_446J3_125_4819_n84, DP_OP_446J3_125_4819_n83, 
      DP_OP_446J3_125_4819_n82, DP_OP_446J3_125_4819_n81, 
      DP_OP_446J3_125_4819_n80, DP_OP_446J3_125_4819_n79, 
      DP_OP_446J3_125_4819_n78, DP_OP_446J3_125_4819_n77, 
      DP_OP_446J3_125_4819_n76, DP_OP_446J3_125_4819_n75, 
      DP_OP_446J3_125_4819_n74, DP_OP_446J3_125_4819_n73, 
      DP_OP_446J3_125_4819_n72, DP_OP_446J3_125_4819_n27, 
      DP_OP_446J3_125_4819_n26, DP_OP_446J3_125_4819_n25, 
      DP_OP_446J3_125_4819_n24, DP_OP_446J3_125_4819_n23, 
      DP_OP_446J3_125_4819_n22, DP_OP_446J3_125_4819_n21, 
      DP_OP_446J3_125_4819_n20, DP_OP_446J3_125_4819_n19, 
      DP_OP_446J3_125_4819_n18, DP_OP_446J3_125_4819_n17, 
      DP_OP_446J3_125_4819_n16, DP_OP_446J3_125_4819_n15, 
      DP_OP_446J3_125_4819_n14, DP_OP_446J3_125_4819_n13, 
      DP_OP_446J3_125_4819_n12, DP_OP_451J3_128_3502_n85, 
      DP_OP_451J3_128_3502_n84, DP_OP_451J3_128_3502_n83, 
      DP_OP_451J3_128_3502_n82, DP_OP_451J3_128_3502_n81, 
      DP_OP_451J3_128_3502_n80, DP_OP_451J3_128_3502_n79, 
      DP_OP_451J3_128_3502_n78, DP_OP_451J3_128_3502_n77, 
      DP_OP_451J3_128_3502_n76, DP_OP_451J3_128_3502_n75, 
      DP_OP_451J3_128_3502_n74, DP_OP_451J3_128_3502_n73, 
      DP_OP_451J3_128_3502_n72, DP_OP_451J3_128_3502_n71, 
      DP_OP_451J3_128_3502_n70, DP_OP_451J3_128_3502_n30, 
      DP_OP_451J3_128_3502_n29, DP_OP_451J3_128_3502_n28, 
      DP_OP_451J3_128_3502_n27, DP_OP_451J3_128_3502_n26, 
      DP_OP_451J3_128_3502_n25, DP_OP_451J3_128_3502_n24, 
      DP_OP_451J3_128_3502_n23, DP_OP_451J3_128_3502_n22, 
      DP_OP_451J3_128_3502_n21, DP_OP_451J3_128_3502_n20, 
      DP_OP_451J3_128_3502_n19, DP_OP_451J3_128_3502_n18, 
      DP_OP_451J3_128_3502_n17, DP_OP_451J3_128_3502_n16, 
      DP_OP_451J3_128_3502_n15, DP_OP_456J3_131_2158_n82, 
      DP_OP_456J3_131_2158_n81, DP_OP_456J3_131_2158_n80, 
      DP_OP_456J3_131_2158_n79, DP_OP_456J3_131_2158_n78, 
      DP_OP_456J3_131_2158_n77, DP_OP_456J3_131_2158_n76, 
      DP_OP_456J3_131_2158_n75, DP_OP_456J3_131_2158_n74, 
      DP_OP_456J3_131_2158_n73, DP_OP_456J3_131_2158_n72, 
      DP_OP_456J3_131_2158_n71, DP_OP_456J3_131_2158_n70, 
      DP_OP_456J3_131_2158_n69, DP_OP_456J3_131_2158_n68, 
      DP_OP_456J3_131_2158_n67, DP_OP_456J3_131_2158_n32, 
      DP_OP_456J3_131_2158_n31, DP_OP_456J3_131_2158_n30, 
      DP_OP_456J3_131_2158_n29, DP_OP_456J3_131_2158_n28, 
      DP_OP_456J3_131_2158_n27, DP_OP_456J3_131_2158_n26, 
      DP_OP_456J3_131_2158_n25, DP_OP_456J3_131_2158_n24, 
      DP_OP_456J3_131_2158_n23, DP_OP_456J3_131_2158_n22, 
      DP_OP_456J3_131_2158_n21, DP_OP_456J3_131_2158_n20, 
      DP_OP_456J3_131_2158_n19, DP_OP_456J3_131_2158_n18, 
      DP_OP_456J3_131_2158_n17, intadd_0_A_16_port, intadd_0_A_12_port, 
      intadd_0_A_11_port, intadd_0_A_10_port, intadd_0_A_9_port, 
      intadd_0_A_8_port, intadd_0_A_7_port, intadd_0_A_6_port, 
      intadd_0_A_5_port, intadd_0_A_4_port, intadd_0_A_3_port, 
      intadd_0_A_2_port, intadd_0_A_1_port, intadd_0_A_0_port, 
      intadd_0_B_14_port, intadd_0_B_13_port, intadd_0_B_12_port, 
      intadd_0_B_11_port, intadd_0_B_10_port, intadd_0_B_9_port, 
      intadd_0_B_8_port, intadd_0_B_7_port, intadd_0_B_6_port, 
      intadd_0_B_5_port, intadd_0_B_4_port, intadd_0_B_3_port, 
      intadd_0_B_2_port, intadd_0_B_1_port, intadd_0_B_0_port, intadd_0_CI, 
      intadd_0_SUM_26_port, intadd_0_SUM_25_port, intadd_0_SUM_24_port, 
      intadd_0_SUM_23_port, intadd_0_SUM_22_port, intadd_0_SUM_21_port, 
      intadd_0_SUM_20_port, intadd_0_SUM_19_port, intadd_0_SUM_18_port, 
      intadd_0_SUM_17_port, intadd_0_SUM_16_port, intadd_0_SUM_15_port, 
      intadd_0_SUM_14_port, intadd_0_SUM_13_port, intadd_0_SUM_12_port, 
      intadd_0_SUM_11_port, intadd_0_SUM_10_port, intadd_0_SUM_9_port, 
      intadd_0_SUM_8_port, intadd_0_SUM_7_port, intadd_0_SUM_6_port, 
      intadd_0_SUM_5_port, intadd_0_SUM_4_port, intadd_0_SUM_3_port, 
      intadd_0_SUM_2_port, intadd_0_SUM_1_port, intadd_0_SUM_0_port, 
      intadd_0_n27, intadd_0_n26, intadd_0_n25, intadd_0_n24, intadd_0_n23, 
      intadd_0_n22, intadd_0_n21, intadd_0_n20, intadd_0_n19, intadd_0_n18, 
      intadd_0_n17, intadd_0_n16, intadd_0_n15, intadd_0_n14, intadd_0_n13, 
      intadd_0_n12, intadd_0_n11, intadd_0_n10, intadd_0_n9, intadd_0_n8, 
      intadd_0_n7, intadd_0_n6, intadd_0_n5, intadd_0_n4, intadd_0_n3, 
      intadd_0_n2, intadd_0_n1, intadd_1_A_0_port, intadd_1_B_18_port, 
      intadd_1_B_14_port, intadd_1_B_13_port, intadd_1_B_12_port, 
      intadd_1_B_11_port, intadd_1_B_10_port, intadd_1_B_9_port, 
      intadd_1_B_8_port, intadd_1_B_7_port, intadd_1_B_6_port, 
      intadd_1_B_5_port, intadd_1_B_4_port, intadd_1_B_3_port, 
      intadd_1_B_2_port, intadd_1_B_1_port, intadd_1_B_0_port, 
      intadd_1_SUM_24_port, intadd_1_SUM_23_port, intadd_1_SUM_22_port, 
      intadd_1_SUM_21_port, intadd_1_SUM_20_port, intadd_1_SUM_19_port, 
      intadd_1_SUM_18_port, intadd_1_SUM_17_port, intadd_1_SUM_16_port, 
      intadd_1_SUM_15_port, intadd_1_SUM_14_port, intadd_1_SUM_13_port, 
      intadd_1_SUM_12_port, intadd_1_SUM_11_port, intadd_1_SUM_10_port, 
      intadd_1_SUM_9_port, intadd_1_SUM_8_port, intadd_1_SUM_7_port, 
      intadd_1_SUM_6_port, intadd_1_SUM_5_port, intadd_1_SUM_4_port, 
      intadd_1_SUM_3_port, intadd_1_SUM_2_port, intadd_1_SUM_1_port, 
      intadd_1_SUM_0_port, intadd_1_n25, intadd_1_n24, intadd_1_n23, 
      intadd_1_n22, intadd_1_n21, intadd_1_n20, intadd_1_n19, intadd_1_n18, 
      intadd_1_n17, intadd_1_n16, intadd_1_n15, intadd_1_n14, intadd_1_n13, 
      intadd_1_n12, intadd_1_n11, intadd_1_n10, intadd_1_n9, intadd_1_n8, 
      intadd_1_n7, intadd_1_n6, intadd_1_n5, intadd_1_n4, intadd_1_n3, 
      intadd_1_n2, intadd_1_n1, intadd_2_A_9_port, intadd_2_A_8_port, 
      intadd_2_A_7_port, intadd_2_A_6_port, intadd_2_A_5_port, 
      intadd_2_A_4_port, intadd_2_A_3_port, intadd_2_A_2_port, 
      intadd_2_A_1_port, intadd_2_A_0_port, intadd_2_B_0_port, 
      intadd_2_SUM_9_port, intadd_2_SUM_8_port, intadd_2_SUM_7_port, 
      intadd_2_SUM_6_port, intadd_2_SUM_5_port, intadd_2_SUM_4_port, 
      intadd_2_SUM_3_port, intadd_2_SUM_2_port, intadd_2_SUM_1_port, 
      intadd_2_SUM_0_port, intadd_2_n10, intadd_2_n9, intadd_2_n8, intadd_2_n7,
      intadd_2_n6, intadd_2_n5, intadd_2_n4, intadd_2_n3, intadd_2_n2, 
      intadd_2_n1, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
      n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96_port, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246_port, n247_port, n248_port, 
      n249_port, n250_port, n251_port, n252_port, n253_port, n254_port, 
      n255_port, n256_port, n257_port, n258_port, n259_port, n260_port, 
      n261_port, n262_port, n263_port, n264_port, n265_port, n266_port, 
      n267_port, n268_port, n269_port, n270_port, n271_port, n272_port, 
      n273_port, n274_port, n275_port, n276_port, n277_port, n278_port, 
      n279_port, n280_port, n281_port, n282_port, n283_port, n284_port, 
      n285_port, n286_port, n287_port, n288_port, n289_port, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
      n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, 
      n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
      n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
      n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
      n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, 
      n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
      n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
      n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n1415, n_1170 : std_logic;

begin
   
   OP_COMPARE_reg_3_inst : DLH_X1 port map( G => N285, D => N289, Q => 
                           OP_COMPARE_3_port);
   OP_COMPARE_reg_2_inst : DLH_X1 port map( G => N285, D => N288, Q => 
                           OP_COMPARE_2_port);
   OP_COMPARE_reg_1_inst : DLH_X1 port map( G => N285, D => N287, Q => 
                           OP_COMPARE_1_port);
   OP_COMPARE_reg_0_inst : DLH_X1 port map( G => N285, D => N286, Q => 
                           OP_COMPARE_0_port);
   OP_A_reg_31_inst : DLH_X1 port map( G => n1412, D => OP1(31), Q => 
                           OP_A_31_port);
   OP_A_reg_30_inst : DLH_X1 port map( G => n1412, D => OP1(30), Q => 
                           OP_A_30_port);
   OP_A_reg_29_inst : DLH_X1 port map( G => n1412, D => OP1(29), Q => 
                           OP_A_29_port);
   OP_A_reg_28_inst : DLH_X1 port map( G => n1412, D => OP1(28), Q => 
                           OP_A_28_port);
   OP_A_reg_27_inst : DLH_X1 port map( G => N246, D => OP1(27), Q => 
                           OP_A_27_port);
   OP_A_reg_26_inst : DLH_X1 port map( G => N246, D => OP1(26), Q => 
                           OP_A_26_port);
   OP_A_reg_25_inst : DLH_X1 port map( G => N246, D => OP1(25), Q => 
                           OP_A_25_port);
   OP_A_reg_24_inst : DLH_X1 port map( G => n1412, D => OP1(24), Q => 
                           OP_A_24_port);
   OP_A_reg_23_inst : DLH_X1 port map( G => N246, D => OP1(23), Q => 
                           OP_A_23_port);
   OP_A_reg_22_inst : DLH_X1 port map( G => n1412, D => OP1(22), Q => 
                           OP_A_22_port);
   OP_A_reg_21_inst : DLH_X1 port map( G => n1412, D => OP1(21), Q => 
                           OP_A_21_port);
   OP_A_reg_20_inst : DLH_X1 port map( G => N246, D => OP1(20), Q => 
                           OP_A_20_port);
   OP_A_reg_19_inst : DLH_X1 port map( G => N246, D => OP1(19), Q => 
                           OP_A_19_port);
   OP_A_reg_18_inst : DLH_X1 port map( G => n1412, D => OP1(18), Q => 
                           OP_A_18_port);
   OP_A_reg_17_inst : DLH_X1 port map( G => n1412, D => OP1(17), Q => 
                           OP_A_17_port);
   OP_A_reg_16_inst : DLH_X1 port map( G => n1412, D => OP1(16), Q => 
                           OP_A_16_port);
   OP_B_reg_31_inst : DLH_X1 port map( G => N246, D => N278, Q => OP_B_31_port)
                           ;
   OP_B_reg_30_inst : DLH_X1 port map( G => n1412, D => N277, Q => OP_B_30_port
                           );
   OP_B_reg_29_inst : DLH_X1 port map( G => N246, D => N276, Q => OP_B_29_port)
                           ;
   OP_B_reg_28_inst : DLH_X1 port map( G => N246, D => N275, Q => OP_B_28_port)
                           ;
   OP_B_reg_27_inst : DLH_X1 port map( G => N246, D => N274, Q => OP_B_27_port)
                           ;
   OP_B_reg_26_inst : DLH_X1 port map( G => N246, D => N273, Q => OP_B_26_port)
                           ;
   OP_B_reg_25_inst : DLH_X1 port map( G => N246, D => N272, Q => OP_B_25_port)
                           ;
   OP_B_reg_24_inst : DLH_X1 port map( G => N246, D => N271, Q => OP_B_24_port)
                           ;
   OP_B_reg_23_inst : DLH_X1 port map( G => N246, D => N270, Q => OP_B_23_port)
                           ;
   OP_B_reg_22_inst : DLH_X1 port map( G => N246, D => N269, Q => OP_B_22_port)
                           ;
   OP_B_reg_21_inst : DLH_X1 port map( G => N246, D => N268, Q => OP_B_21_port)
                           ;
   OP_B_reg_20_inst : DLH_X1 port map( G => N246, D => N267, Q => OP_B_20_port)
                           ;
   OP_B_reg_19_inst : DLH_X1 port map( G => n1412, D => N266, Q => OP_B_19_port
                           );
   OP_B_reg_18_inst : DLH_X1 port map( G => n1412, D => N265, Q => OP_B_18_port
                           );
   OP_B_reg_17_inst : DLH_X1 port map( G => n1412, D => N264, Q => OP_B_17_port
                           );
   OP_B_reg_16_inst : DLH_X1 port map( G => n1412, D => N263, Q => OP_B_16_port
                           );
   OP_B_reg_15_inst : DLH_X1 port map( G => n1412, D => N262, Q => OP_B_15_port
                           );
   OP_B_reg_14_inst : DLH_X1 port map( G => n1412, D => N261, Q => OP_B_14_port
                           );
   OP_B_reg_13_inst : DLH_X1 port map( G => n1412, D => N260, Q => OP_B_13_port
                           );
   OP_B_reg_12_inst : DLH_X1 port map( G => n1412, D => N259, Q => OP_B_12_port
                           );
   OP_B_reg_11_inst : DLH_X1 port map( G => n1412, D => N258, Q => OP_B_11_port
                           );
   OP_B_reg_10_inst : DLH_X1 port map( G => n1412, D => N257, Q => OP_B_10_port
                           );
   OP_B_reg_9_inst : DLH_X1 port map( G => N246, D => N256, Q => OP_B_9_port);
   OP_B_reg_8_inst : DLH_X1 port map( G => N246, D => N255, Q => OP_B_8_port);
   OP_B_reg_7_inst : DLH_X1 port map( G => N246, D => N254, Q => OP_B_7_port);
   OP_B_reg_6_inst : DLH_X1 port map( G => N246, D => N253, Q => OP_B_6_port);
   OP_B_reg_0_inst : DLH_X1 port map( G => n1412, D => N247, Q => OP_B_0_port);
   OP_Ci_reg : DLH_X1 port map( G => N279, D => N280, Q => OP_Ci);
   OP_LOGIC_reg_1_inst : DLH_X1 port map( G => N281, D => N283, Q => 
                           OP_LOGIC_1_port);
   OP_LOGIC_reg_0_inst : DLH_X1 port map( G => N281, D => N282, Q => 
                           OP_LOGIC_0_port);
   OP_SHIFT_reg : DLH_X1 port map( G => N284, D => N96, Q => OP_SHIFT);
   DP_OP_440J3_122_9847_U43 : HA_X1 port map( A => DP_OP_440J3_122_9847_n35, B 
                           => DP_OP_440J3_122_9847_n66, CO => 
                           DP_OP_440J3_122_9847_n34, S => C428_DATA4_1);
   DP_OP_440J3_122_9847_U42 : HA_X1 port map( A => DP_OP_440J3_122_9847_n34, B 
                           => DP_OP_440J3_122_9847_n67, CO => 
                           DP_OP_440J3_122_9847_n33, S => C428_DATA4_2);
   DP_OP_440J3_122_9847_U41 : HA_X1 port map( A => DP_OP_440J3_122_9847_n33, B 
                           => DP_OP_440J3_122_9847_n68, CO => 
                           DP_OP_440J3_122_9847_n32, S => C428_DATA4_3);
   DP_OP_440J3_122_9847_U40 : HA_X1 port map( A => DP_OP_440J3_122_9847_n32, B 
                           => DP_OP_440J3_122_9847_n69, CO => 
                           DP_OP_440J3_122_9847_n31, S => C428_DATA4_4);
   DP_OP_440J3_122_9847_U39 : HA_X1 port map( A => DP_OP_440J3_122_9847_n31, B 
                           => DP_OP_440J3_122_9847_n70, CO => 
                           DP_OP_440J3_122_9847_n30, S => C428_DATA4_5);
   DP_OP_440J3_122_9847_U38 : HA_X1 port map( A => DP_OP_440J3_122_9847_n30, B 
                           => DP_OP_440J3_122_9847_n71, CO => 
                           DP_OP_440J3_122_9847_n29, S => C428_DATA4_6);
   DP_OP_440J3_122_9847_U37 : HA_X1 port map( A => DP_OP_440J3_122_9847_n29, B 
                           => DP_OP_440J3_122_9847_n72, CO => 
                           DP_OP_440J3_122_9847_n28, S => C428_DATA4_7);
   DP_OP_440J3_122_9847_U36 : HA_X1 port map( A => DP_OP_440J3_122_9847_n28, B 
                           => DP_OP_440J3_122_9847_n73, CO => 
                           DP_OP_440J3_122_9847_n27, S => C428_DATA4_8);
   DP_OP_440J3_122_9847_U35 : HA_X1 port map( A => DP_OP_440J3_122_9847_n27, B 
                           => DP_OP_440J3_122_9847_n74, CO => 
                           DP_OP_440J3_122_9847_n26, S => C428_DATA4_9);
   DP_OP_440J3_122_9847_U34 : HA_X1 port map( A => DP_OP_440J3_122_9847_n26, B 
                           => DP_OP_440J3_122_9847_n75, CO => 
                           DP_OP_440J3_122_9847_n25, S => C428_DATA4_10);
   DP_OP_440J3_122_9847_U33 : HA_X1 port map( A => DP_OP_440J3_122_9847_n25, B 
                           => DP_OP_440J3_122_9847_n76, CO => 
                           DP_OP_440J3_122_9847_n24, S => C428_DATA4_11);
   DP_OP_440J3_122_9847_U32 : HA_X1 port map( A => DP_OP_440J3_122_9847_n24, B 
                           => DP_OP_440J3_122_9847_n77, CO => 
                           DP_OP_440J3_122_9847_n23, S => C428_DATA4_12);
   DP_OP_440J3_122_9847_U31 : HA_X1 port map( A => DP_OP_440J3_122_9847_n23, B 
                           => DP_OP_440J3_122_9847_n78, CO => 
                           DP_OP_440J3_122_9847_n22, S => C428_DATA4_13);
   DP_OP_440J3_122_9847_U30 : HA_X1 port map( A => DP_OP_440J3_122_9847_n22, B 
                           => DP_OP_440J3_122_9847_n79, CO => 
                           DP_OP_440J3_122_9847_n21, S => C428_DATA4_14);
   DP_OP_440J3_122_9847_U29 : HA_X1 port map( A => DP_OP_440J3_122_9847_n21, B 
                           => DP_OP_440J3_122_9847_n80, CO => 
                           DP_OP_440J3_122_9847_n20, S => C428_DATA4_15);
   DP_OP_446J3_125_4819_U33 : HA_X1 port map( A => n1414, B => 
                           DP_OP_446J3_125_4819_n72, CO => 
                           DP_OP_446J3_125_4819_n27, S => C2_DATA1_6);
   DP_OP_446J3_125_4819_U32 : HA_X1 port map( A => DP_OP_446J3_125_4819_n27, B 
                           => DP_OP_446J3_125_4819_n73, CO => 
                           DP_OP_446J3_125_4819_n26, S => C429_DATA4_7);
   DP_OP_446J3_125_4819_U31 : HA_X1 port map( A => DP_OP_446J3_125_4819_n26, B 
                           => DP_OP_446J3_125_4819_n74, CO => 
                           DP_OP_446J3_125_4819_n25, S => C429_DATA4_8);
   DP_OP_446J3_125_4819_U30 : HA_X1 port map( A => DP_OP_446J3_125_4819_n25, B 
                           => DP_OP_446J3_125_4819_n75, CO => 
                           DP_OP_446J3_125_4819_n24, S => C429_DATA4_9);
   DP_OP_446J3_125_4819_U29 : HA_X1 port map( A => DP_OP_446J3_125_4819_n24, B 
                           => DP_OP_446J3_125_4819_n76, CO => 
                           DP_OP_446J3_125_4819_n23, S => C429_DATA4_10);
   DP_OP_446J3_125_4819_U28 : HA_X1 port map( A => DP_OP_446J3_125_4819_n23, B 
                           => DP_OP_446J3_125_4819_n77, CO => 
                           DP_OP_446J3_125_4819_n22, S => C429_DATA4_11);
   DP_OP_446J3_125_4819_U27 : HA_X1 port map( A => DP_OP_446J3_125_4819_n22, B 
                           => DP_OP_446J3_125_4819_n78, CO => 
                           DP_OP_446J3_125_4819_n21, S => C429_DATA4_12);
   DP_OP_446J3_125_4819_U26 : HA_X1 port map( A => DP_OP_446J3_125_4819_n21, B 
                           => DP_OP_446J3_125_4819_n79, CO => 
                           DP_OP_446J3_125_4819_n20, S => C429_DATA4_13);
   DP_OP_446J3_125_4819_U25 : HA_X1 port map( A => DP_OP_446J3_125_4819_n20, B 
                           => DP_OP_446J3_125_4819_n80, CO => 
                           DP_OP_446J3_125_4819_n19, S => C429_DATA4_14);
   DP_OP_446J3_125_4819_U24 : HA_X1 port map( A => DP_OP_446J3_125_4819_n19, B 
                           => DP_OP_446J3_125_4819_n81, CO => 
                           DP_OP_446J3_125_4819_n18, S => C429_DATA4_15);
   DP_OP_446J3_125_4819_U23 : HA_X1 port map( A => DP_OP_446J3_125_4819_n18, B 
                           => DP_OP_446J3_125_4819_n82, CO => 
                           DP_OP_446J3_125_4819_n17, S => C429_DATA4_16);
   DP_OP_446J3_125_4819_U22 : HA_X1 port map( A => DP_OP_446J3_125_4819_n17, B 
                           => DP_OP_446J3_125_4819_n83, CO => 
                           DP_OP_446J3_125_4819_n16, S => C429_DATA4_17);
   DP_OP_446J3_125_4819_U21 : HA_X1 port map( A => DP_OP_446J3_125_4819_n16, B 
                           => DP_OP_446J3_125_4819_n84, CO => 
                           DP_OP_446J3_125_4819_n15, S => C429_DATA4_18);
   DP_OP_446J3_125_4819_U20 : HA_X1 port map( A => DP_OP_446J3_125_4819_n15, B 
                           => DP_OP_446J3_125_4819_n85, CO => 
                           DP_OP_446J3_125_4819_n14, S => C429_DATA4_19);
   DP_OP_446J3_125_4819_U19 : HA_X1 port map( A => DP_OP_446J3_125_4819_n14, B 
                           => DP_OP_446J3_125_4819_n86, CO => 
                           DP_OP_446J3_125_4819_n13, S => C429_DATA4_20);
   DP_OP_446J3_125_4819_U18 : HA_X1 port map( A => DP_OP_446J3_125_4819_n13, B 
                           => DP_OP_446J3_125_4819_n87, CO => 
                           DP_OP_446J3_125_4819_n12, S => C429_DATA4_21);
   DP_OP_451J3_128_3502_U37 : HA_X1 port map( A => n1413, B => 
                           DP_OP_451J3_128_3502_n70, CO => 
                           DP_OP_451J3_128_3502_n30, S => C2_DATA1_4);
   DP_OP_451J3_128_3502_U36 : HA_X1 port map( A => DP_OP_451J3_128_3502_n30, B 
                           => DP_OP_451J3_128_3502_n71, CO => 
                           DP_OP_451J3_128_3502_n29, S => C430_DATA4_5);
   DP_OP_451J3_128_3502_U35 : HA_X1 port map( A => DP_OP_451J3_128_3502_n29, B 
                           => DP_OP_451J3_128_3502_n72, CO => 
                           DP_OP_451J3_128_3502_n28, S => C430_DATA4_6);
   DP_OP_451J3_128_3502_U34 : HA_X1 port map( A => DP_OP_451J3_128_3502_n28, B 
                           => DP_OP_451J3_128_3502_n73, CO => 
                           DP_OP_451J3_128_3502_n27, S => C430_DATA4_7);
   DP_OP_451J3_128_3502_U33 : HA_X1 port map( A => DP_OP_451J3_128_3502_n27, B 
                           => DP_OP_451J3_128_3502_n74, CO => 
                           DP_OP_451J3_128_3502_n26, S => C430_DATA4_8);
   DP_OP_451J3_128_3502_U32 : HA_X1 port map( A => DP_OP_451J3_128_3502_n26, B 
                           => DP_OP_451J3_128_3502_n75, CO => 
                           DP_OP_451J3_128_3502_n25, S => C430_DATA4_9);
   DP_OP_451J3_128_3502_U31 : HA_X1 port map( A => DP_OP_451J3_128_3502_n25, B 
                           => DP_OP_451J3_128_3502_n76, CO => 
                           DP_OP_451J3_128_3502_n24, S => C430_DATA4_10);
   DP_OP_451J3_128_3502_U30 : HA_X1 port map( A => DP_OP_451J3_128_3502_n24, B 
                           => DP_OP_451J3_128_3502_n77, CO => 
                           DP_OP_451J3_128_3502_n23, S => C430_DATA4_11);
   DP_OP_451J3_128_3502_U29 : HA_X1 port map( A => DP_OP_451J3_128_3502_n23, B 
                           => DP_OP_451J3_128_3502_n78, CO => 
                           DP_OP_451J3_128_3502_n22, S => C430_DATA4_12);
   DP_OP_451J3_128_3502_U28 : HA_X1 port map( A => DP_OP_451J3_128_3502_n22, B 
                           => DP_OP_451J3_128_3502_n79, CO => 
                           DP_OP_451J3_128_3502_n21, S => C430_DATA4_13);
   DP_OP_451J3_128_3502_U27 : HA_X1 port map( A => DP_OP_451J3_128_3502_n21, B 
                           => DP_OP_451J3_128_3502_n80, CO => 
                           DP_OP_451J3_128_3502_n20, S => C430_DATA4_14);
   DP_OP_451J3_128_3502_U26 : HA_X1 port map( A => DP_OP_451J3_128_3502_n20, B 
                           => DP_OP_451J3_128_3502_n81, CO => 
                           DP_OP_451J3_128_3502_n19, S => C430_DATA4_15);
   DP_OP_451J3_128_3502_U25 : HA_X1 port map( A => DP_OP_451J3_128_3502_n19, B 
                           => DP_OP_451J3_128_3502_n82, CO => 
                           DP_OP_451J3_128_3502_n18, S => C430_DATA4_16);
   DP_OP_451J3_128_3502_U24 : HA_X1 port map( A => DP_OP_451J3_128_3502_n18, B 
                           => DP_OP_451J3_128_3502_n83, CO => 
                           DP_OP_451J3_128_3502_n17, S => C430_DATA4_17);
   DP_OP_451J3_128_3502_U23 : HA_X1 port map( A => DP_OP_451J3_128_3502_n17, B 
                           => DP_OP_451J3_128_3502_n84, CO => 
                           DP_OP_451J3_128_3502_n16, S => C430_DATA4_18);
   DP_OP_451J3_128_3502_U22 : HA_X1 port map( A => DP_OP_451J3_128_3502_n16, B 
                           => DP_OP_451J3_128_3502_n85, CO => 
                           DP_OP_451J3_128_3502_n15, S => C430_DATA4_19);
   DP_OP_456J3_131_2158_U40 : HA_X1 port map( A => n1415, B => 
                           DP_OP_456J3_131_2158_n67, CO => 
                           DP_OP_456J3_131_2158_n32, S => C2_DATA1_2);
   DP_OP_456J3_131_2158_U39 : HA_X1 port map( A => DP_OP_456J3_131_2158_n32, B 
                           => DP_OP_456J3_131_2158_n68, CO => 
                           DP_OP_456J3_131_2158_n31, S => C431_DATA4_3);
   DP_OP_456J3_131_2158_U38 : HA_X1 port map( A => DP_OP_456J3_131_2158_n31, B 
                           => DP_OP_456J3_131_2158_n69, CO => 
                           DP_OP_456J3_131_2158_n30, S => C431_DATA4_4);
   DP_OP_456J3_131_2158_U37 : HA_X1 port map( A => DP_OP_456J3_131_2158_n30, B 
                           => DP_OP_456J3_131_2158_n70, CO => 
                           DP_OP_456J3_131_2158_n29, S => C431_DATA4_5);
   DP_OP_456J3_131_2158_U36 : HA_X1 port map( A => DP_OP_456J3_131_2158_n29, B 
                           => DP_OP_456J3_131_2158_n71, CO => 
                           DP_OP_456J3_131_2158_n28, S => C431_DATA4_6);
   DP_OP_456J3_131_2158_U35 : HA_X1 port map( A => DP_OP_456J3_131_2158_n28, B 
                           => DP_OP_456J3_131_2158_n72, CO => 
                           DP_OP_456J3_131_2158_n27, S => C431_DATA4_7);
   DP_OP_456J3_131_2158_U34 : HA_X1 port map( A => DP_OP_456J3_131_2158_n27, B 
                           => DP_OP_456J3_131_2158_n73, CO => 
                           DP_OP_456J3_131_2158_n26, S => C431_DATA4_8);
   DP_OP_456J3_131_2158_U33 : HA_X1 port map( A => DP_OP_456J3_131_2158_n26, B 
                           => DP_OP_456J3_131_2158_n74, CO => 
                           DP_OP_456J3_131_2158_n25, S => C431_DATA4_9);
   DP_OP_456J3_131_2158_U32 : HA_X1 port map( A => DP_OP_456J3_131_2158_n25, B 
                           => DP_OP_456J3_131_2158_n75, CO => 
                           DP_OP_456J3_131_2158_n24, S => C431_DATA4_10);
   DP_OP_456J3_131_2158_U31 : HA_X1 port map( A => DP_OP_456J3_131_2158_n24, B 
                           => DP_OP_456J3_131_2158_n76, CO => 
                           DP_OP_456J3_131_2158_n23, S => C431_DATA4_11);
   DP_OP_456J3_131_2158_U30 : HA_X1 port map( A => DP_OP_456J3_131_2158_n23, B 
                           => DP_OP_456J3_131_2158_n77, CO => 
                           DP_OP_456J3_131_2158_n22, S => C431_DATA4_12);
   DP_OP_456J3_131_2158_U29 : HA_X1 port map( A => DP_OP_456J3_131_2158_n22, B 
                           => DP_OP_456J3_131_2158_n78, CO => 
                           DP_OP_456J3_131_2158_n21, S => C431_DATA4_13);
   DP_OP_456J3_131_2158_U28 : HA_X1 port map( A => DP_OP_456J3_131_2158_n21, B 
                           => DP_OP_456J3_131_2158_n79, CO => 
                           DP_OP_456J3_131_2158_n20, S => C431_DATA4_14);
   DP_OP_456J3_131_2158_U27 : HA_X1 port map( A => DP_OP_456J3_131_2158_n20, B 
                           => DP_OP_456J3_131_2158_n80, CO => 
                           DP_OP_456J3_131_2158_n19, S => C431_DATA4_15);
   DP_OP_456J3_131_2158_U26 : HA_X1 port map( A => DP_OP_456J3_131_2158_n19, B 
                           => DP_OP_456J3_131_2158_n81, CO => 
                           DP_OP_456J3_131_2158_n18, S => C431_DATA4_16);
   DP_OP_456J3_131_2158_U25 : HA_X1 port map( A => DP_OP_456J3_131_2158_n18, B 
                           => DP_OP_456J3_131_2158_n82, CO => 
                           DP_OP_456J3_131_2158_n17, S => C431_DATA4_17);
   intadd_0_U28 : FA_X1 port map( A => intadd_0_A_0_port, B => 
                           intadd_0_B_0_port, CI => intadd_0_CI, CO => 
                           intadd_0_n27, S => intadd_0_SUM_0_port);
   intadd_0_U27 : FA_X1 port map( A => intadd_0_A_1_port, B => 
                           intadd_0_B_1_port, CI => intadd_0_n27, CO => 
                           intadd_0_n26, S => intadd_0_SUM_1_port);
   intadd_0_U26 : FA_X1 port map( A => intadd_0_A_2_port, B => 
                           intadd_0_B_2_port, CI => intadd_0_n26, CO => 
                           intadd_0_n25, S => intadd_0_SUM_2_port);
   intadd_0_U25 : FA_X1 port map( A => intadd_0_A_3_port, B => 
                           intadd_0_B_3_port, CI => intadd_0_n25, CO => 
                           intadd_0_n24, S => intadd_0_SUM_3_port);
   intadd_0_U24 : FA_X1 port map( A => intadd_0_A_4_port, B => 
                           intadd_0_B_4_port, CI => intadd_0_n24, CO => 
                           intadd_0_n23, S => intadd_0_SUM_4_port);
   intadd_0_U23 : FA_X1 port map( A => intadd_0_A_5_port, B => 
                           intadd_0_B_5_port, CI => intadd_0_n23, CO => 
                           intadd_0_n22, S => intadd_0_SUM_5_port);
   intadd_0_U22 : FA_X1 port map( A => intadd_0_A_6_port, B => 
                           intadd_0_B_6_port, CI => intadd_0_n22, CO => 
                           intadd_0_n21, S => intadd_0_SUM_6_port);
   intadd_0_U21 : FA_X1 port map( A => intadd_0_A_7_port, B => 
                           intadd_0_B_7_port, CI => intadd_0_n21, CO => 
                           intadd_0_n20, S => intadd_0_SUM_7_port);
   intadd_0_U20 : FA_X1 port map( A => intadd_0_A_8_port, B => 
                           intadd_0_B_8_port, CI => intadd_0_n20, CO => 
                           intadd_0_n19, S => intadd_0_SUM_8_port);
   intadd_0_U19 : FA_X1 port map( A => intadd_0_A_9_port, B => 
                           intadd_0_B_9_port, CI => intadd_0_n19, CO => 
                           intadd_0_n18, S => intadd_0_SUM_9_port);
   intadd_0_U18 : FA_X1 port map( A => intadd_0_A_10_port, B => 
                           intadd_0_B_10_port, CI => intadd_0_n18, CO => 
                           intadd_0_n17, S => intadd_0_SUM_10_port);
   intadd_0_U17 : FA_X1 port map( A => intadd_0_A_11_port, B => 
                           intadd_0_B_11_port, CI => intadd_0_n17, CO => 
                           intadd_0_n16, S => intadd_0_SUM_11_port);
   intadd_0_U16 : FA_X1 port map( A => intadd_0_A_12_port, B => 
                           intadd_0_B_12_port, CI => intadd_0_n16, CO => 
                           intadd_0_n15, S => intadd_0_SUM_12_port);
   intadd_0_U15 : FA_X1 port map( A => intadd_0_A_16_port, B => 
                           intadd_0_B_13_port, CI => intadd_0_n15, CO => 
                           intadd_0_n14, S => intadd_0_SUM_13_port);
   intadd_0_U14 : FA_X1 port map( A => intadd_0_A_16_port, B => 
                           intadd_0_B_14_port, CI => intadd_0_n14, CO => 
                           intadd_0_n13, S => intadd_0_SUM_14_port);
   intadd_0_U13 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n13, CO => intadd_0_n12, S => 
                           intadd_0_SUM_15_port);
   intadd_0_U12 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n12, CO => intadd_0_n11, S => 
                           intadd_0_SUM_16_port);
   intadd_0_U11 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n11, CO => intadd_0_n10, S => 
                           intadd_0_SUM_17_port);
   intadd_0_U10 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n10, CO => intadd_0_n9, S => 
                           intadd_0_SUM_18_port);
   intadd_0_U9 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n9, CO => intadd_0_n8, S => 
                           intadd_0_SUM_19_port);
   intadd_0_U8 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n8, CO => intadd_0_n7, S => 
                           intadd_0_SUM_20_port);
   intadd_0_U7 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n7, CO => intadd_0_n6, S => 
                           intadd_0_SUM_21_port);
   intadd_0_U6 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n6, CO => intadd_0_n5, S => 
                           intadd_0_SUM_22_port);
   intadd_0_U5 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n5, CO => intadd_0_n4, S => 
                           intadd_0_SUM_23_port);
   intadd_0_U4 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n4, CO => intadd_0_n3, S => 
                           intadd_0_SUM_24_port);
   intadd_0_U3 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n3, CO => intadd_0_n2, S => 
                           intadd_0_SUM_25_port);
   intadd_0_U2 : FA_X1 port map( A => intadd_0_A_16_port, B => n62, CI => 
                           intadd_0_n2, CO => intadd_0_n1, S => 
                           intadd_0_SUM_26_port);
   intadd_1_U26 : FA_X1 port map( A => intadd_1_A_0_port, B => 
                           intadd_1_B_0_port, CI => intadd_0_SUM_2_port, CO => 
                           intadd_1_n25, S => intadd_1_SUM_0_port);
   intadd_1_U25 : FA_X1 port map( A => intadd_0_SUM_3_port, B => 
                           intadd_1_B_1_port, CI => intadd_1_n25, CO => 
                           intadd_1_n24, S => intadd_1_SUM_1_port);
   intadd_1_U24 : FA_X1 port map( A => intadd_0_SUM_4_port, B => 
                           intadd_1_B_2_port, CI => intadd_1_n24, CO => 
                           intadd_1_n23, S => intadd_1_SUM_2_port);
   intadd_1_U23 : FA_X1 port map( A => intadd_0_SUM_5_port, B => 
                           intadd_1_B_3_port, CI => intadd_1_n23, CO => 
                           intadd_1_n22, S => intadd_1_SUM_3_port);
   intadd_1_U22 : FA_X1 port map( A => intadd_0_SUM_6_port, B => 
                           intadd_1_B_4_port, CI => intadd_1_n22, CO => 
                           intadd_1_n21, S => intadd_1_SUM_4_port);
   intadd_1_U21 : FA_X1 port map( A => intadd_0_SUM_7_port, B => 
                           intadd_1_B_5_port, CI => intadd_1_n21, CO => 
                           intadd_1_n20, S => intadd_1_SUM_5_port);
   intadd_1_U20 : FA_X1 port map( A => intadd_0_SUM_8_port, B => 
                           intadd_1_B_6_port, CI => intadd_1_n20, CO => 
                           intadd_1_n19, S => intadd_1_SUM_6_port);
   intadd_1_U19 : FA_X1 port map( A => intadd_0_SUM_9_port, B => 
                           intadd_1_B_7_port, CI => intadd_1_n19, CO => 
                           intadd_1_n18, S => intadd_1_SUM_7_port);
   intadd_1_U18 : FA_X1 port map( A => intadd_0_SUM_10_port, B => 
                           intadd_1_B_8_port, CI => intadd_1_n18, CO => 
                           intadd_1_n17, S => intadd_1_SUM_8_port);
   intadd_1_U17 : FA_X1 port map( A => intadd_0_SUM_11_port, B => 
                           intadd_1_B_9_port, CI => intadd_1_n17, CO => 
                           intadd_1_n16, S => intadd_1_SUM_9_port);
   intadd_1_U16 : FA_X1 port map( A => intadd_0_SUM_12_port, B => 
                           intadd_1_B_10_port, CI => intadd_1_n16, CO => 
                           intadd_1_n15, S => intadd_1_SUM_10_port);
   intadd_1_U15 : FA_X1 port map( A => intadd_0_SUM_13_port, B => 
                           intadd_1_B_11_port, CI => intadd_1_n15, CO => 
                           intadd_1_n14, S => intadd_1_SUM_11_port);
   intadd_1_U14 : FA_X1 port map( A => intadd_0_SUM_14_port, B => 
                           intadd_1_B_12_port, CI => intadd_1_n14, CO => 
                           intadd_1_n13, S => intadd_1_SUM_12_port);
   intadd_1_U13 : FA_X1 port map( A => intadd_0_SUM_15_port, B => 
                           intadd_1_B_13_port, CI => intadd_1_n13, CO => 
                           intadd_1_n12, S => intadd_1_SUM_13_port);
   intadd_1_U12 : FA_X1 port map( A => intadd_0_SUM_16_port, B => 
                           intadd_1_B_14_port, CI => intadd_1_n12, CO => 
                           intadd_1_n11, S => intadd_1_SUM_14_port);
   intadd_1_U11 : FA_X1 port map( A => intadd_0_SUM_17_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n11, CO => 
                           intadd_1_n10, S => intadd_1_SUM_15_port);
   intadd_1_U10 : FA_X1 port map( A => intadd_0_SUM_18_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n10, CO => 
                           intadd_1_n9, S => intadd_1_SUM_16_port);
   intadd_1_U9 : FA_X1 port map( A => intadd_0_SUM_19_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n9, CO => 
                           intadd_1_n8, S => intadd_1_SUM_17_port);
   intadd_1_U8 : FA_X1 port map( A => intadd_0_SUM_20_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n8, CO => 
                           intadd_1_n7, S => intadd_1_SUM_18_port);
   intadd_1_U7 : FA_X1 port map( A => intadd_0_SUM_21_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n7, CO => 
                           intadd_1_n6, S => intadd_1_SUM_19_port);
   intadd_1_U6 : FA_X1 port map( A => intadd_0_SUM_22_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n6, CO => 
                           intadd_1_n5, S => intadd_1_SUM_20_port);
   intadd_1_U5 : FA_X1 port map( A => intadd_0_SUM_23_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n5, CO => 
                           intadd_1_n4, S => intadd_1_SUM_21_port);
   intadd_1_U4 : FA_X1 port map( A => intadd_0_SUM_24_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n4, CO => 
                           intadd_1_n3, S => intadd_1_SUM_22_port);
   intadd_1_U3 : FA_X1 port map( A => intadd_0_SUM_25_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n3, CO => 
                           intadd_1_n2, S => intadd_1_SUM_23_port);
   intadd_1_U2 : FA_X1 port map( A => intadd_0_SUM_26_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n2, CO => 
                           intadd_1_n1, S => intadd_1_SUM_24_port);
   intadd_2_U11 : FA_X1 port map( A => intadd_2_A_0_port, B => 
                           intadd_2_B_0_port, CI => intadd_1_SUM_2_port, CO => 
                           intadd_2_n10, S => intadd_2_SUM_0_port);
   intadd_2_U10 : FA_X1 port map( A => intadd_2_A_1_port, B => 
                           intadd_1_SUM_3_port, CI => intadd_2_n10, CO => 
                           intadd_2_n9, S => intadd_2_SUM_1_port);
   intadd_2_U9 : FA_X1 port map( A => intadd_2_A_2_port, B => 
                           intadd_1_SUM_4_port, CI => intadd_2_n9, CO => 
                           intadd_2_n8, S => intadd_2_SUM_2_port);
   intadd_2_U8 : FA_X1 port map( A => intadd_2_A_3_port, B => 
                           intadd_1_SUM_5_port, CI => intadd_2_n8, CO => 
                           intadd_2_n7, S => intadd_2_SUM_3_port);
   intadd_2_U7 : FA_X1 port map( A => intadd_2_A_4_port, B => 
                           intadd_1_SUM_6_port, CI => intadd_2_n7, CO => 
                           intadd_2_n6, S => intadd_2_SUM_4_port);
   intadd_2_U6 : FA_X1 port map( A => intadd_2_A_5_port, B => 
                           intadd_1_SUM_7_port, CI => intadd_2_n6, CO => 
                           intadd_2_n5, S => intadd_2_SUM_5_port);
   intadd_2_U5 : FA_X1 port map( A => intadd_2_A_6_port, B => 
                           intadd_1_SUM_8_port, CI => intadd_2_n5, CO => 
                           intadd_2_n4, S => intadd_2_SUM_6_port);
   intadd_2_U4 : FA_X1 port map( A => intadd_2_A_7_port, B => 
                           intadd_1_SUM_9_port, CI => intadd_2_n4, CO => 
                           intadd_2_n3, S => intadd_2_SUM_7_port);
   intadd_2_U3 : FA_X1 port map( A => intadd_2_A_8_port, B => 
                           intadd_1_SUM_10_port, CI => intadd_2_n3, CO => 
                           intadd_2_n2, S => intadd_2_SUM_8_port);
   intadd_2_U2 : FA_X1 port map( A => intadd_2_A_9_port, B => 
                           intadd_1_SUM_11_port, CI => intadd_2_n2, CO => 
                           intadd_2_n1, S => intadd_2_SUM_9_port);
   OP_A_reg_7_inst : DLH_X1 port map( G => N246, D => OP1(7), Q => OP_A_7_port)
                           ;
   OP_A_reg_12_inst : DLH_X1 port map( G => n1412, D => OP1(12), Q => 
                           OP_A_12_port);
   OP_A_reg_13_inst : DLH_X1 port map( G => n1412, D => OP1(13), Q => 
                           OP_A_13_port);
   OP_A_reg_10_inst : DLH_X1 port map( G => n1412, D => OP1(10), Q => 
                           OP_A_10_port);
   OP_A_reg_0_inst : DLH_X1 port map( G => n1412, D => OP1(0), Q => OP_A_0_port
                           );
   OP_A_reg_4_inst : DLH_X1 port map( G => N246, D => OP1(4), Q => OP_A_4_port)
                           ;
   OP_A_reg_8_inst : DLH_X1 port map( G => n1412, D => OP1(8), Q => OP_A_8_port
                           );
   OP_A_reg_6_inst : DLH_X1 port map( G => N246, D => OP1(6), Q => OP_A_6_port)
                           ;
   OP_A_reg_11_inst : DLH_X1 port map( G => n1412, D => OP1(11), Q => 
                           OP_A_11_port);
   OP_A_reg_14_inst : DLH_X1 port map( G => n1412, D => OP1(14), Q => 
                           OP_A_14_port);
   OP_A_reg_1_inst : DLH_X1 port map( G => N246, D => OP1(1), Q => OP_A_1_port)
                           ;
   OP_A_reg_3_inst : DLH_X1 port map( G => N246, D => OP1(3), Q => OP_A_3_port)
                           ;
   OP_A_reg_9_inst : DLH_X1 port map( G => n1412, D => OP1(9), Q => OP_A_9_port
                           );
   OP_A_reg_5_inst : DLH_X1 port map( G => n1412, D => OP1(5), Q => OP_A_5_port
                           );
   OP_B_reg_2_inst : DLH_X1 port map( G => N246, D => N249, Q => OP_B_2_port);
   OP_B_reg_5_inst : DLH_X1 port map( G => n1412, D => N252, Q => OP_B_5_port);
   OP_B_reg_3_inst : DLH_X1 port map( G => N246, D => N250, Q => OP_B_3_port);
   OP_A_reg_15_inst : DLH_X1 port map( G => n1412, D => OP1(15), Q => 
                           OP_A_15_port);
   OP_B_reg_4_inst : DLH_X1 port map( G => N246, D => N251, Q => OP_B_4_port);
   OP_A_reg_2_inst : DLH_X1 port map( G => N246, D => OP1(2), Q => OP_A_2_port)
                           ;
   OP_B_reg_1_inst : DLH_X2 port map( G => N246, D => N248, Q => OP_B_1_port);
   U3 : CLKBUF_X1 port map( A => n148, Z => n60);
   U4 : INV_X1 port map( A => n1368, ZN => n1367);
   U5 : INV_X1 port map( A => n1245, ZN => n1369);
   U6 : INV_X1 port map( A => n1372, ZN => n1344);
   U7 : INV_X2 port map( A => n578, ZN => n55);
   U8 : INV_X2 port map( A => n608, ZN => n56);
   U9 : INV_X2 port map( A => N280, ZN => n196);
   U10 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_15, B1 => 
                           OP_A_11_port, B2 => n159, C1 => n160, C2 => 
                           OP_A_10_port, ZN => intadd_1_B_9_port);
   U11 : AOI211_X1 port map( C1 => n64, C2 => n864, A => n541, B => n540, ZN =>
                           n965);
   U12 : NOR2_X2 port map( A1 => DP_OP_446J3_125_4819_n12, A2 => n1092, ZN => 
                           n57);
   U13 : OR2_X1 port map( A1 => n145, A2 => n114, ZN => n58);
   U14 : OR3_X1 port map( A1 => n1082, A2 => OP_B_7_port, A3 => n161, ZN => n59
                           );
   U15 : NOR2_X2 port map( A1 => OP_B_2_port, A2 => n1160, ZN => n856);
   U16 : NOR2_X2 port map( A1 => OP_B_7_port, A2 => n162, ZN => n1028);
   U17 : NOR2_X2 port map( A1 => n224, A2 => n743, ZN => n147);
   U18 : NOR2_X2 port map( A1 => OP_B_5_port, A2 => n154, ZN => n160);
   U19 : AOI21_X2 port map( B1 => OP_B_3_port, B2 => OP_B_4_port, A => n297, ZN
                           => n1413);
   U20 : NOR2_X2 port map( A1 => OP_B_3_port, A2 => OP_B_2_port, ZN => n895);
   U21 : INV_X1 port map( A => n59, ZN => n61);
   U22 : INV_X1 port map( A => n58, ZN => n62);
   U23 : NOR2_X2 port map( A1 => n901, A2 => n1261, ZN => n1228);
   U24 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n582, ZN => n63);
   U25 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n582, ZN => n64);
   U26 : NOR2_X2 port map( A1 => n1381, A2 => n111, ZN => intadd_1_B_18_port);
   U27 : AOI21_X2 port map( B1 => OP_B_2_port, B2 => OP_B_1_port, A => n1160, 
                           ZN => n1415);
   U28 : NOR3_X4 port map( A1 => n150, A2 => OP_B_5_port, A3 => n153, ZN => 
                           n159);
   U29 : NOR2_X4 port map( A1 => n126, A2 => n109, ZN => intadd_0_A_16_port);
   U30 : NOR3_X4 port map( A1 => n1082, A2 => OP_B_7_port, A3 => n1081, ZN => 
                           n1380);
   U31 : OR2_X1 port map( A1 => n1413, A2 => n1381, ZN => n65);
   U32 : INV_X1 port map( A => OPC(4), ZN => n69);
   U33 : NOR2_X1 port map( A1 => OPC(2), A2 => OPC(1), ZN => n72);
   U34 : INV_X1 port map( A => OPC(6), ZN => n171);
   U35 : NOR3_X1 port map( A1 => OPC(5), A2 => n69, A3 => n171, ZN => n80);
   U36 : NAND2_X1 port map( A1 => OPC(4), A2 => OPC(5), ZN => n81);
   U37 : NOR2_X1 port map( A1 => OPC(6), A2 => n81, ZN => n77);
   U38 : NOR2_X1 port map( A1 => n80, A2 => n77, ZN => n176);
   U39 : INV_X1 port map( A => OPC(3), ZN => n66);
   U40 : INV_X1 port map( A => OPC(0), ZN => n67);
   U41 : NAND3_X1 port map( A1 => n72, A2 => n66, A3 => n67, ZN => n96_port);
   U42 : INV_X1 port map( A => OPC(5), ZN => n68);
   U43 : NAND2_X1 port map( A1 => n69, A2 => n68, ZN => n216);
   U44 : NOR2_X1 port map( A1 => OPC(3), A2 => n67, ZN => n83);
   U45 : NAND2_X1 port map( A1 => n72, A2 => n83, ZN => n1411);
   U46 : OAI22_X1 port map( A1 => n176, A2 => n96_port, B1 => n216, B2 => n1411
                           , ZN => N280);
   U47 : NOR2_X1 port map( A1 => OPC(4), A2 => n68, ZN => n88);
   U48 : NAND2_X1 port map( A1 => n88, A2 => n171, ZN => n172);
   U49 : NOR3_X1 port map( A1 => OPC(6), A2 => OPC(5), A3 => n69, ZN => n100);
   U50 : INV_X1 port map( A => n100, ZN => n1410);
   U51 : NAND3_X1 port map( A1 => OPC(3), A2 => OPC(0), A3 => n72, ZN => n215);
   U52 : OAI22_X1 port map( A1 => n172, A2 => n96_port, B1 => n1410, B2 => n215
                           , ZN => N96);
   U53 : NAND3_X1 port map( A1 => OPC(6), A2 => OPC(5), A3 => n69, ZN => n1406)
                           ;
   U54 : INV_X1 port map( A => n96_port, ZN => n102);
   U55 : INV_X1 port map( A => n216, ZN => n101);
   U56 : NAND2_X1 port map( A1 => OPC(6), A2 => n101, ZN => n1409);
   U57 : INV_X1 port map( A => n1409, ZN => n70);
   U58 : AOI21_X1 port map( B1 => n102, B2 => n70, A => N96, ZN => n71);
   U59 : OAI21_X1 port map( B1 => n1406, B2 => n215, A => n71, ZN => N284);
   U60 : NAND2_X1 port map( A1 => OPC(3), A2 => n72, ZN => n73);
   U61 : NOR2_X1 port map( A1 => OPC(0), A2 => n73, ZN => n86);
   U62 : INV_X1 port map( A => n86, ZN => n1408);
   U63 : INV_X1 port map( A => n215, ZN => n78);
   U64 : NAND2_X1 port map( A1 => OPC(2), A2 => OPC(3), ZN => n74);
   U65 : NOR2_X1 port map( A1 => OPC(0), A2 => n74, ZN => n94);
   U66 : INV_X1 port map( A => OPC(1), ZN => n104);
   U67 : INV_X1 port map( A => OPC(2), ZN => n75);
   U68 : NAND3_X1 port map( A1 => OPC(1), A2 => n83, A3 => n75, ZN => n93);
   U69 : INV_X1 port map( A => n93, ZN => n76);
   U70 : AOI21_X1 port map( B1 => n94, B2 => n104, A => n76, ZN => n179);
   U71 : NOR2_X1 port map( A1 => OPC(4), A2 => n179, ZN => n169);
   U72 : AOI21_X1 port map( B1 => n78, B2 => n77, A => n169, ZN => n79);
   U73 : OAI21_X1 port map( B1 => n1406, B2 => n1408, A => n79, ZN => N286);
   U74 : INV_X1 port map( A => n80, ZN => n217);
   U75 : AOI21_X1 port map( B1 => n172, B2 => n217, A => n1408, ZN => n84);
   U76 : NAND2_X1 port map( A1 => OPC(4), A2 => n171, ZN => n82);
   U77 : OR2_X1 port map( A1 => n171, A2 => n81, ZN => n90);
   U78 : OAI22_X1 port map( A1 => n82, A2 => n1408, B1 => n215, B2 => n90, ZN 
                           => n168);
   U79 : NAND3_X1 port map( A1 => OPC(2), A2 => n83, A3 => n104, ZN => n92);
   U80 : OAI22_X1 port map( A1 => n172, A2 => n92, B1 => n1408, B2 => n90, ZN 
                           => n177);
   U81 : NOR4_X1 port map( A1 => n84, A2 => n168, A3 => N286, A4 => n177, ZN =>
                           n85);
   U82 : OR2_X1 port map( A1 => n216, A2 => n92, ZN => n174);
   U83 : OAI211_X1 port map( C1 => n215, C2 => n217, A => n85, B => n174, ZN =>
                           N285);
   U84 : NAND2_X1 port map( A1 => n101, A2 => n86, ZN => n1407);
   U85 : INV_X1 port map( A => n1411, ZN => n87);
   U86 : OAI21_X1 port map( B1 => n88, B2 => n100, A => n87, ZN => n89);
   U87 : OAI211_X1 port map( C1 => n96_port, C2 => n90, A => n1407, B => n89, 
                           ZN => N281);
   U88 : NAND3_X1 port map( A1 => OPC(2), A2 => OPC(3), A3 => OPC(0), ZN => n91
                           );
   U89 : OAI211_X1 port map( C1 => OPC(1), C2 => n91, A => n93, B => n96_port, 
                           ZN => n99);
   U90 : AOI21_X1 port map( B1 => n93, B2 => n92, A => n217, ZN => n98);
   U91 : NAND3_X1 port map( A1 => OPC(5), A2 => OPC(1), A3 => n94, ZN => n95);
   U92 : OAI21_X1 port map( B1 => n96_port, B2 => n1406, A => n95, ZN => n97);
   U93 : AOI211_X1 port map( C1 => n100, C2 => n99, A => n98, B => n97, ZN => 
                           n115);
   U94 : INV_X1 port map( A => N281, ZN => n219);
   U95 : NAND3_X1 port map( A1 => n102, A2 => n101, A3 => n171, ZN => n103);
   U96 : OAI21_X1 port map( B1 => n215, B2 => n172, A => n103, ZN => n1366);
   U97 : INV_X1 port map( A => n1366, ZN => n901);
   U98 : INV_X1 port map( A => n172, ZN => n106);
   U99 : AOI211_X1 port map( C1 => OPC(3), C2 => OPC(2), A => OPC(0), B => n104
                           , ZN => n105);
   U100 : OAI211_X1 port map( C1 => OPC(2), C2 => OPC(3), A => n106, B => n105,
                           ZN => n1396);
   U101 : NAND4_X1 port map( A1 => n115, A2 => n219, A3 => n901, A4 => n1396, 
                           ZN => n107);
   U102 : NOR3_X2 port map( A1 => N284, A2 => N285, A3 => n107, ZN => n194);
   U103 : CLKBUF_X1 port map( A => n194, Z => n205);
   U104 : NAND2_X1 port map( A1 => n196, A2 => n205, ZN => N246);
   U105 : CLKBUF_X1 port map( A => N246, Z => n1412);
   U106 : INV_X1 port map( A => OP_A_15_port, ZN => n1081);
   U107 : INV_X1 port map( A => OP_B_1_port, ZN => n224);
   U108 : INV_X1 port map( A => OP_B_0_port, ZN => n223);
   U109 : OR2_X1 port map( A1 => OP_B_1_port, A2 => n223, ZN => n510);
   U110 : NOR2_X1 port map( A1 => n1081, A2 => n510, ZN => n126);
   U111 : NOR2_X1 port map( A1 => OP_B_0_port, A2 => n224, ZN => n604);
   U112 : INV_X1 port map( A => n604, ZN => n576);
   U113 : OR2_X1 port map( A1 => n224, A2 => n223, ZN => n578);
   U114 : NAND2_X1 port map( A1 => n55, A2 => n1081, ZN => n116);
   U115 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n576, A => n116, ZN => 
                           n108);
   U116 : INV_X1 port map( A => n108, ZN => n123);
   U117 : NOR2_X1 port map( A1 => DP_OP_440J3_122_9847_n20, A2 => n123, ZN => 
                           n109);
   U118 : INV_X1 port map( A => OP_B_7_port, ZN => n295);
   U119 : AOI21_X1 port map( B1 => OP_B_6_port, B2 => OP_B_5_port, A => n295, 
                           ZN => n1414);
   U120 : INV_X1 port map( A => OP_B_5_port, ZN => n297);
   U121 : INV_X1 port map( A => OP_B_3_port, ZN => n1160);
   U122 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => OP_B_3_port, ZN => n150);
   U123 : NOR3_X1 port map( A1 => n150, A2 => OP_B_5_port, A3 => n1081, ZN => 
                           n1381);
   U124 : NAND2_X1 port map( A1 => n150, A2 => OP_B_5_port, ZN => n121);
   U125 : INV_X1 port map( A => OP_B_4_port, ZN => n1363);
   U126 : NOR2_X1 port map( A1 => n1160, A2 => n1363, ZN => n153);
   U127 : NOR3_X1 port map( A1 => n150, A2 => n153, A3 => n297, ZN => n151);
   U128 : NAND2_X1 port map( A1 => n151, A2 => n1081, ZN => n120);
   U129 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n121, A => n120, ZN => 
                           n110);
   U130 : INV_X1 port map( A => n110, ZN => n157);
   U131 : OR2_X1 port map( A1 => DP_OP_451J3_128_3502_n15, A2 => n157, ZN => 
                           n1383);
   U132 : INV_X1 port map( A => n1383, ZN => n111);
   U133 : INV_X1 port map( A => OP_B_2_port, ZN => n582);
   U134 : AOI211_X1 port map( C1 => n582, C2 => n224, A => OP_B_3_port, B => 
                           n1081, ZN => n145);
   U135 : NAND2_X1 port map( A1 => n856, A2 => n224, ZN => n118);
   U136 : NAND2_X1 port map( A1 => OP_B_3_port, A2 => OP_B_2_port, ZN => n858);
   U137 : NAND2_X1 port map( A1 => OP_B_1_port, A2 => n856, ZN => n112);
   U138 : OAI21_X1 port map( B1 => OP_B_1_port, B2 => n858, A => n112, ZN => 
                           n137);
   U139 : NAND2_X1 port map( A1 => n1081, A2 => n137, ZN => n117);
   U140 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n118, A => n117, ZN => 
                           n113);
   U141 : INV_X1 port map( A => n113, ZN => n142);
   U142 : NOR2_X1 port map( A1 => DP_OP_456J3_131_2158_n17, A2 => n142, ZN => 
                           n114);
   U143 : NAND2_X1 port map( A1 => n196, A2 => n115, ZN => N279);
   U144 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n576, A => n116, ZN => 
                           DP_OP_440J3_122_9847_n80);
   U145 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n578, B1 => OP_A_13_port
                           , B2 => n576, ZN => DP_OP_440J3_122_9847_n79);
   U146 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n578, B1 => OP_A_12_port
                           , B2 => n576, ZN => DP_OP_440J3_122_9847_n78);
   U147 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n576, B1 => OP_A_12_port
                           , B2 => n578, ZN => DP_OP_440J3_122_9847_n77);
   U148 : OAI22_X1 port map( A1 => OP_A_10_port, A2 => n576, B1 => OP_A_11_port
                           , B2 => n578, ZN => DP_OP_440J3_122_9847_n76);
   U149 : OAI22_X1 port map( A1 => OP_A_9_port, A2 => n576, B1 => OP_A_10_port,
                           B2 => n578, ZN => DP_OP_440J3_122_9847_n75);
   U150 : OAI22_X1 port map( A1 => OP_A_8_port, A2 => n576, B1 => OP_A_9_port, 
                           B2 => n578, ZN => DP_OP_440J3_122_9847_n74);
   U151 : OAI22_X1 port map( A1 => OP_A_7_port, A2 => n576, B1 => OP_A_8_port, 
                           B2 => n578, ZN => DP_OP_440J3_122_9847_n73);
   U152 : OAI22_X1 port map( A1 => OP_A_6_port, A2 => n576, B1 => OP_A_7_port, 
                           B2 => n578, ZN => DP_OP_440J3_122_9847_n72);
   U153 : OAI22_X1 port map( A1 => OP_A_5_port, A2 => n576, B1 => OP_A_6_port, 
                           B2 => n578, ZN => DP_OP_440J3_122_9847_n71);
   U154 : OAI22_X1 port map( A1 => OP_A_4_port, A2 => n576, B1 => OP_A_5_port, 
                           B2 => n578, ZN => DP_OP_440J3_122_9847_n70);
   U155 : OAI22_X1 port map( A1 => OP_A_3_port, A2 => n576, B1 => OP_A_4_port, 
                           B2 => n578, ZN => DP_OP_440J3_122_9847_n69);
   U156 : OAI22_X1 port map( A1 => OP_A_2_port, A2 => n576, B1 => OP_A_3_port, 
                           B2 => n578, ZN => DP_OP_440J3_122_9847_n68);
   U157 : OAI22_X1 port map( A1 => OP_A_2_port, A2 => n578, B1 => OP_A_1_port, 
                           B2 => n576, ZN => DP_OP_440J3_122_9847_n67);
   U158 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n578, B1 => OP_A_0_port, 
                           B2 => n576, ZN => DP_OP_440J3_122_9847_n66);
   U159 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n578, A => n576, ZN => 
                           DP_OP_440J3_122_9847_n35);
   U160 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n118, A => n117, ZN => 
                           DP_OP_456J3_131_2158_n82);
   U161 : INV_X1 port map( A => n137, ZN => n119);
   U162 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n119, B1 => OP_A_13_port
                           , B2 => n118, ZN => DP_OP_456J3_131_2158_n81);
   U163 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n119, B1 => OP_A_12_port
                           , B2 => n118, ZN => DP_OP_456J3_131_2158_n80);
   U164 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n118, B1 => OP_A_12_port
                           , B2 => n119, ZN => DP_OP_456J3_131_2158_n79);
   U165 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n119, B1 => OP_A_10_port
                           , B2 => n118, ZN => DP_OP_456J3_131_2158_n78);
   U166 : OAI22_X1 port map( A1 => n119, A2 => OP_A_10_port, B1 => OP_A_9_port,
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n77);
   U167 : OAI22_X1 port map( A1 => n119, A2 => OP_A_9_port, B1 => OP_A_8_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n76);
   U168 : OAI22_X1 port map( A1 => n119, A2 => OP_A_8_port, B1 => OP_A_7_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n75);
   U169 : OAI22_X1 port map( A1 => n119, A2 => OP_A_7_port, B1 => OP_A_6_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n74);
   U170 : OAI22_X1 port map( A1 => n119, A2 => OP_A_6_port, B1 => OP_A_5_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n73);
   U171 : OAI22_X1 port map( A1 => n119, A2 => OP_A_5_port, B1 => OP_A_4_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n72);
   U172 : OAI22_X1 port map( A1 => n119, A2 => OP_A_4_port, B1 => OP_A_3_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n71);
   U173 : OAI22_X1 port map( A1 => n119, A2 => OP_A_3_port, B1 => OP_A_2_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n70);
   U174 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n118, B1 => n119, B2 => 
                           OP_A_2_port, ZN => DP_OP_456J3_131_2158_n69);
   U175 : OAI22_X1 port map( A1 => n119, A2 => OP_A_1_port, B1 => OP_A_0_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n68);
   U176 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n119, A => n118, ZN => 
                           DP_OP_456J3_131_2158_n67);
   U177 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n121, A => n120, ZN => 
                           DP_OP_451J3_128_3502_n85);
   U178 : INV_X1 port map( A => n151, ZN => n122);
   U179 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n122, B1 => OP_A_13_port
                           , B2 => n121, ZN => DP_OP_451J3_128_3502_n84);
   U180 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n122, B1 => OP_A_12_port
                           , B2 => n121, ZN => DP_OP_451J3_128_3502_n83);
   U181 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n121, B1 => OP_A_12_port
                           , B2 => n122, ZN => DP_OP_451J3_128_3502_n82);
   U182 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n122, B1 => OP_A_10_port
                           , B2 => n121, ZN => DP_OP_451J3_128_3502_n81);
   U183 : OAI22_X1 port map( A1 => OP_A_10_port, A2 => n122, B1 => OP_A_9_port,
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n80);
   U184 : OAI22_X1 port map( A1 => OP_A_9_port, A2 => n122, B1 => OP_A_8_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n79);
   U185 : OAI22_X1 port map( A1 => OP_A_8_port, A2 => n122, B1 => OP_A_7_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n78);
   U186 : OAI22_X1 port map( A1 => OP_A_7_port, A2 => n122, B1 => OP_A_6_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n77);
   U187 : OAI22_X1 port map( A1 => OP_A_6_port, A2 => n122, B1 => OP_A_5_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n76);
   U188 : OAI22_X1 port map( A1 => OP_A_5_port, A2 => n122, B1 => OP_A_4_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n75);
   U189 : OAI22_X1 port map( A1 => OP_A_4_port, A2 => n122, B1 => OP_A_3_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n74);
   U190 : OAI22_X1 port map( A1 => OP_A_3_port, A2 => n122, B1 => OP_A_2_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n73);
   U191 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n121, B1 => OP_A_2_port, 
                           B2 => n122, ZN => DP_OP_451J3_128_3502_n72);
   U192 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n122, B1 => OP_A_0_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n71);
   U193 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n122, A => n121, ZN => 
                           DP_OP_451J3_128_3502_n70);
   U194 : XNOR2_X1 port map( A => DP_OP_440J3_122_9847_n20, B => n123, ZN => 
                           n124);
   U195 : INV_X1 port map( A => n126, ZN => n891);
   U196 : NAND2_X1 port map( A1 => n224, A2 => n891, ZN => n125);
   U197 : OAI21_X1 port map( B1 => n126, B2 => n124, A => n125, ZN => 
                           intadd_0_A_12_port);
   U198 : OAI21_X1 port map( B1 => n126, B2 => C428_DATA4_15, A => n125, ZN => 
                           intadd_0_A_11_port);
   U199 : INV_X1 port map( A => n510, ZN => n543);
   U200 : NAND2_X1 port map( A1 => n543, A2 => OP_A_14_port, ZN => n853);
   U201 : INV_X1 port map( A => n853, ZN => n127);
   U202 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_14, A => n127,
                           ZN => intadd_0_A_10_port);
   U203 : INV_X1 port map( A => n510, ZN => n492);
   U204 : NAND2_X1 port map( A1 => n492, A2 => OP_A_13_port, ZN => n820);
   U205 : INV_X1 port map( A => n820, ZN => n128);
   U206 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_13, A => n128,
                           ZN => intadd_0_A_9_port);
   U207 : NAND2_X1 port map( A1 => n543, A2 => OP_A_12_port, ZN => n805);
   U208 : INV_X1 port map( A => n805, ZN => n129);
   U209 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_12, A => n129,
                           ZN => intadd_0_A_8_port);
   U210 : NAND2_X1 port map( A1 => n543, A2 => OP_A_11_port, ZN => n770);
   U211 : INV_X1 port map( A => n770, ZN => n130);
   U212 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_11, A => n130,
                           ZN => intadd_0_A_7_port);
   U213 : NAND2_X1 port map( A1 => n543, A2 => OP_A_10_port, ZN => n741);
   U214 : INV_X1 port map( A => n741, ZN => n131);
   U215 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_10, A => n131,
                           ZN => intadd_0_A_6_port);
   U216 : NAND2_X1 port map( A1 => n492, A2 => OP_A_9_port, ZN => n727);
   U217 : INV_X1 port map( A => n727, ZN => n132);
   U218 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_9, A => n132, 
                           ZN => intadd_0_A_5_port);
   U219 : NAND2_X1 port map( A1 => n543, A2 => OP_A_8_port, ZN => n697);
   U220 : INV_X1 port map( A => n697, ZN => n133);
   U221 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_8, A => n133, 
                           ZN => intadd_0_A_4_port);
   U222 : NAND2_X1 port map( A1 => n543, A2 => OP_A_7_port, ZN => n676);
   U223 : INV_X1 port map( A => n676, ZN => n134);
   U224 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_7, A => n134, 
                           ZN => intadd_0_A_3_port);
   U225 : NAND2_X1 port map( A1 => n543, A2 => OP_A_6_port, ZN => n659);
   U226 : INV_X1 port map( A => n659, ZN => n135);
   U227 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_6, A => n135, 
                           ZN => intadd_0_A_2_port);
   U228 : NAND2_X1 port map( A1 => n492, A2 => OP_A_5_port, ZN => n629);
   U229 : INV_X1 port map( A => n629, ZN => n136);
   U230 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_5, A => n136, 
                           ZN => intadd_0_A_1_port);
   U231 : INV_X1 port map( A => n895, ZN => n766);
   U232 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n582, ZN => n854);
   U233 : INV_X1 port map( A => n854, ZN => n743);
   U234 : AOI22_X1 port map( A1 => OP_B_1_port, A2 => n766, B1 => n743, B2 => 
                           n224, ZN => n148);
   U235 : AND2_X1 port map( A1 => n137, A2 => C2_DATA1_2, ZN => n138);
   U236 : AOI21_X1 port map( B1 => n60, B2 => OP_A_0_port, A => n138, ZN => 
                           n526);
   U237 : INV_X1 port map( A => OP_A_2_port, ZN => n577);
   U238 : NOR2_X1 port map( A1 => n510, A2 => n577, ZN => n553);
   U239 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_2, A => n553, 
                           ZN => n527);
   U240 : NOR2_X1 port map( A1 => n526, A2 => n527, ZN => n538);
   U241 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_3, B1 => 
                           OP_A_0_port, B2 => n147, C1 => n60, C2 => 
                           OP_A_1_port, ZN => n140);
   U242 : INV_X1 port map( A => n140, ZN => n535);
   U243 : INV_X1 port map( A => n538, ZN => n139);
   U244 : INV_X1 port map( A => OP_A_3_port, ZN => n551);
   U245 : NOR2_X1 port map( A1 => n510, A2 => n551, ZN => n581);
   U246 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_3, A => n581, 
                           ZN => n536);
   U247 : OAI21_X1 port map( B1 => n140, B2 => n139, A => n536, ZN => n141);
   U248 : OAI21_X1 port map( B1 => n538, B2 => n535, A => n141, ZN => 
                           intadd_0_A_0_port);
   U249 : XNOR2_X1 port map( A => DP_OP_456J3_131_2158_n17, B => n142, ZN => 
                           n144);
   U250 : OR2_X1 port map( A1 => n145, A2 => n1415, ZN => n143);
   U251 : OAI21_X1 port map( B1 => n145, B2 => n144, A => n143, ZN => 
                           intadd_0_B_14_port);
   U252 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_17, B1 => 
                           OP_A_15_port, B2 => n60, C1 => OP_A_14_port, C2 => 
                           n147, ZN => intadd_0_B_13_port);
   U253 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_16, B1 => 
                           OP_A_13_port, B2 => n147, C1 => OP_A_14_port, C2 => 
                           n60, ZN => intadd_0_B_12_port);
   U254 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_15, B1 => 
                           OP_A_12_port, B2 => n147, C1 => OP_A_13_port, C2 => 
                           n60, ZN => intadd_0_B_11_port);
   U255 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_14, B1 => 
                           OP_A_12_port, B2 => n60, C1 => OP_A_11_port, C2 => 
                           n147, ZN => intadd_0_B_10_port);
   U256 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_13, B1 => 
                           OP_A_11_port, B2 => n60, C1 => n147, C2 => 
                           OP_A_10_port, ZN => intadd_0_B_9_port);
   U257 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_12, B1 => n60, B2 
                           => OP_A_10_port, C1 => n147, C2 => OP_A_9_port, ZN 
                           => intadd_0_B_8_port);
   U258 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_11, B1 => n60, B2 
                           => OP_A_9_port, C1 => n147, C2 => OP_A_8_port, ZN =>
                           intadd_0_B_7_port);
   U259 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_10, B1 => n60, B2 
                           => OP_A_8_port, C1 => n147, C2 => OP_A_7_port, ZN =>
                           intadd_0_B_6_port);
   U260 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_9, B1 => n60, B2 =>
                           OP_A_7_port, C1 => n147, C2 => OP_A_6_port, ZN => 
                           intadd_0_B_5_port);
   U261 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_8, B1 => n60, B2 =>
                           OP_A_6_port, C1 => n147, C2 => OP_A_5_port, ZN => 
                           intadd_0_B_4_port);
   U262 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_7, B1 => n60, B2 =>
                           OP_A_5_port, C1 => n147, C2 => OP_A_4_port, ZN => 
                           intadd_0_B_3_port);
   U263 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_6, B1 => n60, B2 =>
                           OP_A_4_port, C1 => n147, C2 => OP_A_3_port, ZN => 
                           intadd_0_B_2_port);
   U264 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_5, B1 => n60, B2 =>
                           OP_A_3_port, C1 => n147, C2 => OP_A_2_port, ZN => 
                           intadd_0_B_1_port);
   U265 : NAND2_X1 port map( A1 => n543, A2 => OP_A_4_port, ZN => n605);
   U266 : INV_X1 port map( A => n605, ZN => n146);
   U267 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_4, A => n146, 
                           ZN => intadd_0_B_0_port);
   U268 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_4, B1 => n60, B2 =>
                           OP_A_2_port, C1 => n147, C2 => OP_A_1_port, ZN => 
                           intadd_0_CI);
   U269 : NOR2_X1 port map( A1 => OP_B_5_port, A2 => OP_B_6_port, ZN => n1082);
   U270 : NAND2_X1 port map( A1 => n1082, A2 => OP_B_7_port, ZN => n1079);
   U271 : INV_X1 port map( A => OP_B_6_port, ZN => n378);
   U272 : NOR2_X1 port map( A1 => n297, A2 => n378, ZN => n161);
   U273 : NOR3_X1 port map( A1 => n1082, A2 => n161, A3 => n295, ZN => n163);
   U274 : NAND2_X1 port map( A1 => n163, A2 => n1081, ZN => n1078);
   U275 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n1079, A => n1078, ZN =>
                           DP_OP_446J3_125_4819_n87);
   U276 : INV_X1 port map( A => n163, ZN => n149);
   U277 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n149, B1 => OP_A_13_port
                           , B2 => n1079, ZN => DP_OP_446J3_125_4819_n86);
   U278 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n149, B1 => OP_A_12_port
                           , B2 => n1079, ZN => DP_OP_446J3_125_4819_n85);
   U279 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n1079, B1 => 
                           OP_A_12_port, B2 => n149, ZN => 
                           DP_OP_446J3_125_4819_n84);
   U280 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n149, B1 => OP_A_10_port
                           , B2 => n1079, ZN => DP_OP_446J3_125_4819_n83);
   U281 : OAI22_X1 port map( A1 => OP_A_10_port, A2 => n149, B1 => OP_A_9_port,
                           B2 => n1079, ZN => DP_OP_446J3_125_4819_n82);
   U282 : OAI22_X1 port map( A1 => OP_A_9_port, A2 => n149, B1 => OP_A_8_port, 
                           B2 => n1079, ZN => DP_OP_446J3_125_4819_n81);
   U283 : OAI22_X1 port map( A1 => OP_A_8_port, A2 => n149, B1 => OP_A_7_port, 
                           B2 => n1079, ZN => DP_OP_446J3_125_4819_n80);
   U284 : OAI22_X1 port map( A1 => OP_A_7_port, A2 => n149, B1 => OP_A_6_port, 
                           B2 => n1079, ZN => DP_OP_446J3_125_4819_n79);
   U285 : OAI22_X1 port map( A1 => OP_A_6_port, A2 => n149, B1 => OP_A_5_port, 
                           B2 => n1079, ZN => DP_OP_446J3_125_4819_n78);
   U286 : OAI22_X1 port map( A1 => OP_A_5_port, A2 => n149, B1 => OP_A_4_port, 
                           B2 => n1079, ZN => DP_OP_446J3_125_4819_n77);
   U287 : OAI22_X1 port map( A1 => OP_A_4_port, A2 => n149, B1 => OP_A_3_port, 
                           B2 => n1079, ZN => DP_OP_446J3_125_4819_n76);
   U288 : OAI22_X1 port map( A1 => OP_A_3_port, A2 => n149, B1 => OP_A_2_port, 
                           B2 => n1079, ZN => DP_OP_446J3_125_4819_n75);
   U289 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n1079, B1 => OP_A_2_port,
                           B2 => n149, ZN => DP_OP_446J3_125_4819_n74);
   U290 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n149, B1 => OP_A_0_port, 
                           B2 => n1079, ZN => DP_OP_446J3_125_4819_n73);
   U291 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n149, A => n1079, ZN => 
                           DP_OP_446J3_125_4819_n72);
   U292 : AND2_X1 port map( A1 => C2_DATA1_4, A2 => n151, ZN => n152);
   U293 : AOI21_X1 port map( B1 => n159, B2 => OP_A_0_port, A => n152, ZN => 
                           n566);
   U294 : NOR2_X1 port map( A1 => intadd_0_SUM_0_port, A2 => n566, ZN => n565);
   U295 : INV_X1 port map( A => intadd_0_SUM_1_port, ZN => n156);
   U296 : INV_X1 port map( A => n565, ZN => n591);
   U297 : INV_X1 port map( A => n153, ZN => n154);
   U298 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_5, B1 => 
                           OP_A_0_port, B2 => n160, C1 => OP_A_1_port, C2 => 
                           n159, ZN => n592);
   U299 : OAI21_X1 port map( B1 => intadd_0_SUM_1_port, B2 => n591, A => n592, 
                           ZN => n155);
   U300 : OAI21_X1 port map( B1 => n565, B2 => n156, A => n155, ZN => 
                           intadd_1_A_0_port);
   U301 : XNOR2_X1 port map( A => DP_OP_451J3_128_3502_n15, B => n157, ZN => 
                           n158);
   U302 : OAI21_X1 port map( B1 => n1381, B2 => n158, A => n65, ZN => 
                           intadd_1_B_14_port);
   U303 : AOI222_X1 port map( A1 => OP_A_15_port, A2 => n159, B1 => n1413, B2 
                           => C430_DATA4_19, C1 => OP_A_14_port, C2 => n160, ZN
                           => intadd_1_B_13_port);
   U304 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_18, B1 => 
                           OP_A_13_port, B2 => n160, C1 => OP_A_14_port, C2 => 
                           n159, ZN => intadd_1_B_12_port);
   U305 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_17, B1 => 
                           OP_A_12_port, B2 => n160, C1 => OP_A_13_port, C2 => 
                           n159, ZN => intadd_1_B_11_port);
   U306 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_16, B1 => 
                           OP_A_12_port, B2 => n159, C1 => OP_A_11_port, C2 => 
                           n160, ZN => intadd_1_B_10_port);
   U307 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_14, B1 => n159, B2 
                           => OP_A_10_port, C1 => n160, C2 => OP_A_9_port, ZN 
                           => intadd_1_B_8_port);
   U308 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_13, B1 => n159, B2 
                           => OP_A_9_port, C1 => n160, C2 => OP_A_8_port, ZN =>
                           intadd_1_B_7_port);
   U309 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_12, B1 => n159, B2 
                           => OP_A_8_port, C1 => n160, C2 => OP_A_7_port, ZN =>
                           intadd_1_B_6_port);
   U310 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_11, B1 => n159, B2 
                           => OP_A_7_port, C1 => n160, C2 => OP_A_6_port, ZN =>
                           intadd_1_B_5_port);
   U311 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_10, B1 => n159, B2 
                           => OP_A_6_port, C1 => n160, C2 => OP_A_5_port, ZN =>
                           intadd_1_B_4_port);
   U312 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_9, B1 => n159, B2 
                           => OP_A_5_port, C1 => n160, C2 => OP_A_4_port, ZN =>
                           intadd_1_B_3_port);
   U313 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_8, B1 => n159, B2 
                           => OP_A_4_port, C1 => n160, C2 => OP_A_3_port, ZN =>
                           intadd_1_B_2_port);
   U314 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_7, B1 => n159, B2 
                           => OP_A_3_port, C1 => n160, C2 => OP_A_2_port, ZN =>
                           intadd_1_B_1_port);
   U315 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_6, B1 => 
                           OP_A_1_port, B2 => n160, C1 => n159, C2 => 
                           OP_A_2_port, ZN => intadd_1_B_0_port);
   U316 : CLKBUF_X1 port map( A => n1414, Z => n167);
   U317 : INV_X1 port map( A => n161, ZN => n162);
   U318 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_17, B1 => n61, B2 =>
                           OP_A_11_port, C1 => n1028, C2 => OP_A_10_port, ZN =>
                           intadd_2_A_9_port);
   U319 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_16, B1 => n61, B2 =>
                           OP_A_10_port, C1 => n1028, C2 => OP_A_9_port, ZN => 
                           intadd_2_A_8_port);
   U320 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_15, B1 => n61, B2 =>
                           OP_A_9_port, C1 => n1028, C2 => OP_A_8_port, ZN => 
                           intadd_2_A_7_port);
   U321 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_14, B1 => n61, B2 =>
                           OP_A_8_port, C1 => n1028, C2 => OP_A_7_port, ZN => 
                           intadd_2_A_6_port);
   U322 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_13, B1 => n61, B2 =>
                           OP_A_7_port, C1 => n1028, C2 => OP_A_6_port, ZN => 
                           intadd_2_A_5_port);
   U323 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_12, B1 => n61, B2 =>
                           OP_A_6_port, C1 => n1028, C2 => OP_A_5_port, ZN => 
                           intadd_2_A_4_port);
   U324 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_11, B1 => n61, B2 =>
                           OP_A_5_port, C1 => n1028, C2 => OP_A_4_port, ZN => 
                           intadd_2_A_3_port);
   U325 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_10, B1 => n61, B2 =>
                           OP_A_4_port, C1 => n1028, C2 => OP_A_3_port, ZN => 
                           intadd_2_A_2_port);
   U326 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_9, B1 => n61, B2 => 
                           OP_A_3_port, C1 => n1028, C2 => OP_A_2_port, ZN => 
                           intadd_2_A_1_port);
   U327 : AND2_X1 port map( A1 => C2_DATA1_6, A2 => n163, ZN => n164);
   U328 : AOI21_X1 port map( B1 => OP_A_0_port, B2 => n61, A => n164, ZN => 
                           n621);
   U329 : NOR2_X1 port map( A1 => intadd_1_SUM_0_port, A2 => n621, ZN => n620);
   U330 : INV_X1 port map( A => intadd_1_SUM_1_port, ZN => n166);
   U331 : INV_X1 port map( A => n620, ZN => n642);
   U332 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_7, B1 => n61, B2 => 
                           OP_A_1_port, C1 => n1028, C2 => OP_A_0_port, ZN => 
                           n643);
   U333 : OAI21_X1 port map( B1 => intadd_1_SUM_1_port, B2 => n642, A => n643, 
                           ZN => n165);
   U334 : OAI21_X1 port map( B1 => n620, B2 => n166, A => n165, ZN => 
                           intadd_2_A_0_port);
   U335 : AOI222_X1 port map( A1 => n167, A2 => C429_DATA4_8, B1 => n61, B2 => 
                           OP_A_2_port, C1 => n1028, C2 => OP_A_1_port, ZN => 
                           intadd_2_B_0_port);
   U336 : AOI21_X1 port map( B1 => n169, B2 => n171, A => n168, ZN => n170);
   U337 : OAI21_X1 port map( B1 => n174, B2 => n171, A => n170, ZN => N287);
   U338 : AOI21_X1 port map( B1 => n172, B2 => n1409, A => n179, ZN => n173);
   U339 : INV_X1 port map( A => n173, ZN => n175);
   U340 : OAI211_X1 port map( C1 => n176, C2 => n1408, A => n175, B => n174, ZN
                           => N288);
   U341 : INV_X1 port map( A => n177, ZN => n178);
   U342 : OAI21_X1 port map( B1 => n179, B2 => n1406, A => n178, ZN => N289);
   U343 : INV_X1 port map( A => OP2(0), ZN => n218);
   U344 : AOI22_X1 port map( A1 => OP2(0), A2 => n194, B1 => n196, B2 => n218, 
                           ZN => N247);
   U345 : INV_X1 port map( A => OP2(1), ZN => n484);
   U346 : AOI22_X1 port map( A1 => OP2(1), A2 => n194, B1 => n196, B2 => n484, 
                           ZN => N248);
   U347 : INV_X1 port map( A => OP2(2), ZN => n180);
   U348 : AOI22_X1 port map( A1 => OP2(2), A2 => n194, B1 => n196, B2 => n180, 
                           ZN => N249);
   U349 : INV_X1 port map( A => OP2(3), ZN => n181);
   U350 : AOI22_X1 port map( A1 => OP2(3), A2 => n194, B1 => n196, B2 => n181, 
                           ZN => N250);
   U351 : INV_X1 port map( A => OP2(4), ZN => n182);
   U352 : AOI22_X1 port map( A1 => OP2(4), A2 => n194, B1 => n196, B2 => n182, 
                           ZN => N251);
   U353 : INV_X1 port map( A => OP2(5), ZN => n613);
   U354 : AOI22_X1 port map( A1 => OP2(5), A2 => n194, B1 => n196, B2 => n613, 
                           ZN => N252);
   U355 : INV_X1 port map( A => OP2(6), ZN => n183);
   U356 : AOI22_X1 port map( A1 => OP2(6), A2 => n194, B1 => n196, B2 => n183, 
                           ZN => N253);
   U357 : INV_X1 port map( A => OP2(7), ZN => n665);
   U358 : AOI22_X1 port map( A1 => OP2(7), A2 => n205, B1 => n196, B2 => n665, 
                           ZN => N254);
   U359 : INV_X1 port map( A => OP2(8), ZN => n184);
   U360 : AOI22_X1 port map( A1 => OP2(8), A2 => n205, B1 => n196, B2 => n184, 
                           ZN => N255);
   U361 : INV_X1 port map( A => OP2(9), ZN => n692);
   U362 : AOI22_X1 port map( A1 => OP2(9), A2 => n205, B1 => n196, B2 => n692, 
                           ZN => N256);
   U363 : INV_X1 port map( A => OP2(10), ZN => n185);
   U364 : AOI22_X1 port map( A1 => OP2(10), A2 => n205, B1 => n196, B2 => n185,
                           ZN => N257);
   U365 : INV_X1 port map( A => OP2(11), ZN => n186);
   U366 : AOI22_X1 port map( A1 => OP2(11), A2 => n205, B1 => n196, B2 => n186,
                           ZN => N258);
   U367 : INV_X1 port map( A => OP2(12), ZN => n777);
   U368 : AOI22_X1 port map( A1 => OP2(12), A2 => n205, B1 => n196, B2 => n777,
                           ZN => N259);
   U369 : INV_X1 port map( A => OP2(13), ZN => n801);
   U370 : AOI22_X1 port map( A1 => OP2(13), A2 => n205, B1 => n196, B2 => n801,
                           ZN => N260);
   U371 : INV_X1 port map( A => OP2(14), ZN => n187);
   U372 : AOI22_X1 port map( A1 => OP2(14), A2 => n205, B1 => n196, B2 => n187,
                           ZN => N261);
   U373 : INV_X1 port map( A => OP2(15), ZN => n860);
   U374 : AOI22_X1 port map( A1 => OP2(15), A2 => n205, B1 => n196, B2 => n860,
                           ZN => N262);
   U375 : INV_X1 port map( A => OP2(16), ZN => n188);
   U376 : AOI22_X1 port map( A1 => OP2(16), A2 => n205, B1 => n196, B2 => n188,
                           ZN => N263);
   U377 : INV_X1 port map( A => OP2(17), ZN => n189);
   U378 : AOI22_X1 port map( A1 => OP2(17), A2 => n194, B1 => n196, B2 => n189,
                           ZN => N264);
   U379 : INV_X1 port map( A => OP2(18), ZN => n190);
   U380 : AOI22_X1 port map( A1 => OP2(18), A2 => n194, B1 => n196, B2 => n190,
                           ZN => N265);
   U381 : INV_X1 port map( A => OP2(19), ZN => n191);
   U382 : AOI22_X1 port map( A1 => OP2(19), A2 => n194, B1 => n196, B2 => n191,
                           ZN => N266);
   U383 : INV_X1 port map( A => OP2(20), ZN => n192);
   U384 : AOI22_X1 port map( A1 => OP2(20), A2 => n194, B1 => n196, B2 => n192,
                           ZN => N267);
   U385 : INV_X1 port map( A => OP2(21), ZN => n193);
   U386 : AOI22_X1 port map( A1 => OP2(21), A2 => n194, B1 => n196, B2 => n193,
                           ZN => N268);
   U387 : INV_X1 port map( A => OP2(22), ZN => n195);
   U388 : AOI22_X1 port map( A1 => OP2(22), A2 => n205, B1 => n196, B2 => n195,
                           ZN => N269);
   U389 : INV_X1 port map( A => OP2(23), ZN => n197);
   U390 : AOI22_X1 port map( A1 => OP2(23), A2 => n205, B1 => n196, B2 => n197,
                           ZN => N270);
   U391 : INV_X1 port map( A => OP2(24), ZN => n1138);
   U392 : AOI22_X1 port map( A1 => OP2(24), A2 => n205, B1 => n196, B2 => n1138
                           , ZN => N271);
   U393 : INV_X1 port map( A => OP2(25), ZN => n198);
   U394 : AOI22_X1 port map( A1 => OP2(25), A2 => n205, B1 => n196, B2 => n198,
                           ZN => N272);
   U395 : INV_X1 port map( A => OP2(26), ZN => n199);
   U396 : AOI22_X1 port map( A1 => OP2(26), A2 => n205, B1 => n196, B2 => n199,
                           ZN => N273);
   U397 : INV_X1 port map( A => OP2(27), ZN => n200);
   U398 : AOI22_X1 port map( A1 => OP2(27), A2 => n205, B1 => n196, B2 => n200,
                           ZN => N274);
   U399 : INV_X1 port map( A => OP2(28), ZN => n201);
   U400 : AOI22_X1 port map( A1 => OP2(28), A2 => n205, B1 => n196, B2 => n201,
                           ZN => N275);
   U401 : INV_X1 port map( A => OP2(29), ZN => n202);
   U402 : AOI22_X1 port map( A1 => OP2(29), A2 => n205, B1 => n196, B2 => n202,
                           ZN => N276);
   U403 : INV_X1 port map( A => OP2(30), ZN => n203);
   U404 : AOI22_X1 port map( A1 => OP2(30), A2 => n205, B1 => n196, B2 => n203,
                           ZN => N277);
   U405 : INV_X1 port map( A => OP2(31), ZN => n204);
   U406 : AOI22_X1 port map( A1 => OP2(31), A2 => n205, B1 => n196, B2 => n204,
                           ZN => N278);
   U407 : INV_X1 port map( A => N284, ZN => n1159);
   U408 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => n55, ZN => n1204);
   U409 : NAND2_X1 port map( A1 => n543, A2 => OP_A_21_port, ZN => n1059);
   U410 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => n604, ZN => n1133);
   U411 : OR2_X1 port map( A1 => OP_B_1_port, A2 => OP_B_0_port, ZN => n608);
   U412 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => n56, ZN => n1003);
   U413 : AND4_X1 port map( A1 => n1204, A2 => n1059, A3 => n1133, A4 => n1003,
                           ZN => n785);
   U414 : NAND2_X1 port map( A1 => n492, A2 => OP_A_25_port, ZN => n1205);
   U415 : NAND2_X1 port map( A1 => OP_A_27_port, A2 => n55, ZN => n1318);
   U416 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => n56, ZN => n1130);
   U417 : CLKBUF_X1 port map( A => n604, Z => n554);
   U418 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => n554, ZN => n1272);
   U419 : NAND4_X1 port map( A1 => n1205, A2 => n1318, A3 => n1130, A4 => n1272
                           , ZN => n782);
   U420 : INV_X1 port map( A => n858, ZN => n511);
   U421 : INV_X1 port map( A => OP_A_31_port, ZN => n1370);
   U422 : AOI22_X1 port map( A1 => OP_A_30_port, A2 => n604, B1 => OP_A_28_port
                           , B2 => n56, ZN => n206);
   U423 : NAND2_X1 port map( A1 => n492, A2 => OP_A_29_port, ZN => n1319);
   U424 : OAI211_X1 port map( C1 => n578, C2 => n1370, A => n206, B => n1319, 
                           ZN => n1265);
   U425 : AOI22_X1 port map( A1 => n856, A2 => n782, B1 => n511, B2 => n1265, 
                           ZN => n208);
   U426 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => n55, ZN => n1058);
   U427 : NAND2_X1 port map( A1 => n492, A2 => OP_A_17_port, ZN => n938);
   U428 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => n554, ZN => n1006);
   U429 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n56, ZN => n888);
   U430 : NAND4_X1 port map( A1 => n1058, A2 => n938, A3 => n1006, A4 => n888, 
                           ZN => n778);
   U431 : NAND2_X1 port map( A1 => n895, A2 => n778, ZN => n207);
   U432 : OAI211_X1 port map( C1 => n785, C2 => n743, A => n208, B => n207, ZN 
                           => n899);
   U433 : NAND2_X1 port map( A1 => OP_A_15_port, A2 => n55, ZN => n937);
   U434 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => n56, ZN => n768);
   U435 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => n554, ZN => n890);
   U436 : AND4_X1 port map( A1 => n820, A2 => n937, A3 => n768, A4 => n890, ZN 
                           => n772);
   U437 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n858, ZN => n1352);
   U438 : INV_X1 port map( A => n1352, ZN => n892);
   U439 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => n55, ZN => n818);
   U440 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => n554, ZN => n769);
   U441 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => n56, ZN => n673);
   U442 : AND4_X1 port map( A1 => n818, A2 => n727, A3 => n769, A4 => n673, ZN 
                           => n682);
   U443 : INV_X1 port map( A => n856, ZN => n742);
   U444 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n742, ZN => n1350);
   U445 : INV_X1 port map( A => n1350, ZN => n567);
   U446 : OAI22_X1 port map( A1 => n772, A2 => n892, B1 => n682, B2 => n567, ZN
                           => n214);
   U447 : NAND2_X1 port map( A1 => OP_A_3_port, A2 => n55, ZN => n627);
   U448 : NAND2_X1 port map( A1 => n492, A2 => OP_A_1_port, ZN => n508);
   U449 : NAND2_X1 port map( A1 => OP_A_0_port, A2 => n56, ZN => n896);
   U450 : NAND2_X1 port map( A1 => OP_A_2_port, A2 => n554, ZN => n209);
   U451 : AND4_X1 port map( A1 => n627, A2 => n508, A3 => n896, A4 => n209, ZN 
                           => n212);
   U452 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n766, ZN => n1360);
   U453 : INV_X1 port map( A => n1360, ZN => n1261);
   U454 : NAND2_X1 port map( A1 => OP_A_7_port, A2 => n55, ZN => n726);
   U455 : NAND2_X1 port map( A1 => OP_A_4_port, A2 => n56, ZN => n210);
   U456 : NAND2_X1 port map( A1 => OP_A_6_port, A2 => n554, ZN => n675);
   U457 : NAND4_X1 port map( A1 => n726, A2 => n629, A3 => n210, A4 => n675, ZN
                           => n583);
   U458 : INV_X1 port map( A => n583, ZN => n211);
   U459 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n743, ZN => n1358);
   U460 : INV_X1 port map( A => n1358, ZN => n900);
   U461 : OAI22_X1 port map( A1 => n212, A2 => n1261, B1 => n211, B2 => n900, 
                           ZN => n213);
   U462 : AOI211_X1 port map( C1 => OP_B_4_port, C2 => n899, A => n214, B => 
                           n213, ZN => n482);
   U463 : NOR2_X1 port map( A1 => n216, A2 => n215, ZN => n1347);
   U464 : CLKBUF_X1 port map( A => n1347, Z => n1330);
   U465 : NAND2_X1 port map( A1 => OP_B_0_port, A2 => OP_A_0_port, ZN => n293);
   U466 : OR2_X1 port map( A1 => n217, A2 => n1411, ZN => n1139);
   U467 : OAI22_X1 port map( A1 => n1396, A2 => n293, B1 => n1139, B2 => n218, 
                           ZN => n221);
   U468 : NOR2_X1 port map( A1 => n219, A2 => OP_LOGIC_0_port, ZN => n475);
   U469 : INV_X1 port map( A => OP_LOGIC_1_port, ZN => n222);
   U470 : AND2_X1 port map( A1 => n475, A2 => n222, ZN => n1245);
   U471 : INV_X1 port map( A => n1228, ZN => n1062);
   U472 : OAI22_X1 port map( A1 => n293, A2 => n1369, B1 => n896, B2 => n1062, 
                           ZN => n220);
   U473 : AOI211_X1 port map( C1 => n1330, C2 => OP1(0), A => n221, B => n220, 
                           ZN => n481);
   U474 : NAND3_X1 port map( A1 => N281, A2 => n222, A3 => OP_LOGIC_0_port, ZN 
                           => n1368);
   U475 : INV_X1 port map( A => OP_A_0_port, ZN => n550);
   U476 : NAND2_X1 port map( A1 => n223, A2 => n550, ZN => n488);
   U477 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n551, ZN => n365);
   U478 : INV_X1 port map( A => n365, ZN => n316);
   U479 : INV_X1 port map( A => OP_A_5_port, ZN => n607);
   U480 : NAND2_X1 port map( A1 => n607, A2 => OP_B_5_port, ZN => n369);
   U481 : OAI21_X1 port map( B1 => n1363, B2 => OP_A_4_port, A => n369, ZN => 
                           n320);
   U482 : INV_X1 port map( A => OP_A_1_port, ZN => n579);
   U483 : OAI21_X1 port map( B1 => n224, B2 => OP_A_1_port, A => OP_A_0_port, 
                           ZN => n315);
   U484 : OAI211_X1 port map( C1 => n579, C2 => n55, A => n608, B => n315, ZN 
                           => n366);
   U485 : NOR2_X1 port map( A1 => OP_A_3_port, A2 => n1160, ZN => n302);
   U486 : AOI21_X1 port map( B1 => n577, B2 => OP_B_2_port, A => n302, ZN => 
                           n364);
   U487 : INV_X1 port map( A => n302, ZN => n317);
   U488 : NOR2_X1 port map( A1 => n577, A2 => OP_B_2_port, ZN => n225);
   U489 : AOI22_X1 port map( A1 => n366, A2 => n364, B1 => n317, B2 => n225, ZN
                           => n227);
   U490 : INV_X1 port map( A => OP_A_4_port, ZN => n368);
   U491 : NOR2_X1 port map( A1 => n368, A2 => OP_B_4_port, ZN => n226);
   U492 : NOR2_X1 port map( A1 => n607, A2 => OP_B_5_port, ZN => n371);
   U493 : AOI21_X1 port map( B1 => n369, B2 => n226, A => n371, ZN => n319);
   U494 : OAI221_X1 port map( B1 => n316, B2 => n320, C1 => n227, C2 => n320, A
                           => n319, ZN => n233);
   U495 : NAND2_X1 port map( A1 => n378, A2 => OP_A_6_port, ZN => n228);
   U496 : NOR2_X1 port map( A1 => n295, A2 => OP_A_7_port, ZN => n379);
   U497 : NAND2_X1 port map( A1 => n295, A2 => OP_A_7_port, ZN => n380);
   U498 : OAI21_X1 port map( B1 => n228, B2 => n379, A => n380, ZN => n322);
   U499 : INV_X1 port map( A => OP_A_6_port, ZN => n372);
   U500 : AOI21_X1 port map( B1 => n372, B2 => OP_B_6_port, A => n379, ZN => 
                           n324);
   U501 : INV_X1 port map( A => OP_A_12_port, ZN => n234);
   U502 : NAND2_X1 port map( A1 => n234, A2 => OP_B_12_port, ZN => n333);
   U503 : INV_X1 port map( A => OP_A_13_port, ZN => n235);
   U504 : INV_X1 port map( A => OP_B_14_port, ZN => n229);
   U505 : NAND2_X1 port map( A1 => n1081, A2 => OP_B_15_port, ZN => n349);
   U506 : OAI21_X1 port map( B1 => n229, B2 => OP_A_14_port, A => n349, ZN => 
                           n230);
   U507 : AOI21_X1 port map( B1 => n235, B2 => OP_B_13_port, A => n230, ZN => 
                           n241);
   U508 : AND2_X1 port map( A1 => n333, A2 => n241, ZN => n231);
   U509 : INV_X1 port map( A => OP_A_10_port, ZN => n336);
   U510 : INV_X1 port map( A => OP_A_11_port, ZN => n236);
   U511 : NAND2_X1 port map( A1 => n236, A2 => OP_B_11_port, ZN => n343);
   U512 : INV_X1 port map( A => n343, ZN => n240);
   U513 : AOI21_X1 port map( B1 => OP_B_10_port, B2 => n336, A => n240, ZN => 
                           n238);
   U514 : INV_X1 port map( A => OP_A_9_port, ZN => n303);
   U515 : INV_X1 port map( A => OP_A_8_port, ZN => n237);
   U516 : AOI22_X1 port map( A1 => OP_B_9_port, A2 => n303, B1 => OP_B_8_port, 
                           B2 => n237, ZN => n339);
   U517 : NAND3_X1 port map( A1 => n231, A2 => n238, A3 => n339, ZN => n326);
   U518 : INV_X1 port map( A => n326, ZN => n232);
   U519 : OAI221_X1 port map( B1 => n233, B2 => n322, C1 => n324, C2 => n322, A
                           => n232, ZN => n249_port);
   U520 : INV_X1 port map( A => OP_A_14_port, ZN => n332);
   U521 : NOR2_X1 port map( A1 => n332, A2 => OP_B_14_port, ZN => n346);
   U522 : OAI22_X1 port map( A1 => OP_B_13_port, A2 => n235, B1 => OP_B_12_port
                           , B2 => n234, ZN => n335);
   U523 : OR2_X1 port map( A1 => n336, A2 => OP_B_10_port, ZN => n337);
   U524 : NOR2_X1 port map( A1 => n236, A2 => OP_B_11_port, ZN => n345);
   U525 : INV_X1 port map( A => n345, ZN => n338);
   U526 : INV_X1 port map( A => OP_B_9_port, ZN => n340);
   U527 : OAI22_X1 port map( A1 => OP_B_8_port, A2 => n237, B1 => OP_B_9_port, 
                           B2 => n303, ZN => n357);
   U528 : OAI211_X1 port map( C1 => OP_A_9_port, C2 => n340, A => n238, B => 
                           n357, ZN => n239);
   U529 : OAI211_X1 port map( C1 => n240, C2 => n337, A => n338, B => n239, ZN 
                           => n242);
   U530 : OAI221_X1 port map( B1 => n335, B2 => n333, C1 => n335, C2 => n242, A
                           => n241, ZN => n243);
   U531 : INV_X1 port map( A => n243, ZN => n244);
   U532 : NOR2_X1 port map( A1 => n1081, A2 => OP_B_15_port, ZN => n352);
   U533 : AOI211_X1 port map( C1 => n349, C2 => n346, A => n244, B => n352, ZN 
                           => n327);
   U534 : INV_X1 port map( A => OP_B_17_port, ZN => n256_port);
   U535 : NOR2_X1 port map( A1 => OP_A_17_port, A2 => n256_port, ZN => n394);
   U536 : INV_X1 port map( A => OP_B_16_port, ZN => n257_port);
   U537 : NOR2_X1 port map( A1 => OP_A_16_port, A2 => n257_port, ZN => n395);
   U538 : INV_X1 port map( A => OP_B_18_port, ZN => n358);
   U539 : INV_X1 port map( A => OP_A_19_port, ZN => n255_port);
   U540 : NAND2_X1 port map( A1 => OP_B_19_port, A2 => n255_port, ZN => n397);
   U541 : OAI21_X1 port map( B1 => OP_A_18_port, B2 => n358, A => n397, ZN => 
                           n258_port);
   U542 : INV_X1 port map( A => OP_A_21_port, ZN => n246_port);
   U543 : INV_X1 port map( A => OP_B_22_port, ZN => n390);
   U544 : INV_X1 port map( A => OP_A_23_port, ZN => n253_port);
   U545 : NAND2_X1 port map( A1 => OP_B_23_port, A2 => n253_port, ZN => n408);
   U546 : OAI21_X1 port map( B1 => OP_A_22_port, B2 => n390, A => n408, ZN => 
                           n245);
   U547 : AOI21_X1 port map( B1 => OP_B_21_port, B2 => n246_port, A => n245, ZN
                           => n247_port);
   U548 : INV_X1 port map( A => n247_port, ZN => n261_port);
   U549 : INV_X1 port map( A => OP_B_20_port, ZN => n254_port);
   U550 : NOR2_X1 port map( A1 => n254_port, A2 => OP_A_20_port, ZN => n400);
   U551 : OR2_X1 port map( A1 => n261_port, A2 => n400, ZN => n248_port);
   U552 : OR4_X1 port map( A1 => n394, A2 => n395, A3 => n258_port, A4 => 
                           n248_port, ZN => n325);
   U553 : AOI21_X1 port map( B1 => n249_port, B2 => n327, A => n325, ZN => 
                           n250_port);
   U554 : INV_X1 port map( A => n250_port, ZN => n285_port);
   U555 : INV_X1 port map( A => OP_B_24_port, ZN => n417);
   U556 : INV_X1 port map( A => OP_A_25_port, ZN => n266_port);
   U557 : NAND2_X1 port map( A1 => n266_port, A2 => OP_B_25_port, ZN => n418);
   U558 : INV_X1 port map( A => OP_A_26_port, ZN => n423);
   U559 : INV_X1 port map( A => OP_A_27_port, ZN => n1248);
   U560 : NAND2_X1 port map( A1 => OP_B_27_port, A2 => n1248, ZN => n425);
   U561 : INV_X1 port map( A => n425, ZN => n271_port);
   U562 : AOI21_X1 port map( B1 => n423, B2 => OP_B_26_port, A => n271_port, ZN
                           => n267_port);
   U563 : OAI211_X1 port map( C1 => n417, C2 => OP_A_24_port, A => n418, B => 
                           n267_port, ZN => n277_port);
   U564 : INV_X1 port map( A => OP_B_28_port, ZN => n275_port);
   U565 : INV_X1 port map( A => OP_A_29_port, ZN => n1297);
   U566 : NAND2_X1 port map( A1 => n1297, A2 => OP_B_29_port, ZN => n413);
   U567 : NOR2_X1 port map( A1 => OP_B_31_port, A2 => n1370, ZN => n428);
   U568 : INV_X1 port map( A => OP_A_30_port, ZN => n252_port);
   U569 : NAND2_X1 port map( A1 => OP_B_30_port, A2 => n252_port, ZN => n452);
   U570 : INV_X1 port map( A => n452, ZN => n411);
   U571 : NOR2_X1 port map( A1 => n428, A2 => n411, ZN => n272_port);
   U572 : OAI211_X1 port map( C1 => n275_port, C2 => OP_A_28_port, A => n413, B
                           => n272_port, ZN => n251_port);
   U573 : OR2_X1 port map( A1 => n277_port, A2 => n251_port, ZN => n463);
   U574 : NOR2_X1 port map( A1 => OP_B_30_port, A2 => n252_port, ZN => n440);
   U575 : INV_X1 port map( A => n428, ZN => n450);
   U576 : NAND2_X1 port map( A1 => n1370, A2 => OP_B_31_port, ZN => n306);
   U577 : INV_X1 port map( A => n306, ZN => n453);
   U578 : AND2_X1 port map( A1 => n390, A2 => OP_A_22_port, ZN => n264_port);
   U579 : NOR2_X1 port map( A1 => OP_B_23_port, A2 => n253_port, ZN => n409);
   U580 : INV_X1 port map( A => OP_B_21_port, ZN => n402);
   U581 : AOI22_X1 port map( A1 => OP_A_21_port, A2 => n402, B1 => OP_A_20_port
                           , B2 => n254_port, ZN => n404);
   U582 : INV_X1 port map( A => OP_A_18_port, ZN => n391);
   U583 : NOR2_X1 port map( A1 => OP_B_18_port, A2 => n391, ZN => n260_port);
   U584 : NOR2_X1 port map( A1 => OP_B_19_port, A2 => n255_port, ZN => n398);
   U585 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n256_port, ZN => n393);
   U586 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n257_port, ZN => n360);
   U587 : AOI211_X1 port map( C1 => n393, C2 => n360, A => n394, B => n258_port
                           , ZN => n259_port);
   U588 : AOI211_X1 port map( C1 => n260_port, C2 => n397, A => n398, B => 
                           n259_port, ZN => n262_port);
   U589 : AOI221_X1 port map( B1 => n400, B2 => n404, C1 => n262_port, C2 => 
                           n404, A => n261_port, ZN => n263_port);
   U590 : AOI211_X1 port map( C1 => n264_port, C2 => n408, A => n409, B => 
                           n263_port, ZN => n283_port);
   U591 : INV_X1 port map( A => n413, ZN => n289_port);
   U592 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n275_port, ZN => 
                           n265_port);
   U593 : NOR2_X1 port map( A1 => OP_B_29_port, A2 => n1297, ZN => n415);
   U594 : INV_X1 port map( A => n415, ZN => n362);
   U595 : OAI21_X1 port map( B1 => n289_port, B2 => n265_port, A => n362, ZN =>
                           n281_port);
   U596 : INV_X1 port map( A => OP_A_28_port, ZN => n412);
   U597 : AOI21_X1 port map( B1 => OP_B_28_port, B2 => n412, A => n289_port, ZN
                           => n280_port);
   U598 : OR2_X1 port map( A1 => n423, A2 => OP_B_26_port, ZN => n270_port);
   U599 : NOR2_X1 port map( A1 => OP_B_25_port, A2 => n266_port, ZN => n419);
   U600 : AND2_X1 port map( A1 => n417, A2 => OP_A_24_port, ZN => n268_port);
   U601 : OAI211_X1 port map( C1 => n419, C2 => n268_port, A => n418, B => 
                           n267_port, ZN => n269_port);
   U602 : OR2_X1 port map( A1 => n1248, A2 => OP_B_27_port, ZN => n422);
   U603 : OAI211_X1 port map( C1 => n271_port, C2 => n270_port, A => n269_port,
                           B => n422, ZN => n279_port);
   U604 : OAI221_X1 port map( B1 => n281_port, B2 => n280_port, C1 => n281_port
                           , C2 => n279_port, A => n272_port, ZN => n273_port);
   U605 : OAI21_X1 port map( B1 => n283_port, B2 => n463, A => n273_port, ZN =>
                           n274_port);
   U606 : AOI211_X1 port map( C1 => n440, C2 => n450, A => n453, B => n274_port
                           , ZN => n461);
   U607 : OAI21_X1 port map( B1 => n285_port, B2 => n463, A => n461, ZN => 
                           n287_port);
   U608 : NOR2_X1 port map( A1 => OP_COMPARE_1_port, A2 => OP_COMPARE_2_port, 
                           ZN => n438);
   U609 : NOR2_X1 port map( A1 => n453, A2 => n411, ZN => n278_port);
   U610 : OAI211_X1 port map( C1 => n275_port, C2 => OP_A_28_port, A => n413, B
                           => n278_port, ZN => n276_port);
   U611 : OR2_X1 port map( A1 => n277_port, A2 => n276_port, ZN => n330);
   U612 : OAI221_X1 port map( B1 => n281_port, B2 => n280_port, C1 => n281_port
                           , C2 => n279_port, A => n278_port, ZN => n282_port);
   U613 : OAI21_X1 port map( B1 => n283_port, B2 => n330, A => n282_port, ZN =>
                           n284_port);
   U614 : AOI211_X1 port map( C1 => n440, C2 => n306, A => n428, B => n284_port
                           , ZN => n329);
   U615 : OAI211_X1 port map( C1 => n330, C2 => n285_port, A => 
                           OP_COMPARE_0_port, B => n329, ZN => n286_port);
   U616 : OAI211_X1 port map( C1 => OP_COMPARE_0_port, C2 => n287_port, A => 
                           n438, B => n286_port, ZN => n474);
   U617 : INV_X1 port map( A => OP_COMPARE_3_port, ZN => n473);
   U618 : NAND2_X1 port map( A1 => n425, A2 => n422, ZN => n1241);
   U619 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => OP_B_19_port, ZN => n976
                           );
   U620 : OR2_X1 port map( A1 => OP_A_19_port, A2 => OP_B_19_port, ZN => n992);
   U621 : NAND2_X1 port map( A1 => n976, A2 => n992, ZN => n975);
   U622 : INV_X1 port map( A => n975, ZN => n984);
   U623 : NOR2_X1 port map( A1 => OP_A_23_port, A2 => OP_B_23_port, ZN => n1108
                           );
   U624 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => OP_B_23_port, ZN => 
                           n1123);
   U625 : INV_X1 port map( A => n1123, ZN => n288_port);
   U626 : NOR2_X1 port map( A1 => n1108, A2 => n288_port, ZN => n1106);
   U627 : AND2_X1 port map( A1 => OP_A_15_port, A2 => OP_B_15_port, ZN => n878)
                           ;
   U628 : NOR2_X1 port map( A1 => OP_A_15_port, A2 => OP_B_15_port, ZN => n863)
                           ;
   U629 : NOR2_X1 port map( A1 => n878, A2 => n863, ZN => n874);
   U630 : OR4_X1 port map( A1 => n1241, A2 => n984, A3 => n1106, A4 => n874, ZN
                           => n301);
   U631 : NOR2_X1 port map( A1 => n289_port, A2 => n415, ZN => n1302);
   U632 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => OP_B_26_port, ZN => 
                           n1237);
   U633 : OAI21_X1 port map( B1 => OP_A_26_port, B2 => OP_B_26_port, A => n1237
                           , ZN => n1200);
   U634 : NOR2_X1 port map( A1 => OP_A_30_port, A2 => OP_B_30_port, ZN => n1375
                           );
   U635 : NAND2_X1 port map( A1 => OP_A_30_port, A2 => OP_B_30_port, ZN => 
                           n1377);
   U636 : INV_X1 port map( A => n1377, ZN => n290);
   U637 : NOR2_X1 port map( A1 => n1375, A2 => n290, ZN => n1343);
   U638 : INV_X1 port map( A => n1343, ZN => n1333);
   U639 : NOR2_X1 port map( A1 => OP_A_28_port, A2 => OP_B_28_port, ZN => n1299
                           );
   U640 : INV_X1 port map( A => n1299, ZN => n291);
   U641 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => OP_B_28_port, ZN => 
                           n1301);
   U642 : NAND2_X1 port map( A1 => n291, A2 => n1301, ZN => n1267);
   U643 : NAND4_X1 port map( A1 => n1302, A2 => n1200, A3 => n1333, A4 => n1267
                           , ZN => n300);
   U644 : NAND2_X1 port map( A1 => n1363, A2 => n368, ZN => n598);
   U645 : NAND2_X1 port map( A1 => OP_B_4_port, A2 => OP_A_4_port, ZN => n571);
   U646 : NAND2_X1 port map( A1 => n598, A2 => n571, ZN => n574);
   U647 : NAND2_X1 port map( A1 => n582, A2 => n577, ZN => n547);
   U648 : NOR2_X1 port map( A1 => n582, A2 => n577, ZN => n507);
   U649 : INV_X1 port map( A => n507, ZN => n292);
   U650 : NAND2_X1 port map( A1 => n547, A2 => n292, ZN => n524);
   U651 : NOR2_X1 port map( A1 => OP_B_1_port, A2 => OP_A_1_port, ZN => n521);
   U652 : INV_X1 port map( A => n521, ZN => n503);
   U653 : NAND2_X1 port map( A1 => OP_B_1_port, A2 => OP_A_1_port, ZN => n520);
   U654 : NAND2_X1 port map( A1 => n503, A2 => n520, ZN => n506);
   U655 : NAND2_X1 port map( A1 => n293, A2 => n488, ZN => n476);
   U656 : NAND4_X1 port map( A1 => n574, A2 => n524, A3 => n506, A4 => n476, ZN
                           => n299);
   U657 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => OP_B_11_port, ZN => n750
                           );
   U658 : OR2_X1 port map( A1 => OP_A_11_port, A2 => OP_B_11_port, ZN => n774);
   U659 : NAND2_X1 port map( A1 => n750, A2 => n774, ZN => n755);
   U660 : NAND2_X1 port map( A1 => OP_B_7_port, A2 => OP_A_7_port, ZN => n646);
   U661 : INV_X1 port map( A => OP_A_7_port, ZN => n294);
   U662 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => n679);
   U663 : NAND2_X1 port map( A1 => n646, A2 => n679, ZN => n654);
   U664 : NAND2_X1 port map( A1 => OP_B_6_port, A2 => OP_A_6_port, ZN => n650);
   U665 : NOR2_X1 port map( A1 => OP_B_6_port, A2 => OP_A_6_port, ZN => n652);
   U666 : INV_X1 port map( A => n652, ZN => n296);
   U667 : NAND2_X1 port map( A1 => n650, A2 => n296, ZN => n637);
   U668 : NAND2_X1 port map( A1 => OP_B_5_port, A2 => OP_A_5_port, ZN => n594);
   U669 : NAND2_X1 port map( A1 => n297, A2 => n607, ZN => n633);
   U670 : NAND2_X1 port map( A1 => n594, A2 => n633, ZN => n601);
   U671 : NAND4_X1 port map( A1 => n755, A2 => n654, A3 => n637, A4 => n601, ZN
                           => n298);
   U672 : NOR4_X1 port map( A1 => n301, A2 => n300, A3 => n299, A4 => n298, ZN 
                           => n314);
   U673 : NOR2_X1 port map( A1 => n365, A2 => n302, ZN => n558);
   U674 : NOR2_X1 port map( A1 => OP_A_13_port, A2 => OP_B_13_port, ZN => n832)
                           ;
   U675 : INV_X1 port map( A => n832, ZN => n794);
   U676 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => OP_B_13_port, ZN => n830
                           );
   U677 : NAND2_X1 port map( A1 => n794, A2 => n830, ZN => n799);
   U678 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => OP_B_8_port, ZN => n712);
   U679 : NOR2_X1 port map( A1 => OP_A_8_port, A2 => OP_B_8_port, ZN => n716);
   U680 : INV_X1 port map( A => n716, ZN => n672);
   U681 : NAND2_X1 port map( A1 => n712, A2 => n672, ZN => n681);
   U682 : NOR2_X1 port map( A1 => OP_A_9_port, A2 => OP_B_9_port, ZN => n715);
   U683 : NOR2_X1 port map( A1 => n303, A2 => n340, ZN => n699);
   U684 : NOR2_X1 port map( A1 => n715, A2 => n699, ZN => n703);
   U685 : INV_X1 port map( A => n703, ZN => n304);
   U686 : NAND4_X1 port map( A1 => n558, A2 => n799, A3 => n681, A4 => n304, ZN
                           => n312);
   U687 : NOR2_X1 port map( A1 => OP_A_21_port, A2 => OP_B_21_port, ZN => n1051
                           );
   U688 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => OP_B_21_port, ZN => 
                           n1049);
   U689 : INV_X1 port map( A => n1049, ZN => n1022);
   U690 : NOR2_X1 port map( A1 => n1051, A2 => n1022, ZN => n1021);
   U691 : NOR2_X1 port map( A1 => OP_A_25_port, A2 => OP_B_25_port, ZN => n1196
                           );
   U692 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => OP_B_25_port, ZN => 
                           n1194);
   U693 : INV_X1 port map( A => n1194, ZN => n305);
   U694 : NOR2_X1 port map( A1 => n1196, A2 => n305, ZN => n1165);
   U695 : NOR2_X1 port map( A1 => OP_A_17_port, A2 => OP_B_17_port, ZN => n954)
                           ;
   U696 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => OP_B_17_port, ZN => n952
                           );
   U697 : INV_X1 port map( A => n952, ZN => n929);
   U698 : NOR2_X1 port map( A1 => n954, A2 => n929, ZN => n919);
   U699 : NAND2_X1 port map( A1 => n306, A2 => n450, ZN => n1371);
   U700 : OR4_X1 port map( A1 => n1021, A2 => n1165, A3 => n919, A4 => n1371, 
                           ZN => n311);
   U701 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => OP_B_18_port, ZN => n981
                           );
   U702 : INV_X1 port map( A => n981, ZN => n949);
   U703 : NOR2_X1 port map( A1 => OP_A_18_port, A2 => OP_B_18_port, ZN => n983)
                           ;
   U704 : NOR2_X1 port map( A1 => n949, A2 => n983, ZN => n959);
   U705 : INV_X1 port map( A => n959, ZN => n307);
   U706 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => OP_B_20_port, ZN => 
                           n1047);
   U707 : NOR2_X1 port map( A1 => OP_A_20_port, A2 => OP_B_20_port, ZN => n1050
                           );
   U708 : INV_X1 port map( A => n1050, ZN => n1008);
   U709 : NAND2_X1 port map( A1 => n1047, A2 => n1008, ZN => n1019);
   U710 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => OP_B_22_port, ZN => 
                           n1124);
   U711 : OAI21_X1 port map( B1 => OP_A_22_port, B2 => OP_B_22_port, A => n1124
                           , ZN => n1125);
   U712 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => OP_B_24_port, ZN => 
                           n1193);
   U713 : NOR2_X1 port map( A1 => OP_A_24_port, A2 => OP_B_24_port, ZN => n1195
                           );
   U714 : INV_X1 port map( A => n1195, ZN => n1142);
   U715 : NAND2_X1 port map( A1 => n1193, A2 => n1142, ZN => n1129);
   U716 : NAND4_X1 port map( A1 => n307, A2 => n1019, A3 => n1125, A4 => n1129,
                           ZN => n310);
   U717 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => OP_B_10_port, ZN => n756
                           );
   U718 : OAI21_X1 port map( B1 => OP_A_10_port, B2 => OP_B_10_port, A => n756,
                           ZN => n720);
   U719 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => OP_B_12_port, ZN => n828
                           );
   U720 : NOR2_X1 port map( A1 => OP_A_12_port, A2 => OP_B_12_port, ZN => n831)
                           ;
   U721 : INV_X1 port map( A => n831, ZN => n781);
   U722 : NAND2_X1 port map( A1 => n828, A2 => n781, ZN => n780);
   U723 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => OP_B_14_port, ZN => n871
                           );
   U724 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => OP_B_14_port, A => n871,
                           ZN => n836);
   U725 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => OP_B_16_port, ZN => n950
                           );
   U726 : NOR2_X1 port map( A1 => OP_A_16_port, A2 => OP_B_16_port, ZN => n953)
                           ;
   U727 : INV_X1 port map( A => n953, ZN => n308);
   U728 : NAND2_X1 port map( A1 => n950, A2 => n308, ZN => n905);
   U729 : NAND4_X1 port map( A1 => n720, A2 => n780, A3 => n836, A4 => n905, ZN
                           => n309);
   U730 : NOR4_X1 port map( A1 => n312, A2 => n311, A3 => n310, A4 => n309, ZN 
                           => n313);
   U731 : AOI211_X1 port map( C1 => n314, C2 => n313, A => OP_COMPARE_1_port, B
                           => OP_COMPARE_2_port, ZN => n470);
   U732 : OAI22_X1 port map( A1 => OP_B_0_port, A2 => n315, B1 => OP_B_1_port, 
                           B2 => n579, ZN => n318);
   U733 : OAI21_X1 port map( B1 => OP_B_2_port, B2 => n577, A => n316, ZN => 
                           n367);
   U734 : AOI22_X1 port map( A1 => n364, A2 => n318, B1 => n317, B2 => n367, ZN
                           => n321);
   U735 : OAI21_X1 port map( B1 => n321, B2 => n320, A => n319, ZN => n323);
   U736 : AOI21_X1 port map( B1 => n324, B2 => n323, A => n322, ZN => n361);
   U737 : AOI221_X1 port map( B1 => n361, B2 => n327, C1 => n326, C2 => n327, A
                           => n325, ZN => n328);
   U738 : INV_X1 port map( A => n328, ZN => n462);
   U739 : INV_X1 port map( A => OP_COMPARE_1_port, ZN => n460);
   U740 : OAI211_X1 port map( C1 => n330, C2 => n462, A => n460, B => n329, ZN 
                           => n331);
   U741 : INV_X1 port map( A => n331, ZN => n437);
   U742 : NAND2_X1 port map( A1 => OP_B_14_port, A2 => n332, ZN => n351);
   U743 : INV_X1 port map( A => OP_B_13_port, ZN => n334);
   U744 : AOI222_X1 port map( A1 => OP_A_13_port, A2 => n334, B1 => 
                           OP_A_13_port, B2 => n333, C1 => n334, C2 => n333, ZN
                           => n348);
   U745 : INV_X1 port map( A => n335, ZN => n354);
   U746 : NAND2_X1 port map( A1 => OP_B_10_port, A2 => n336, ZN => n344);
   U747 : NAND2_X1 port map( A1 => n338, A2 => n337, ZN => n355);
   U748 : AOI211_X1 port map( C1 => n340, C2 => OP_A_9_port, A => n355, B => 
                           n339, ZN => n341);
   U749 : INV_X1 port map( A => n341, ZN => n342);
   U750 : OAI211_X1 port map( C1 => n345, C2 => n344, A => n343, B => n342, ZN 
                           => n347);
   U751 : NOR2_X1 port map( A1 => n352, A2 => n346, ZN => n353);
   U752 : OAI221_X1 port map( B1 => n348, B2 => n354, C1 => n348, C2 => n347, A
                           => n353, ZN => n350);
   U753 : OAI211_X1 port map( C1 => n352, C2 => n351, A => n350, B => n349, ZN 
                           => n388);
   U754 : NAND2_X1 port map( A1 => n354, A2 => n353, ZN => n356);
   U755 : NOR3_X1 port map( A1 => n357, A2 => n356, A3 => n355, ZN => n382);
   U756 : AOI21_X1 port map( B1 => OP_A_22_port, B2 => n390, A => n409, ZN => 
                           n403);
   U757 : AND2_X1 port map( A1 => n404, A2 => n403, ZN => n359);
   U758 : AOI21_X1 port map( B1 => n358, B2 => OP_A_18_port, A => n398, ZN => 
                           n392);
   U759 : AND4_X1 port map( A1 => n393, A2 => n360, A3 => n359, A4 => n392, ZN 
                           => n386);
   U760 : OAI221_X1 port map( B1 => n388, B2 => n382, C1 => n388, C2 => n361, A
                           => n386, ZN => n444);
   U761 : OAI21_X1 port map( B1 => OP_B_26_port, B2 => n423, A => n422, ZN => 
                           n426);
   U762 : AOI211_X1 port map( C1 => OP_A_24_port, C2 => n417, A => n419, B => 
                           n426, ZN => n439);
   U763 : OAI21_X1 port map( B1 => OP_B_28_port, B2 => n412, A => n362, ZN => 
                           n416);
   U764 : NOR3_X1 port map( A1 => n428, A2 => n440, A3 => n416, ZN => n363);
   U765 : NAND2_X1 port map( A1 => n439, A2 => n363, ZN => n432);
   U766 : OAI21_X1 port map( B1 => n444, B2 => n432, A => OP_COMPARE_1_port, ZN
                           => n435);
   U767 : OAI22_X1 port map( A1 => n367, A2 => n366, B1 => n365, B2 => n364, ZN
                           => n377);
   U768 : NAND2_X1 port map( A1 => OP_B_4_port, A2 => n368, ZN => n370);
   U769 : OAI21_X1 port map( B1 => n371, B2 => n370, A => n369, ZN => n376);
   U770 : AOI21_X1 port map( B1 => OP_A_4_port, B2 => n1363, A => n371, ZN => 
                           n375);
   U771 : OAI21_X1 port map( B1 => OP_B_6_port, B2 => n372, A => n380, ZN => 
                           n373);
   U772 : INV_X1 port map( A => n373, ZN => n374);
   U773 : OAI221_X1 port map( B1 => n377, B2 => n376, C1 => n375, C2 => n376, A
                           => n374, ZN => n385);
   U774 : NOR2_X1 port map( A1 => OP_A_6_port, A2 => n378, ZN => n381);
   U775 : AOI21_X1 port map( B1 => n381, B2 => n380, A => n379, ZN => n384);
   U776 : INV_X1 port map( A => n382, ZN => n383);
   U777 : AOI21_X1 port map( B1 => n385, B2 => n384, A => n383, ZN => n387);
   U778 : OAI21_X1 port map( B1 => n388, B2 => n387, A => n386, ZN => n389);
   U779 : INV_X1 port map( A => n389, ZN => n443);
   U780 : OR2_X1 port map( A1 => OP_A_22_port, A2 => n390, ZN => n410);
   U781 : NAND2_X1 port map( A1 => n391, A2 => OP_B_18_port, ZN => n399);
   U782 : OAI211_X1 port map( C1 => n395, C2 => n394, A => n393, B => n392, ZN 
                           => n396);
   U783 : OAI211_X1 port map( C1 => n399, C2 => n398, A => n397, B => n396, ZN 
                           => n406);
   U784 : INV_X1 port map( A => n400, ZN => n401);
   U785 : OAI222_X1 port map( A1 => n402, A2 => n401, B1 => n402, B2 => 
                           OP_A_21_port, C1 => n401, C2 => OP_A_21_port, ZN => 
                           n405);
   U786 : OAI221_X1 port map( B1 => n406, B2 => n405, C1 => n404, C2 => n405, A
                           => n403, ZN => n407);
   U787 : OAI211_X1 port map( C1 => n410, C2 => n409, A => n408, B => n407, ZN 
                           => n455);
   U788 : INV_X1 port map( A => n455, ZN => n433);
   U789 : AOI21_X1 port map( B1 => n411, B2 => n450, A => n453, ZN => n431);
   U790 : NAND2_X1 port map( A1 => OP_B_28_port, A2 => n412, ZN => n414);
   U791 : OAI21_X1 port map( B1 => n415, B2 => n414, A => n413, ZN => n449);
   U792 : INV_X1 port map( A => n416, ZN => n448);
   U793 : OR2_X1 port map( A1 => OP_A_24_port, A2 => n417, ZN => n420);
   U794 : OAI21_X1 port map( B1 => n420, B2 => n419, A => n418, ZN => n421);
   U795 : INV_X1 port map( A => n421, ZN => n427);
   U796 : NAND3_X1 port map( A1 => OP_B_26_port, A2 => n423, A3 => n422, ZN => 
                           n424);
   U797 : OAI211_X1 port map( C1 => n427, C2 => n426, A => n425, B => n424, ZN 
                           => n447);
   U798 : NOR2_X1 port map( A1 => n428, A2 => n440, ZN => n429);
   U799 : OAI221_X1 port map( B1 => n449, B2 => n448, C1 => n449, C2 => n447, A
                           => n429, ZN => n430);
   U800 : OAI211_X1 port map( C1 => n433, C2 => n432, A => n431, B => n430, ZN 
                           => n434);
   U801 : AOI221_X1 port map( B1 => OP_COMPARE_2_port, B2 => n435, C1 => n443, 
                           C2 => n435, A => n434, ZN => n436);
   U802 : OAI21_X1 port map( B1 => n437, B2 => n436, A => OP_COMPARE_0_port, ZN
                           => n469);
   U803 : INV_X1 port map( A => n438, ZN => n467);
   U804 : INV_X1 port map( A => n439, ZN => n442);
   U805 : NOR2_X1 port map( A1 => n453, A2 => n440, ZN => n446);
   U806 : NAND2_X1 port map( A1 => n448, A2 => n446, ZN => n441);
   U807 : NOR2_X1 port map( A1 => n442, A2 => n441, ZN => n456);
   U808 : AOI21_X1 port map( B1 => n443, B2 => n456, A => OP_COMPARE_2_port, ZN
                           => n459);
   U809 : INV_X1 port map( A => n444, ZN => n445);
   U810 : AOI21_X1 port map( B1 => n445, B2 => n456, A => n460, ZN => n458);
   U811 : OAI221_X1 port map( B1 => n449, B2 => n448, C1 => n449, C2 => n447, A
                           => n446, ZN => n451);
   U812 : OAI211_X1 port map( C1 => n453, C2 => n452, A => n451, B => n450, ZN 
                           => n454);
   U813 : AOI21_X1 port map( B1 => n456, B2 => n455, A => n454, ZN => n457);
   U814 : OAI21_X1 port map( B1 => n459, B2 => n458, A => n457, ZN => n465);
   U815 : OAI211_X1 port map( C1 => n463, C2 => n462, A => n461, B => n460, ZN 
                           => n464);
   U816 : AOI21_X1 port map( B1 => n465, B2 => n464, A => OP_COMPARE_0_port, ZN
                           => n466);
   U817 : OAI21_X1 port map( B1 => n470, B2 => n467, A => n466, ZN => n468);
   U818 : OAI21_X1 port map( B1 => n470, B2 => n469, A => n468, ZN => n472);
   U819 : INV_X1 port map( A => N285, ZN => n471);
   U820 : AOI221_X1 port map( B1 => OP_COMPARE_3_port, B2 => n474, C1 => n473, 
                           C2 => n472, A => n471, ZN => n479);
   U821 : INV_X1 port map( A => N279, ZN => n1398);
   U822 : XOR2_X1 port map( A => n476, B => OP_Ci, Z => n477);
   U823 : NAND2_X1 port map( A1 => OP_LOGIC_1_port, A2 => n475, ZN => n1372);
   U824 : OAI22_X1 port map( A1 => n1398, A2 => n477, B1 => n1372, B2 => n476, 
                           ZN => n478);
   U825 : AOI211_X1 port map( C1 => n1367, C2 => n488, A => n479, B => n478, ZN
                           => n480);
   U826 : OAI211_X1 port map( C1 => n1159, C2 => n482, A => n481, B => n480, ZN
                           => Y(0));
   U827 : INV_X1 port map( A => n508, ZN => n483);
   U828 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_1, A => n483, 
                           ZN => n485);
   U829 : OAI22_X1 port map( A1 => n1396, A2 => n485, B1 => n1139, B2 => n484, 
                           ZN => n487);
   U830 : AOI22_X1 port map( A1 => n543, A2 => OP_A_0_port, B1 => OP_A_1_port, 
                           B2 => n56, ZN => n921);
   U831 : OAI22_X1 port map( A1 => n921, A2 => n1062, B1 => n520, B2 => n1369, 
                           ZN => n486);
   U832 : AOI211_X1 port map( C1 => n1330, C2 => OP1(1), A => n487, B => n486, 
                           ZN => n505);
   U833 : AOI22_X1 port map( A1 => OP_B_0_port, A2 => OP_A_0_port, B1 => OP_Ci,
                           B2 => n488, ZN => n522);
   U834 : INV_X1 port map( A => n522, ZN => n490);
   U835 : INV_X1 port map( A => n506, ZN => n489);
   U836 : AOI221_X1 port map( B1 => n522, B2 => n506, C1 => n490, C2 => n489, A
                           => n1398, ZN => n502);
   U837 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n55, ZN => n1353);
   U838 : NAND2_X1 port map( A1 => n492, A2 => OP_A_26_port, ZN => n1226);
   U839 : NAND2_X1 port map( A1 => OP_A_27_port, A2 => n554, ZN => n1289);
   U840 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => n56, ZN => n1166);
   U841 : NAND4_X1 port map( A1 => n1353, A2 => n1226, A3 => n1289, A4 => n1166
                           , ZN => n792);
   U842 : NAND2_X1 port map( A1 => n492, A2 => OP_A_30_port, ZN => n1354);
   U843 : NAND2_X1 port map( A1 => OP_A_29_port, A2 => n56, ZN => n1290);
   U844 : OAI211_X1 port map( C1 => n576, C2 => n1370, A => n1354, B => n1290, 
                           ZN => n491);
   U845 : AOI21_X1 port map( B1 => OP_SHIFT, B2 => n55, A => n491, ZN => n1298)
                           ;
   U846 : INV_X1 port map( A => n1298, ZN => n798);
   U847 : AOI22_X1 port map( A1 => n856, A2 => n792, B1 => n511, B2 => n798, ZN
                           => n494);
   U848 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => n55, ZN => n1225);
   U849 : NAND2_X1 port map( A1 => n492, A2 => OP_A_22_port, ZN => n1098);
   U850 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => n554, ZN => n1169);
   U851 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => n56, ZN => n1034);
   U852 : NAND4_X1 port map( A1 => n1225, A2 => n1098, A3 => n1169, A4 => n1034
                           , ZN => n793);
   U853 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => n55, ZN => n1097);
   U854 : NAND2_X1 port map( A1 => n543, A2 => OP_A_18_port, ZN => n972);
   U855 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => n554, ZN => n1037);
   U856 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n56, ZN => n913);
   U857 : NAND4_X1 port map( A1 => n1097, A2 => n972, A3 => n1037, A4 => n913, 
                           ZN => n795);
   U858 : AOI22_X1 port map( A1 => n64, A2 => n793, B1 => n895, B2 => n795, ZN 
                           => n493);
   U859 : NAND2_X1 port map( A1 => n494, A2 => n493, ZN => n923);
   U860 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => n55, ZN => n739);
   U861 : NAND2_X1 port map( A1 => OP_A_7_port, A2 => n554, ZN => n694);
   U862 : NAND2_X1 port map( A1 => OP_A_5_port, A2 => n56, ZN => n495);
   U863 : NAND4_X1 port map( A1 => n739, A2 => n659, A3 => n694, A4 => n495, ZN
                           => n597);
   U864 : AOI22_X1 port map( A1 => OP_B_4_port, A2 => n923, B1 => n1358, B2 => 
                           n597, ZN => n500);
   U865 : NAND2_X1 port map( A1 => OP_A_4_port, A2 => n55, ZN => n657);
   U866 : NAND2_X1 port map( A1 => OP_A_1_port, A2 => n56, ZN => n496);
   U867 : OAI211_X1 port map( C1 => n576, C2 => n551, A => n657, B => n496, ZN 
                           => n498);
   U868 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n55, ZN => n971);
   U869 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => n56, ZN => n803);
   U870 : NAND2_X1 port map( A1 => OP_A_15_port, A2 => n554, ZN => n916);
   U871 : NAND4_X1 port map( A1 => n853, A2 => n971, A3 => n803, A4 => n916, ZN
                           => n610);
   U872 : INV_X1 port map( A => n610, ZN => n796);
   U873 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => n55, ZN => n851);
   U874 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => n554, ZN => n804);
   U875 : NAND2_X1 port map( A1 => OP_A_9_port, A2 => n56, ZN => n695);
   U876 : AND4_X1 port map( A1 => n851, A2 => n741, A3 => n804, A4 => n695, ZN 
                           => n700);
   U877 : OAI22_X1 port map( A1 => n796, A2 => n892, B1 => n700, B2 => n567, ZN
                           => n497);
   U878 : AOI221_X1 port map( B1 => n553, B2 => n1360, C1 => n498, C2 => n1360,
                           A => n497, ZN => n499);
   U879 : AOI21_X1 port map( B1 => n500, B2 => n499, A => n1159, ZN => n501);
   U880 : AOI211_X1 port map( C1 => n1367, C2 => n503, A => n502, B => n501, ZN
                           => n504);
   U881 : OAI211_X1 port map( C1 => n1372, C2 => n506, A => n505, B => n504, ZN
                           => Y(1));
   U882 : INV_X1 port map( A => n524, ZN => n523);
   U883 : AOI22_X1 port map( A1 => n507, A2 => n1245, B1 => n1344, B2 => n523, 
                           ZN => n534);
   U884 : INV_X1 port map( A => n1139, ZN => n1348);
   U885 : NAND2_X1 port map( A1 => OP_A_2_port, A2 => n56, ZN => n516);
   U886 : OAI211_X1 port map( C1 => n576, C2 => n550, A => n508, B => n516, ZN 
                           => n821);
   U887 : AOI22_X1 port map( A1 => n1348, A2 => OP2(2), B1 => n1228, B2 => n821
                           , ZN => n533);
   U888 : AOI22_X1 port map( A1 => OP1(2), A2 => n1330, B1 => n1367, B2 => n547
                           , ZN => n532);
   U889 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => n56, ZN => n817);
   U890 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n604, ZN => n939);
   U891 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n55, ZN => n1004);
   U892 : NAND4_X1 port map( A1 => n891, A2 => n817, A3 => n939, A4 => n1004, 
                           ZN => n842);
   U893 : INV_X1 port map( A => n842, ZN => n729);
   U894 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => n604, ZN => n724);
   U895 : NAND2_X1 port map( A1 => OP_A_6_port, A2 => n56, ZN => n626);
   U896 : NAND2_X1 port map( A1 => OP_A_9_port, A2 => n55, ZN => n767);
   U897 : NAND4_X1 port map( A1 => n724, A2 => n626, A3 => n767, A4 => n676, ZN
                           => n619);
   U898 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => n604, ZN => n819);
   U899 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => n56, ZN => n725);
   U900 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => n55, ZN => n889);
   U901 : NAND4_X1 port map( A1 => n819, A2 => n725, A3 => n770, A4 => n889, ZN
                           => n722);
   U902 : AOI22_X1 port map( A1 => n1358, A2 => n619, B1 => n1350, B2 => n722, 
                           ZN => n519);
   U903 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => n604, ZN => n1206);
   U904 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => n56, ZN => n1057);
   U905 : NAND2_X1 port map( A1 => n543, A2 => OP_A_23_port, ZN => n1132);
   U906 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => n55, ZN => n1270);
   U907 : AND4_X1 port map( A1 => n1206, A2 => n1057, A3 => n1132, A4 => n1270,
                           ZN => n825);
   U908 : AOI22_X1 port map( A1 => OP_B_1_port, A2 => OP_SHIFT, B1 => 
                           OP_A_30_port, B2 => n56, ZN => n509);
   U909 : OAI21_X1 port map( B1 => n510, B2 => n1370, A => n509, ZN => n1328);
   U910 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => n604, ZN => n1060);
   U911 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => n56, ZN => n936);
   U912 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => n55, ZN => n1131);
   U913 : NAND2_X1 port map( A1 => n543, A2 => OP_A_19_port, ZN => n1005);
   U914 : NAND4_X1 port map( A1 => n1060, A2 => n936, A3 => n1131, A4 => n1005,
                           ZN => n827);
   U915 : AOI22_X1 port map( A1 => n511, A2 => n1328, B1 => n895, B2 => n827, 
                           ZN => n514);
   U916 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => n56, ZN => n1203);
   U917 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n554, ZN => n1320);
   U918 : NAND2_X1 port map( A1 => n543, A2 => OP_A_27_port, ZN => n1271);
   U919 : NAND2_X1 port map( A1 => OP_A_29_port, A2 => n55, ZN => n512);
   U920 : NAND4_X1 port map( A1 => n1203, A2 => n1320, A3 => n1271, A4 => n512,
                           ZN => n838);
   U921 : NAND2_X1 port map( A1 => n856, A2 => n838, ZN => n513);
   U922 : OAI211_X1 port map( C1 => n825, C2 => n743, A => n514, B => n513, ZN 
                           => n935);
   U923 : NAND2_X1 port map( A1 => OP_A_4_port, A2 => n554, ZN => n628);
   U924 : INV_X1 port map( A => n581, ZN => n515);
   U925 : NAND2_X1 port map( A1 => OP_A_5_port, A2 => n55, ZN => n674);
   U926 : NAND4_X1 port map( A1 => n628, A2 => n516, A3 => n515, A4 => n674, ZN
                           => n517);
   U927 : AOI22_X1 port map( A1 => OP_B_4_port, A2 => n935, B1 => n1360, B2 => 
                           n517, ZN => n518);
   U928 : OAI211_X1 port map( C1 => n729, C2 => n892, A => n519, B => n518, ZN 
                           => n530);
   U929 : OAI21_X1 port map( B1 => n522, B2 => n521, A => n520, ZN => n548);
   U930 : INV_X1 port map( A => n548, ZN => n525);
   U931 : AOI221_X1 port map( B1 => n525, B2 => n524, C1 => n548, C2 => n523, A
                           => n1398, ZN => n529);
   U932 : AOI211_X1 port map( C1 => n527, C2 => n526, A => n538, B => n1396, ZN
                           => n528);
   U933 : AOI211_X1 port map( C1 => N284, C2 => n530, A => n529, B => n528, ZN 
                           => n531);
   U934 : NAND4_X1 port map( A1 => n534, A2 => n533, A3 => n532, A4 => n531, ZN
                           => Y(2));
   U935 : XNOR2_X1 port map( A => n536, B => n535, ZN => n537);
   U936 : XNOR2_X1 port map( A => n538, B => n537, ZN => n564);
   U937 : INV_X1 port map( A => n1396, ZN => n987);
   U938 : INV_X1 port map( A => n987, ZN => n1284);
   U939 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => n554, ZN => n1227);
   U940 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => n56, ZN => n1096);
   U941 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => n55, ZN => n1287);
   U942 : NAND2_X1 port map( A1 => n543, A2 => OP_A_24_port, ZN => n1168);
   U943 : NAND4_X1 port map( A1 => n1227, A2 => n1096, A3 => n1287, A4 => n1168
                           , ZN => n864);
   U944 : NAND2_X1 port map( A1 => OP_A_29_port, A2 => n554, ZN => n1355);
   U945 : NAND2_X1 port map( A1 => OP_A_27_port, A2 => n56, ZN => n1224);
   U946 : NAND2_X1 port map( A1 => n543, A2 => OP_A_28_port, ZN => n1288);
   U947 : NAND3_X1 port map( A1 => n1355, A2 => n1224, A3 => n1288, ZN => n539)
                           ;
   U948 : AOI21_X1 port map( B1 => OP_A_30_port, B2 => n55, A => n539, ZN => 
                           n870);
   U949 : NOR2_X1 port map( A1 => n870, A2 => n742, ZN => n541);
   U950 : AOI22_X1 port map( A1 => n56, A2 => OP_A_31_port, B1 => OP_SHIFT, B2 
                           => n608, ZN => n1374);
   U951 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => n554, ZN => n1099);
   U952 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => n56, ZN => n970);
   U953 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => n55, ZN => n1167);
   U954 : NAND2_X1 port map( A1 => n543, A2 => OP_A_20_port, ZN => n1036);
   U955 : NAND4_X1 port map( A1 => n1099, A2 => n970, A3 => n1167, A4 => n1036,
                           ZN => n866);
   U956 : INV_X1 port map( A => n866, ZN => n749);
   U957 : OAI22_X1 port map( A1 => n1374, A2 => n858, B1 => n749, B2 => n766, 
                           ZN => n540);
   U958 : NAND2_X1 port map( A1 => OP_A_9_port, A2 => n554, ZN => n738);
   U959 : NAND2_X1 port map( A1 => OP_A_7_port, A2 => n56, ZN => n656);
   U960 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => n55, ZN => n802);
   U961 : NAND4_X1 port map( A1 => n738, A2 => n656, A3 => n802, A4 => n697, ZN
                           => n649);
   U962 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => n554, ZN => n852);
   U963 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => n56, ZN => n740);
   U964 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => n55, ZN => n914);
   U965 : NAND4_X1 port map( A1 => n852, A2 => n740, A3 => n805, A4 => n914, ZN
                           => n645);
   U966 : AOI22_X1 port map( A1 => n1358, A2 => n649, B1 => n1350, B2 => n645, 
                           ZN => n546);
   U967 : NAND2_X1 port map( A1 => OP_A_5_port, A2 => n554, ZN => n658);
   U968 : NAND2_X1 port map( A1 => OP_A_3_port, A2 => n56, ZN => n542);
   U969 : NAND2_X1 port map( A1 => OP_A_6_port, A2 => n55, ZN => n696);
   U970 : NAND4_X1 port map( A1 => n658, A2 => n542, A3 => n696, A4 => n605, ZN
                           => n544);
   U971 : NAND2_X1 port map( A1 => OP_A_15_port, A2 => n56, ZN => n850);
   U972 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n554, ZN => n973);
   U973 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => n55, ZN => n1035);
   U974 : NAND2_X1 port map( A1 => n543, A2 => OP_A_16_port, ZN => n915);
   U975 : NAND4_X1 port map( A1 => n850, A2 => n973, A3 => n1035, A4 => n915, 
                           ZN => n875);
   U976 : AOI22_X1 port map( A1 => n1360, A2 => n544, B1 => n1352, B2 => n875, 
                           ZN => n545);
   U977 : OAI211_X1 port map( C1 => n965, C2 => n1363, A => n546, B => n545, ZN
                           => n561);
   U978 : AOI22_X1 port map( A1 => OP_B_2_port, A2 => OP_A_2_port, B1 => n548, 
                           B2 => n547, ZN => n549);
   U979 : NOR2_X1 port map( A1 => n558, A2 => n549, ZN => n572);
   U980 : AOI211_X1 port map( C1 => n558, C2 => n549, A => n1398, B => n572, ZN
                           => n560);
   U981 : AOI22_X1 port map( A1 => n1348, A2 => OP2(3), B1 => n1347, B2 => 
                           OP1(3), ZN => n557);
   U982 : OAI22_X1 port map( A1 => n551, A2 => n608, B1 => n550, B2 => n578, ZN
                           => n552);
   U983 : AOI211_X1 port map( C1 => n554, C2 => OP_A_1_port, A => n553, B => 
                           n552, ZN => n967);
   U984 : INV_X1 port map( A => n967, ZN => n555);
   U985 : AOI22_X1 port map( A1 => OP_B_3_port, A2 => n1367, B1 => n1228, B2 =>
                           n555, ZN => n556);
   U986 : OAI211_X1 port map( C1 => n558, C2 => n1372, A => n557, B => n556, ZN
                           => n559);
   U987 : AOI211_X1 port map( C1 => N284, C2 => n561, A => n560, B => n559, ZN 
                           => n563);
   U988 : OAI221_X1 port map( B1 => n1367, B2 => OP_B_3_port, C1 => n1367, C2 
                           => n1245, A => OP_A_3_port, ZN => n562);
   U989 : OAI211_X1 port map( C1 => n564, C2 => n1284, A => n563, B => n562, ZN
                           => Y(3));
   U990 : NAND2_X1 port map( A1 => n1352, A2 => N284, ZN => n869);
   U991 : INV_X1 port map( A => n869, ZN => n839);
   U992 : AOI211_X1 port map( C1 => n566, C2 => intadd_0_SUM_0_port, A => n565,
                           B => n1396, ZN => n569);
   U993 : NOR2_X1 port map( A1 => n1159, A2 => n567, ZN => n865);
   U994 : INV_X1 port map( A => n865, ZN => n824);
   U995 : NOR2_X1 port map( A1 => n1159, A2 => n900, ZN => n867);
   U996 : INV_X1 port map( A => n867, ZN => n728);
   U997 : OAI22_X1 port map( A1 => n772, A2 => n824, B1 => n682, B2 => n728, ZN
                           => n568);
   U998 : AOI211_X1 port map( C1 => n839, C2 => n778, A => n569, B => n568, ZN 
                           => n590);
   U999 : INV_X1 port map( A => n574, ZN => n573);
   U1000 : NAND2_X1 port map( A1 => OP_B_4_port, A2 => N284, ZN => n765);
   U1001 : INV_X1 port map( A => n765, ZN => n745);
   U1002 : AOI22_X1 port map( A1 => n856, A2 => n1265, B1 => n63, B2 => n782, 
                           ZN => n570);
   U1003 : INV_X1 port map( A => OP_SHIFT, ZN => n1158);
   U1004 : NOR2_X1 port map( A1 => n858, A2 => n1158, ZN => n661);
   U1005 : INV_X1 port map( A => n661, ZN => n624);
   U1006 : OAI211_X1 port map( C1 => n785, C2 => n766, A => n570, B => n624, ZN
                           => n1009);
   U1007 : AOI22_X1 port map( A1 => n1344, A2 => n573, B1 => n745, B2 => n1009,
                           ZN => n589);
   U1008 : INV_X1 port map( A => n571, ZN => n599);
   U1009 : AOI22_X1 port map( A1 => n1245, A2 => n599, B1 => n1367, B2 => n598,
                           ZN => n588);
   U1010 : AOI21_X1 port map( B1 => OP_A_3_port, B2 => OP_B_3_port, A => n572, 
                           ZN => n575);
   U1011 : INV_X1 port map( A => n575, ZN => n600);
   U1012 : AOI221_X1 port map( B1 => n575, B2 => n574, C1 => n600, C2 => n573, 
                           A => n1398, ZN => n586);
   U1013 : OAI22_X1 port map( A1 => n579, A2 => n578, B1 => n577, B2 => n576, 
                           ZN => n580);
   U1014 : AOI211_X1 port map( C1 => n56, C2 => OP_A_4_port, A => n581, B => 
                           n580, ZN => n893);
   U1015 : AOI22_X1 port map( A1 => OP_B_2_port, A2 => n896, B1 => n893, B2 => 
                           n582, ZN => n771);
   U1016 : NAND2_X1 port map( A1 => n771, A2 => n1160, ZN => n1012);
   U1017 : NAND2_X1 port map( A1 => n1363, A2 => n1366, ZN => n886);
   U1018 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n1159, ZN => n1252);
   U1019 : NAND2_X1 port map( A1 => n895, A2 => n1252, ZN => n1373);
   U1020 : INV_X1 port map( A => n1373, ZN => n1329);
   U1021 : AOI22_X1 port map( A1 => n1330, A2 => OP1(4), B1 => n1329, B2 => 
                           n583, ZN => n584);
   U1022 : OAI21_X1 port map( B1 => n1012, B2 => n886, A => n584, ZN => n585);
   U1023 : AOI211_X1 port map( C1 => n1348, C2 => OP2(4), A => n586, B => n585,
                           ZN => n587);
   U1024 : NAND4_X1 port map( A1 => n590, A2 => n589, A3 => n588, A4 => n587, 
                           ZN => Y(4));
   U1025 : XNOR2_X1 port map( A => n592, B => n591, ZN => n593);
   U1026 : XNOR2_X1 port map( A => intadd_0_SUM_1_port, B => n593, ZN => n618);
   U1027 : INV_X1 port map( A => n795, ZN => n704);
   U1028 : OAI22_X1 port map( A1 => n704, A2 => n869, B1 => n700, B2 => n728, 
                           ZN => n596);
   U1029 : OAI22_X1 port map( A1 => n594, A2 => n1369, B1 => n1372, B2 => n601,
                           ZN => n595);
   U1030 : AOI211_X1 port map( C1 => n1329, C2 => n597, A => n596, B => n595, 
                           ZN => n617);
   U1031 : OAI21_X1 port map( B1 => n600, B2 => n599, A => n598, ZN => n602);
   U1032 : INV_X1 port map( A => n602, ZN => n634);
   U1033 : INV_X1 port map( A => n601, ZN => n603);
   U1034 : AOI221_X1 port map( B1 => n634, B2 => n603, C1 => n602, C2 => n601, 
                           A => n1398, ZN => n615);
   U1035 : INV_X1 port map( A => n886, ZN => n744);
   U1036 : AOI22_X1 port map( A1 => OP_A_3_port, A2 => n604, B1 => OP_A_2_port,
                           B2 => n55, ZN => n606);
   U1037 : OAI211_X1 port map( C1 => n608, C2 => n607, A => n606, B => n605, ZN
                           => n920);
   U1038 : INV_X1 port map( A => n920, ZN => n698);
   U1039 : OAI22_X1 port map( A1 => n698, A2 => n766, B1 => n921, B2 => n743, 
                           ZN => n1030);
   U1040 : AOI22_X1 port map( A1 => n1330, A2 => OP1(5), B1 => n744, B2 => 
                           n1030, ZN => n612);
   U1041 : AOI22_X1 port map( A1 => n854, A2 => n792, B1 => n895, B2 => n793, 
                           ZN => n609);
   U1042 : OAI211_X1 port map( C1 => n1298, C2 => n742, A => n609, B => n624, 
                           ZN => n1039);
   U1043 : AOI22_X1 port map( A1 => n745, A2 => n1039, B1 => n865, B2 => n610, 
                           ZN => n611);
   U1044 : OAI211_X1 port map( C1 => n1139, C2 => n613, A => n612, B => n611, 
                           ZN => n614);
   U1045 : AOI211_X1 port map( C1 => n1367, C2 => n633, A => n615, B => n614, 
                           ZN => n616);
   U1046 : OAI211_X1 port map( C1 => n1284, C2 => n618, A => n617, B => n616, 
                           ZN => Y(5));
   U1047 : INV_X1 port map( A => n637, ZN => n635);
   U1048 : AOI22_X1 port map( A1 => n1329, A2 => n619, B1 => n1344, B2 => n635,
                           ZN => n641);
   U1049 : AOI211_X1 port map( C1 => n621, C2 => intadd_1_SUM_0_port, A => n620
                           , B => n1396, ZN => n623);
   U1050 : OAI22_X1 port map( A1 => n652, A2 => n1368, B1 => n729, B2 => n824, 
                           ZN => n622);
   U1051 : AOI211_X1 port map( C1 => n867, C2 => n722, A => n623, B => n622, ZN
                           => n640);
   U1052 : AOI22_X1 port map( A1 => n856, A2 => n1328, B1 => n64, B2 => n838, 
                           ZN => n625);
   U1053 : OAI211_X1 port map( C1 => n825, C2 => n766, A => n625, B => n624, ZN
                           => n1066);
   U1054 : NAND4_X1 port map( A1 => n629, A2 => n628, A3 => n627, A4 => n626, 
                           ZN => n941);
   U1055 : AOI22_X1 port map( A1 => n63, A2 => n821, B1 => n895, B2 => n941, ZN
                           => n1063);
   U1056 : AOI22_X1 port map( A1 => n1348, A2 => OP2(6), B1 => n1330, B2 => 
                           OP1(6), ZN => n630);
   U1057 : OAI21_X1 port map( B1 => n1063, B2 => n886, A => n630, ZN => n632);
   U1058 : INV_X1 port map( A => n827, ZN => n730);
   U1059 : OAI22_X1 port map( A1 => n730, A2 => n869, B1 => n650, B2 => n1369, 
                           ZN => n631);
   U1060 : AOI211_X1 port map( C1 => n745, C2 => n1066, A => n632, B => n631, 
                           ZN => n639);
   U1061 : AOI22_X1 port map( A1 => OP_B_5_port, A2 => OP_A_5_port, B1 => n634,
                           B2 => n633, ZN => n651);
   U1062 : INV_X1 port map( A => n651, ZN => n636);
   U1063 : OAI221_X1 port map( B1 => n651, B2 => n637, C1 => n636, C2 => n635, 
                           A => N279, ZN => n638);
   U1064 : NAND4_X1 port map( A1 => n641, A2 => n640, A3 => n639, A4 => n638, 
                           ZN => Y(6));
   U1065 : XNOR2_X1 port map( A => n643, B => n642, ZN => n644);
   U1066 : XNOR2_X1 port map( A => intadd_1_SUM_1_port, B => n644, ZN => n670);
   U1067 : INV_X1 port map( A => n645, ZN => n748);
   U1068 : OAI22_X1 port map( A1 => n749, A2 => n869, B1 => n748, B2 => n728, 
                           ZN => n648);
   U1069 : OAI22_X1 port map( A1 => n646, A2 => n1369, B1 => n1372, B2 => n654,
                           ZN => n647);
   U1070 : AOI211_X1 port map( C1 => n1329, C2 => n649, A => n648, B => n647, 
                           ZN => n669);
   U1071 : OAI21_X1 port map( B1 => n652, B2 => n651, A => n650, ZN => n678);
   U1072 : INV_X1 port map( A => n678, ZN => n655);
   U1073 : INV_X1 port map( A => n654, ZN => n653);
   U1074 : AOI221_X1 port map( B1 => n655, B2 => n654, C1 => n678, C2 => n653, 
                           A => n1398, ZN => n667);
   U1075 : NAND4_X1 port map( A1 => n659, A2 => n658, A3 => n657, A4 => n656, 
                           ZN => n855);
   U1076 : INV_X1 port map( A => n855, ZN => n964);
   U1077 : OAI22_X1 port map( A1 => n964, A2 => n766, B1 => n967, B2 => n743, 
                           ZN => n1100);
   U1078 : AOI22_X1 port map( A1 => n1330, A2 => OP1(7), B1 => n744, B2 => 
                           n1100, ZN => n664);
   U1079 : OAI22_X1 port map( A1 => n1374, A2 => n742, B1 => n870, B2 => n743, 
                           ZN => n660);
   U1080 : AOI211_X1 port map( C1 => n895, C2 => n864, A => n661, B => n660, ZN
                           => n1107);
   U1081 : INV_X1 port map( A => n1107, ZN => n662);
   U1082 : AOI22_X1 port map( A1 => n745, A2 => n662, B1 => n865, B2 => n875, 
                           ZN => n663);
   U1083 : OAI211_X1 port map( C1 => n1139, C2 => n665, A => n664, B => n663, 
                           ZN => n666);
   U1084 : AOI211_X1 port map( C1 => n1367, C2 => n679, A => n667, B => n666, 
                           ZN => n668);
   U1085 : OAI211_X1 port map( C1 => n1284, C2 => n670, A => n669, B => n668, 
                           ZN => Y(7));
   U1086 : AOI22_X1 port map( A1 => n64, A2 => n1265, B1 => n895, B2 => n782, 
                           ZN => n671);
   U1087 : OAI21_X1 port map( B1 => n1160, B2 => n1158, A => n671, ZN => n1135)
                           ;
   U1088 : AOI22_X1 port map( A1 => n745, A2 => n1135, B1 => n1367, B2 => n672,
                           ZN => n691);
   U1089 : INV_X1 port map( A => n712, ZN => n677);
   U1090 : NAND4_X1 port map( A1 => n676, A2 => n675, A3 => n674, A4 => n673, 
                           ZN => n1007);
   U1091 : INV_X1 port map( A => n1007, ZN => n906);
   U1092 : OAI222_X1 port map( A1 => n896, A2 => n742, B1 => n766, B2 => n906, 
                           C1 => n743, C2 => n893, ZN => n1134);
   U1093 : AOI22_X1 port map( A1 => n677, A2 => n1245, B1 => n744, B2 => n1134,
                           ZN => n690);
   U1094 : AOI22_X1 port map( A1 => OP_B_7_port, A2 => OP_A_7_port, B1 => n679,
                           B2 => n678, ZN => n713);
   U1095 : NOR2_X1 port map( A1 => n713, A2 => n681, ZN => n680);
   U1096 : AOI211_X1 port map( C1 => n713, C2 => n681, A => n1398, B => n680, 
                           ZN => n688);
   U1097 : OAI22_X1 port map( A1 => n682, A2 => n1373, B1 => n681, B2 => n1372,
                           ZN => n687);
   U1098 : AOI22_X1 port map( A1 => n1348, A2 => OP2(8), B1 => n1330, B2 => 
                           OP1(8), ZN => n685);
   U1099 : OAI22_X1 port map( A1 => n785, A2 => n869, B1 => n772, B2 => n728, 
                           ZN => n683);
   U1100 : AOI21_X1 port map( B1 => n865, B2 => n778, A => n683, ZN => n684);
   U1101 : OAI211_X1 port map( C1 => intadd_2_SUM_0_port, C2 => n1284, A => 
                           n685, B => n684, ZN => n686);
   U1102 : NOR3_X1 port map( A1 => n688, A2 => n687, A3 => n686, ZN => n689);
   U1103 : NAND3_X1 port map( A1 => n691, A2 => n690, A3 => n689, ZN => Y(8));
   U1104 : OAI22_X1 port map( A1 => intadd_2_SUM_1_port, A2 => n1284, B1 => 
                           n1139, B2 => n692, ZN => n693);
   U1105 : AOI21_X1 port map( B1 => n703, B2 => n1344, A => n693, ZN => n711);
   U1106 : NAND4_X1 port map( A1 => n697, A2 => n696, A3 => n695, A4 => n694, 
                           ZN => n1038);
   U1107 : INV_X1 port map( A => n1038, ZN => n932);
   U1108 : OAI222_X1 port map( A1 => n743, A2 => n698, B1 => n766, B2 => n932, 
                           C1 => n742, C2 => n921, ZN => n1161);
   U1109 : AOI22_X1 port map( A1 => n1330, A2 => OP1(9), B1 => n744, B2 => 
                           n1161, ZN => n710);
   U1110 : NOR2_X1 port map( A1 => n1158, A2 => n765, ZN => n1121);
   U1111 : INV_X1 port map( A => n1121, ZN => n1109);
   U1112 : NOR2_X1 port map( A1 => n1160, A2 => n1109, ZN => n754);
   U1113 : INV_X1 port map( A => n699, ZN => n714);
   U1114 : OAI22_X1 port map( A1 => n700, A2 => n1373, B1 => n714, B2 => n1369,
                           ZN => n701);
   U1115 : AOI211_X1 port map( C1 => n839, C2 => n793, A => n754, B => n701, ZN
                           => n709);
   U1116 : AOI21_X1 port map( B1 => n713, B2 => n712, A => n716, ZN => n702);
   U1117 : XOR2_X1 port map( A => n703, B => n702, Z => n707);
   U1118 : OAI22_X1 port map( A1 => n704, A2 => n824, B1 => n715, B2 => n1368, 
                           ZN => n706);
   U1119 : AOI22_X1 port map( A1 => n854, A2 => n798, B1 => n895, B2 => n792, 
                           ZN => n1174);
   U1120 : OAI22_X1 port map( A1 => n1174, A2 => n765, B1 => n796, B2 => n728, 
                           ZN => n705);
   U1121 : AOI211_X1 port map( C1 => n707, C2 => N279, A => n706, B => n705, ZN
                           => n708);
   U1122 : NAND4_X1 port map( A1 => n711, A2 => n710, A3 => n709, A4 => n708, 
                           ZN => Y(9));
   U1123 : NAND2_X1 port map( A1 => n714, A2 => n712, ZN => n719);
   U1124 : INV_X1 port map( A => n713, ZN => n718);
   U1125 : OAI21_X1 port map( B1 => n716, B2 => n715, A => n714, ZN => n717);
   U1126 : OAI21_X1 port map( B1 => n719, B2 => n718, A => n717, ZN => n757);
   U1127 : XNOR2_X1 port map( A => n720, B => n757, ZN => n737);
   U1128 : NOR2_X1 port map( A1 => OP_A_10_port, A2 => OP_B_10_port, ZN => n758
                           );
   U1129 : OAI22_X1 port map( A1 => n758, A2 => n1368, B1 => n1372, B2 => n720,
                           ZN => n721);
   U1130 : AOI211_X1 port map( C1 => n1329, C2 => n722, A => n754, B => n721, 
                           ZN => n736);
   U1131 : AOI22_X1 port map( A1 => n1348, A2 => OP2(10), B1 => n1347, B2 => 
                           OP1(10), ZN => n723);
   U1132 : OAI21_X1 port map( B1 => n756, B2 => n1369, A => n723, ZN => n734);
   U1133 : OAI22_X1 port map( A1 => n825, A2 => n869, B1 => intadd_2_SUM_2_port
                           , B2 => n1284, ZN => n733);
   U1134 : NAND4_X1 port map( A1 => n727, A2 => n726, A3 => n725, A4 => n724, 
                           ZN => n940);
   U1135 : AOI222_X1 port map( A1 => n821, A2 => n856, B1 => n941, B2 => n854, 
                           C1 => n940, C2 => n895, ZN => n1212);
   U1136 : AOI22_X1 port map( A1 => n63, A2 => n1328, B1 => n895, B2 => n838, 
                           ZN => n1182);
   U1137 : OAI22_X1 port map( A1 => n1212, A2 => n886, B1 => n1182, B2 => n765,
                           ZN => n732);
   U1138 : OAI22_X1 port map( A1 => n730, A2 => n824, B1 => n729, B2 => n728, 
                           ZN => n731);
   U1139 : NOR4_X1 port map( A1 => n734, A2 => n733, A3 => n732, A4 => n731, ZN
                           => n735);
   U1140 : OAI211_X1 port map( C1 => n1398, C2 => n737, A => n736, B => n735, 
                           ZN => Y(10));
   U1141 : AOI22_X1 port map( A1 => n867, A2 => n875, B1 => n839, B2 => n864, 
                           ZN => n764);
   U1142 : OAI22_X1 port map( A1 => n1374, A2 => n743, B1 => n870, B2 => n766, 
                           ZN => n1251);
   U1143 : NAND4_X1 port map( A1 => n741, A2 => n740, A3 => n739, A4 => n738, 
                           ZN => n974);
   U1144 : INV_X1 port map( A => n974, ZN => n1112);
   U1145 : OAI222_X1 port map( A1 => n743, A2 => n964, B1 => n766, B2 => n1112,
                           C1 => n742, C2 => n967, ZN => n1243);
   U1146 : AOI22_X1 port map( A1 => n745, A2 => n1251, B1 => n744, B2 => n1243,
                           ZN => n763);
   U1147 : AOI22_X1 port map( A1 => OP1(11), A2 => n1330, B1 => n1367, B2 => 
                           n774, ZN => n747);
   U1148 : NAND2_X1 port map( A1 => n1348, A2 => OP2(11), ZN => n746);
   U1149 : OAI211_X1 port map( C1 => intadd_2_SUM_3_port, C2 => n1284, A => 
                           n747, B => n746, ZN => n753);
   U1150 : OAI22_X1 port map( A1 => n749, A2 => n824, B1 => n748, B2 => n1373, 
                           ZN => n752);
   U1151 : OAI22_X1 port map( A1 => n750, A2 => n1369, B1 => n1372, B2 => n755,
                           ZN => n751);
   U1152 : NOR4_X1 port map( A1 => n754, A2 => n753, A3 => n752, A4 => n751, ZN
                           => n762);
   U1153 : INV_X1 port map( A => n755, ZN => n760);
   U1154 : OAI21_X1 port map( B1 => n758, B2 => n757, A => n756, ZN => n775);
   U1155 : AOI21_X1 port map( B1 => n760, B2 => n775, A => n1398, ZN => n759);
   U1156 : OAI21_X1 port map( B1 => n760, B2 => n775, A => n759, ZN => n761);
   U1157 : NAND4_X1 port map( A1 => n764, A2 => n763, A3 => n762, A4 => n761, 
                           ZN => Y(11));
   U1158 : NOR2_X1 port map( A1 => n766, A2 => n765, ZN => n877);
   U1159 : NAND4_X1 port map( A1 => n770, A2 => n769, A3 => n768, A4 => n767, 
                           ZN => n1119);
   U1160 : AOI222_X1 port map( A1 => n1007, A2 => n63, B1 => OP_B_3_port, B2 =>
                           n771, C1 => n1119, C2 => n895, ZN => n1278);
   U1161 : OAI22_X1 port map( A1 => n1278, A2 => n886, B1 => n772, B2 => n1373,
                           ZN => n773);
   U1162 : AOI21_X1 port map( B1 => n877, B2 => n1265, A => n773, ZN => n791);
   U1163 : AOI22_X1 port map( A1 => OP_A_11_port, A2 => OP_B_11_port, B1 => 
                           n775, B2 => n774, ZN => n829);
   U1164 : NOR2_X1 port map( A1 => n829, A2 => n780, ZN => n776);
   U1165 : AOI211_X1 port map( C1 => n829, C2 => n780, A => n1398, B => n776, 
                           ZN => n789);
   U1166 : OAI22_X1 port map( A1 => intadd_2_SUM_4_port, A2 => n1284, B1 => 
                           n1139, B2 => n777, ZN => n788);
   U1167 : AOI22_X1 port map( A1 => n1330, A2 => OP1(12), B1 => n867, B2 => 
                           n778, ZN => n779);
   U1168 : OAI21_X1 port map( B1 => n780, B2 => n1372, A => n779, ZN => n787);
   U1169 : AOI22_X1 port map( A1 => n839, A2 => n782, B1 => n1367, B2 => n781, 
                           ZN => n784);
   U1170 : NOR2_X1 port map( A1 => n895, A2 => n1109, ZN => n862);
   U1171 : INV_X1 port map( A => n862, ZN => n783);
   U1172 : OAI211_X1 port map( C1 => n785, C2 => n824, A => n784, B => n783, ZN
                           => n786);
   U1173 : NOR4_X1 port map( A1 => n789, A2 => n788, A3 => n787, A4 => n786, ZN
                           => n790);
   U1174 : OAI211_X1 port map( C1 => n828, C2 => n1369, A => n791, B => n790, 
                           ZN => Y(12));
   U1175 : AOI22_X1 port map( A1 => n865, A2 => n793, B1 => n839, B2 => n792, 
                           ZN => n816);
   U1176 : AOI22_X1 port map( A1 => n867, A2 => n795, B1 => n1367, B2 => n794, 
                           ZN => n815);
   U1177 : OAI22_X1 port map( A1 => n796, A2 => n1373, B1 => n830, B2 => n1369,
                           ZN => n797);
   U1178 : AOI211_X1 port map( C1 => n877, C2 => n798, A => n862, B => n797, ZN
                           => n814);
   U1179 : INV_X1 port map( A => n799, ZN => n808);
   U1180 : AOI21_X1 port map( B1 => n829, B2 => n828, A => n831, ZN => n800);
   U1181 : XOR2_X1 port map( A => n808, B => n800, Z => n812);
   U1182 : OAI22_X1 port map( A1 => intadd_2_SUM_5_port, A2 => n1284, B1 => 
                           n1139, B2 => n801, ZN => n811);
   U1183 : NAND4_X1 port map( A1 => n805, A2 => n804, A3 => n803, A4 => n802, 
                           ZN => n1170);
   U1184 : AOI22_X1 port map( A1 => n856, A2 => n920, B1 => n854, B2 => n1038, 
                           ZN => n806);
   U1185 : OAI21_X1 port map( B1 => n921, B2 => n858, A => n806, ZN => n807);
   U1186 : AOI21_X1 port map( B1 => n895, B2 => n1170, A => n807, ZN => n1295);
   U1187 : AOI22_X1 port map( A1 => n808, A2 => n1344, B1 => n1347, B2 => 
                           OP1(13), ZN => n809);
   U1188 : OAI21_X1 port map( B1 => n1295, B2 => n886, A => n809, ZN => n810);
   U1189 : AOI211_X1 port map( C1 => n812, C2 => N279, A => n811, B => n810, ZN
                           => n813);
   U1190 : NAND4_X1 port map( A1 => n816, A2 => n815, A3 => n814, A4 => n813, 
                           ZN => Y(13));
   U1191 : NOR2_X1 port map( A1 => OP_A_14_port, A2 => OP_B_14_port, ZN => n873
                           );
   U1192 : NAND4_X1 port map( A1 => n820, A2 => n819, A3 => n818, A4 => n817, 
                           ZN => n1207);
   U1193 : INV_X1 port map( A => n821, ZN => n933);
   U1194 : AOI22_X1 port map( A1 => n856, A2 => n941, B1 => n63, B2 => n940, ZN
                           => n822);
   U1195 : OAI21_X1 port map( B1 => n933, B2 => n858, A => n822, ZN => n823);
   U1196 : AOI21_X1 port map( B1 => n895, B2 => n1207, A => n823, ZN => n1326);
   U1197 : OAI22_X1 port map( A1 => n825, A2 => n824, B1 => n1326, B2 => n886, 
                           ZN => n826);
   U1198 : AOI21_X1 port map( B1 => n867, B2 => n827, A => n826, ZN => n849);
   U1199 : INV_X1 port map( A => n836, ZN => n843);
   U1200 : NAND2_X1 port map( A1 => n830, A2 => n828, ZN => n835);
   U1201 : INV_X1 port map( A => n829, ZN => n834);
   U1202 : OAI21_X1 port map( B1 => n832, B2 => n831, A => n830, ZN => n833);
   U1203 : OAI21_X1 port map( B1 => n835, B2 => n834, A => n833, ZN => n872);
   U1204 : INV_X1 port map( A => n872, ZN => n837);
   U1205 : AOI221_X1 port map( B1 => n843, B2 => n837, C1 => n836, C2 => n872, 
                           A => n1398, ZN => n847);
   U1206 : AOI22_X1 port map( A1 => n1348, A2 => OP2(14), B1 => n1347, B2 => 
                           OP1(14), ZN => n841);
   U1207 : AOI22_X1 port map( A1 => n839, A2 => n838, B1 => n877, B2 => n1328, 
                           ZN => n840);
   U1208 : OAI211_X1 port map( C1 => intadd_2_SUM_6_port, C2 => n1284, A => 
                           n841, B => n840, ZN => n846);
   U1209 : AOI22_X1 port map( A1 => n843, A2 => n1344, B1 => n1329, B2 => n842,
                           ZN => n844);
   U1210 : OAI21_X1 port map( B1 => n871, B2 => n1369, A => n844, ZN => n845);
   U1211 : NOR4_X1 port map( A1 => n862, A2 => n847, A3 => n846, A4 => n845, ZN
                           => n848);
   U1212 : OAI211_X1 port map( C1 => n873, C2 => n1368, A => n849, B => n848, 
                           ZN => Y(14));
   U1213 : NAND4_X1 port map( A1 => n853, A2 => n852, A3 => n851, A4 => n850, 
                           ZN => n1229);
   U1214 : AOI22_X1 port map( A1 => n856, A2 => n855, B1 => n64, B2 => n974, ZN
                           => n857);
   U1215 : OAI21_X1 port map( B1 => n967, B2 => n858, A => n857, ZN => n859);
   U1216 : AOI21_X1 port map( B1 => n895, B2 => n1229, A => n859, ZN => n1364);
   U1217 : OAI22_X1 port map( A1 => intadd_2_SUM_7_port, A2 => n1284, B1 => 
                           n1139, B2 => n860, ZN => n861);
   U1218 : AOI211_X1 port map( C1 => n1330, C2 => OP1(15), A => n862, B => n861
                           , ZN => n885);
   U1219 : INV_X1 port map( A => n863, ZN => n902);
   U1220 : AOI22_X1 port map( A1 => n867, A2 => n866, B1 => n865, B2 => n864, 
                           ZN => n868);
   U1221 : OAI21_X1 port map( B1 => n870, B2 => n869, A => n868, ZN => n883);
   U1222 : OAI21_X1 port map( B1 => n873, B2 => n872, A => n871, ZN => n903);
   U1223 : XNOR2_X1 port map( A => n874, B => n903, ZN => n881);
   U1224 : AOI22_X1 port map( A1 => n1329, A2 => n875, B1 => n1344, B2 => n874,
                           ZN => n880);
   U1225 : INV_X1 port map( A => n1374, ZN => n876);
   U1226 : AOI22_X1 port map( A1 => n878, A2 => n1245, B1 => n877, B2 => n876, 
                           ZN => n879);
   U1227 : OAI211_X1 port map( C1 => n1398, C2 => n881, A => n880, B => n879, 
                           ZN => n882);
   U1228 : AOI211_X1 port map( C1 => n1367, C2 => n902, A => n883, B => n882, 
                           ZN => n884);
   U1229 : OAI211_X1 port map( C1 => n1364, C2 => n886, A => n885, B => n884, 
                           ZN => Y(15));
   U1230 : AOI22_X1 port map( A1 => n1348, A2 => OP2(16), B1 => n1347, B2 => 
                           OP1(16), ZN => n912);
   U1231 : OAI22_X1 port map( A1 => intadd_2_SUM_8_port, A2 => n1284, B1 => 
                           n950, B2 => n1369, ZN => n887);
   U1232 : NOR2_X1 port map( A1 => n1121, A2 => n887, ZN => n911);
   U1233 : NAND4_X1 port map( A1 => n891, A2 => n890, A3 => n889, A4 => n888, 
                           ZN => n1268);
   U1234 : INV_X1 port map( A => n1268, ZN => n894);
   U1235 : NOR2_X1 port map( A1 => n901, A2 => n892, ZN => n1230);
   U1236 : INV_X1 port map( A => n1230, ZN => n1111);
   U1237 : OAI22_X1 port map( A1 => n894, A2 => n1062, B1 => n893, B2 => n1111,
                           ZN => n898);
   U1238 : NOR2_X1 port map( A1 => n901, A2 => n1363, ZN => n1244);
   U1239 : NAND2_X1 port map( A1 => n895, A2 => n1244, ZN => n966);
   U1240 : OAI22_X1 port map( A1 => n953, A2 => n1368, B1 => n966, B2 => n896, 
                           ZN => n897);
   U1241 : AOI211_X1 port map( C1 => n1252, C2 => n899, A => n898, B => n897, 
                           ZN => n910);
   U1242 : NOR2_X1 port map( A1 => n901, A2 => n900, ZN => n1242);
   U1243 : AOI22_X1 port map( A1 => OP_A_15_port, A2 => OP_B_15_port, B1 => 
                           n903, B2 => n902, ZN => n951);
   U1244 : NOR2_X1 port map( A1 => n951, A2 => n905, ZN => n904);
   U1245 : AOI211_X1 port map( C1 => n951, C2 => n905, A => n1398, B => n904, 
                           ZN => n908);
   U1246 : NAND2_X1 port map( A1 => n1350, A2 => n1366, ZN => n1233);
   U1247 : OAI22_X1 port map( A1 => n906, A2 => n1233, B1 => n905, B2 => n1372,
                           ZN => n907);
   U1248 : AOI211_X1 port map( C1 => n1242, C2 => n1119, A => n908, B => n907, 
                           ZN => n909);
   U1249 : NAND4_X1 port map( A1 => n912, A2 => n911, A3 => n910, A4 => n909, 
                           ZN => Y(16));
   U1250 : NAND4_X1 port map( A1 => n916, A2 => n915, A3 => n914, A4 => n913, 
                           ZN => n1285);
   U1251 : AOI22_X1 port map( A1 => n919, A2 => n1344, B1 => n1228, B2 => n1285
                           , ZN => n931);
   U1252 : AOI22_X1 port map( A1 => n1348, A2 => OP2(17), B1 => n1347, B2 => 
                           OP1(17), ZN => n917);
   U1253 : OAI211_X1 port map( C1 => intadd_2_SUM_9_port, C2 => n1284, A => 
                           n917, B => n1109, ZN => n928);
   U1254 : AOI21_X1 port map( B1 => n951, B2 => n950, A => n953, ZN => n918);
   U1255 : XNOR2_X1 port map( A => n919, B => n918, ZN => n926);
   U1256 : AOI22_X1 port map( A1 => n1230, A2 => n920, B1 => n1242, B2 => n1170
                           , ZN => n925);
   U1257 : OAI22_X1 port map( A1 => n921, A2 => n966, B1 => n954, B2 => n1368, 
                           ZN => n922);
   U1258 : AOI21_X1 port map( B1 => n1252, B2 => n923, A => n922, ZN => n924);
   U1259 : OAI211_X1 port map( C1 => n1398, C2 => n926, A => n925, B => n924, 
                           ZN => n927);
   U1260 : AOI211_X1 port map( C1 => n929, C2 => n1245, A => n928, B => n927, 
                           ZN => n930);
   U1261 : OAI211_X1 port map( C1 => n932, C2 => n1233, A => n931, B => n930, 
                           ZN => Y(17));
   U1262 : OAI22_X1 port map( A1 => n933, A2 => n966, B1 => n983, B2 => n1368, 
                           ZN => n934);
   U1263 : AOI211_X1 port map( C1 => n1252, C2 => n935, A => n1121, B => n934, 
                           ZN => n962);
   U1264 : NAND4_X1 port map( A1 => n939, A2 => n938, A3 => n937, A4 => n936, 
                           ZN => n1316);
   U1265 : INV_X1 port map( A => n1316, ZN => n1210);
   U1266 : INV_X1 port map( A => n940, ZN => n1069);
   U1267 : OAI22_X1 port map( A1 => n1210, A2 => n1062, B1 => n1069, B2 => 
                           n1233, ZN => n948);
   U1268 : INV_X1 port map( A => n941, ZN => n946);
   U1269 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_18, B1 => 
                           OP_A_12_port, B2 => n61, C1 => OP_A_11_port, C2 => 
                           n1028, ZN => n979);
   U1270 : XOR2_X1 port map( A => n979, B => intadd_1_SUM_12_port, Z => n942);
   U1271 : XNOR2_X1 port map( A => intadd_2_n1, B => n942, ZN => n943);
   U1272 : AOI22_X1 port map( A1 => n987, A2 => n943, B1 => n1242, B2 => n1207,
                           ZN => n945);
   U1273 : AOI22_X1 port map( A1 => n1348, A2 => OP2(18), B1 => n1347, B2 => 
                           OP1(18), ZN => n944);
   U1274 : OAI211_X1 port map( C1 => n946, C2 => n1111, A => n945, B => n944, 
                           ZN => n947);
   U1275 : AOI211_X1 port map( C1 => n949, C2 => n1245, A => n948, B => n947, 
                           ZN => n961);
   U1276 : NAND2_X1 port map( A1 => n952, A2 => n950, ZN => n957);
   U1277 : INV_X1 port map( A => n951, ZN => n956);
   U1278 : OAI21_X1 port map( B1 => n954, B2 => n953, A => n952, ZN => n955);
   U1279 : OAI21_X1 port map( B1 => n957, B2 => n956, A => n955, ZN => n982);
   U1280 : XNOR2_X1 port map( A => n959, B => n982, ZN => n958);
   U1281 : AOI22_X1 port map( A1 => n959, A2 => n1344, B1 => N279, B2 => n958, 
                           ZN => n960);
   U1282 : NAND3_X1 port map( A1 => n962, A2 => n961, A3 => n960, ZN => Y(18));
   U1283 : AOI22_X1 port map( A1 => n1348, A2 => OP2(19), B1 => n1347, B2 => 
                           OP1(19), ZN => n963);
   U1284 : OAI21_X1 port map( B1 => n964, B2 => n1111, A => n963, ZN => n969);
   U1285 : INV_X1 port map( A => n1252, ZN => n1181);
   U1286 : OAI22_X1 port map( A1 => n967, A2 => n966, B1 => n965, B2 => n1181, 
                           ZN => n968);
   U1287 : AOI211_X1 port map( C1 => n1367, C2 => n992, A => n969, B => n968, 
                           ZN => n991);
   U1288 : NAND4_X1 port map( A1 => n973, A2 => n972, A3 => n971, A4 => n970, 
                           ZN => n1351);
   U1289 : INV_X1 port map( A => n1233, ZN => n1122);
   U1290 : AOI22_X1 port map( A1 => n1228, A2 => n1351, B1 => n1122, B2 => n974
                           , ZN => n990);
   U1291 : OAI22_X1 port map( A1 => n976, A2 => n1369, B1 => n1372, B2 => n975,
                           ZN => n977);
   U1292 : AOI211_X1 port map( C1 => n1242, C2 => n1229, A => n1121, B => n977,
                           ZN => n989);
   U1293 : AND2_X1 port map( A1 => intadd_1_SUM_12_port, A2 => intadd_2_n1, ZN 
                           => n978);
   U1294 : OAI22_X1 port map( A1 => n979, A2 => n978, B1 => 
                           intadd_1_SUM_12_port, B2 => intadd_2_n1, ZN => n995)
                           ;
   U1295 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_19, B1 => 
                           OP_A_12_port, B2 => n1028, C1 => n61, C2 => 
                           OP_A_13_port, ZN => n998);
   U1296 : XNOR2_X1 port map( A => intadd_1_SUM_13_port, B => n998, ZN => n980)
                           ;
   U1297 : XNOR2_X1 port map( A => n995, B => n980, ZN => n986);
   U1298 : OAI21_X1 port map( B1 => n983, B2 => n982, A => n981, ZN => n993);
   U1299 : XOR2_X1 port map( A => n984, B => n993, Z => n985);
   U1300 : AOI22_X1 port map( A1 => n987, A2 => n986, B1 => n985, B2 => N279, 
                           ZN => n988);
   U1301 : NAND4_X1 port map( A1 => n991, A2 => n990, A3 => n989, A4 => n988, 
                           ZN => Y(19));
   U1302 : AOI22_X1 port map( A1 => n1242, A2 => n1268, B1 => n1122, B2 => 
                           n1119, ZN => n1018);
   U1303 : AOI22_X1 port map( A1 => OP_A_19_port, A2 => OP_B_19_port, B1 => 
                           n993, B2 => n992, ZN => n1048);
   U1304 : NOR2_X1 port map( A1 => n1048, A2 => n1019, ZN => n994);
   U1305 : AOI211_X1 port map( C1 => n1048, C2 => n1019, A => n1398, B => n994,
                           ZN => n1016);
   U1306 : INV_X1 port map( A => n995, ZN => n999);
   U1307 : INV_X1 port map( A => intadd_1_SUM_13_port, ZN => n996);
   U1308 : NAND2_X1 port map( A1 => n996, A2 => n995, ZN => n997);
   U1309 : AOI22_X1 port map( A1 => intadd_1_SUM_13_port, A2 => n999, B1 => 
                           n998, B2 => n997, ZN => n1027);
   U1310 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_20, B1 => n61, B2 
                           => OP_A_14_port, C1 => n1028, C2 => OP_A_13_port, ZN
                           => n1023);
   U1311 : INV_X1 port map( A => intadd_1_SUM_14_port, ZN => n1026);
   U1312 : XNOR2_X1 port map( A => n1023, B => n1026, ZN => n1000);
   U1313 : XNOR2_X1 port map( A => n1027, B => n1000, ZN => n1001);
   U1314 : NOR2_X1 port map( A1 => n1001, A2 => n1284, ZN => n1015);
   U1315 : AOI22_X1 port map( A1 => n1348, A2 => OP2(20), B1 => n1347, B2 => 
                           OP1(20), ZN => n1002);
   U1316 : OAI211_X1 port map( C1 => n1369, C2 => n1047, A => n1002, B => n1109
                           , ZN => n1014);
   U1317 : INV_X1 port map( A => n1244, ZN => n1211);
   U1318 : NAND4_X1 port map( A1 => n1006, A2 => n1005, A3 => n1004, A4 => 
                           n1003, ZN => n1269);
   U1319 : AOI22_X1 port map( A1 => n1228, A2 => n1269, B1 => n1230, B2 => 
                           n1007, ZN => n1011);
   U1320 : AOI22_X1 port map( A1 => n1252, A2 => n1009, B1 => n1367, B2 => 
                           n1008, ZN => n1010);
   U1321 : OAI211_X1 port map( C1 => n1211, C2 => n1012, A => n1011, B => n1010
                           , ZN => n1013);
   U1322 : NOR4_X1 port map( A1 => n1016, A2 => n1015, A3 => n1014, A4 => n1013
                           , ZN => n1017);
   U1323 : OAI211_X1 port map( C1 => n1019, C2 => n1372, A => n1018, B => n1017
                           , ZN => Y(20));
   U1324 : AOI21_X1 port map( B1 => n1048, B2 => n1047, A => n1050, ZN => n1020
                           );
   U1325 : XNOR2_X1 port map( A => n1021, B => n1020, ZN => n1046);
   U1326 : AOI22_X1 port map( A1 => n1022, A2 => n1245, B1 => n1021, B2 => 
                           n1344, ZN => n1045);
   U1327 : INV_X1 port map( A => n1027, ZN => n1024);
   U1328 : OAI21_X1 port map( B1 => intadd_1_SUM_14_port, B2 => n1024, A => 
                           n1023, ZN => n1025);
   U1329 : OAI21_X1 port map( B1 => n1027, B2 => n1026, A => n1025, ZN => n1077
                           );
   U1330 : INV_X1 port map( A => n1077, ZN => n1074);
   U1331 : AOI222_X1 port map( A1 => OP_A_15_port, A2 => n61, B1 => n1414, B2 
                           => C429_DATA4_21, C1 => n1028, C2 => OP_A_14_port, 
                           ZN => n1076);
   U1332 : INV_X1 port map( A => intadd_1_SUM_15_port, ZN => n1073);
   U1333 : XNOR2_X1 port map( A => n1076, B => n1073, ZN => n1029);
   U1334 : XNOR2_X1 port map( A => n1074, B => n1029, ZN => n1033);
   U1335 : AOI22_X1 port map( A1 => n1348, A2 => OP2(21), B1 => n1330, B2 => 
                           OP1(21), ZN => n1032);
   U1336 : AOI22_X1 port map( A1 => n1244, A2 => n1030, B1 => n1242, B2 => 
                           n1285, ZN => n1031);
   U1337 : OAI211_X1 port map( C1 => n1033, C2 => n1284, A => n1032, B => n1031
                           , ZN => n1043);
   U1338 : NAND4_X1 port map( A1 => n1037, A2 => n1036, A3 => n1035, A4 => 
                           n1034, ZN => n1286);
   U1339 : AOI22_X1 port map( A1 => n1228, A2 => n1286, B1 => n1230, B2 => 
                           n1038, ZN => n1041);
   U1340 : AOI21_X1 port map( B1 => n1252, B2 => n1039, A => n1121, ZN => n1040
                           );
   U1341 : OAI211_X1 port map( C1 => n1051, C2 => n1368, A => n1041, B => n1040
                           , ZN => n1042);
   U1342 : AOI211_X1 port map( C1 => n1122, C2 => n1170, A => n1043, B => n1042
                           , ZN => n1044);
   U1343 : OAI211_X1 port map( C1 => n1398, C2 => n1046, A => n1045, B => n1044
                           , ZN => Y(21));
   U1344 : INV_X1 port map( A => n1125, ZN => n1056);
   U1345 : NAND2_X1 port map( A1 => n1049, A2 => n1047, ZN => n1054);
   U1346 : INV_X1 port map( A => n1048, ZN => n1053);
   U1347 : OAI21_X1 port map( B1 => n1051, B2 => n1050, A => n1049, ZN => n1052
                           );
   U1348 : OAI21_X1 port map( B1 => n1054, B2 => n1053, A => n1052, ZN => n1126
                           );
   U1349 : INV_X1 port map( A => n1126, ZN => n1055);
   U1350 : AOI221_X1 port map( B1 => n1056, B2 => n1055, C1 => n1125, C2 => 
                           n1126, A => n1398, ZN => n1072);
   U1351 : NOR2_X1 port map( A1 => OP_A_22_port, A2 => OP_B_22_port, ZN => 
                           n1104);
   U1352 : OAI22_X1 port map( A1 => n1104, A2 => n1368, B1 => n1124, B2 => 
                           n1369, ZN => n1071);
   U1353 : AOI22_X1 port map( A1 => n1348, A2 => OP2(22), B1 => n1330, B2 => 
                           OP1(22), ZN => n1068);
   U1354 : NAND4_X1 port map( A1 => n1060, A2 => n1059, A3 => n1058, A4 => 
                           n1057, ZN => n1317);
   U1355 : INV_X1 port map( A => n1317, ZN => n1184);
   U1356 : INV_X1 port map( A => n1207, ZN => n1061);
   U1357 : OAI22_X1 port map( A1 => n1184, A2 => n1062, B1 => n1061, B2 => 
                           n1233, ZN => n1065);
   U1358 : INV_X1 port map( A => n1242, ZN => n1183);
   U1359 : OAI22_X1 port map( A1 => n1210, A2 => n1183, B1 => n1063, B2 => 
                           n1211, ZN => n1064);
   U1360 : AOI211_X1 port map( C1 => n1252, C2 => n1066, A => n1065, B => n1064
                           , ZN => n1067);
   U1361 : OAI211_X1 port map( C1 => n1069, C2 => n1111, A => n1068, B => n1067
                           , ZN => n1070);
   U1362 : NOR4_X1 port map( A1 => n1121, A2 => n1072, A3 => n1071, A4 => n1070
                           , ZN => n1088);
   U1363 : NAND2_X1 port map( A1 => n1074, A2 => n1073, ZN => n1075);
   U1364 : AOI22_X1 port map( A1 => intadd_1_SUM_15_port, A2 => n1077, B1 => 
                           n1076, B2 => n1075, ZN => n1091);
   U1365 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n1079, A => n1078, ZN 
                           => n1080);
   U1366 : INV_X1 port map( A => n1080, ZN => n1092);
   U1367 : XNOR2_X1 port map( A => DP_OP_446J3_125_4819_n12, B => n1092, ZN => 
                           n1083);
   U1368 : AOI21_X1 port map( B1 => n1414, B2 => n1083, A => n1380, ZN => n1084
                           );
   U1369 : INV_X1 port map( A => n1084, ZN => n1090);
   U1370 : XNOR2_X1 port map( A => n1091, B => n1090, ZN => n1086);
   U1371 : AOI21_X1 port map( B1 => intadd_1_SUM_16_port, B2 => n1086, A => 
                           n1284, ZN => n1085);
   U1372 : OAI21_X1 port map( B1 => intadd_1_SUM_16_port, B2 => n1086, A => 
                           n1085, ZN => n1087);
   U1373 : OAI211_X1 port map( C1 => n1372, C2 => n1125, A => n1088, B => n1087
                           , ZN => Y(22));
   U1374 : INV_X1 port map( A => intadd_1_SUM_16_port, ZN => n1089);
   U1375 : FA_X1 port map( A => n1091, B => n1090, CI => n1089, CO => n1093, S 
                           => n_1170);
   U1376 : NOR3_X1 port map( A1 => n1093, A2 => n57, A3 => n1380, ZN => n1143);
   U1377 : INV_X1 port map( A => n1143, ZN => n1094);
   U1378 : OAI21_X1 port map( B1 => n1380, B2 => n57, A => n1093, ZN => n1144);
   U1379 : NAND2_X1 port map( A1 => n1094, A2 => n1144, ZN => n1095);
   U1380 : XNOR2_X1 port map( A => intadd_1_SUM_17_port, B => n1095, ZN => 
                           n1118);
   U1381 : NAND4_X1 port map( A1 => n1099, A2 => n1098, A3 => n1097, A4 => 
                           n1096, ZN => n1349);
   U1382 : AOI22_X1 port map( A1 => n1228, A2 => n1349, B1 => n1122, B2 => 
                           n1229, ZN => n1102);
   U1383 : AOI22_X1 port map( A1 => n1244, A2 => n1100, B1 => n1242, B2 => 
                           n1351, ZN => n1101);
   U1384 : OAI211_X1 port map( C1 => n1123, C2 => n1369, A => n1102, B => n1101
                           , ZN => n1103);
   U1385 : AOI21_X1 port map( B1 => n1344, B2 => n1106, A => n1103, ZN => n1117
                           );
   U1386 : OAI21_X1 port map( B1 => n1104, B2 => n1126, A => n1124, ZN => n1105
                           );
   U1387 : XOR2_X1 port map( A => n1106, B => n1105, Z => n1115);
   U1388 : OAI22_X1 port map( A1 => n1108, A2 => n1368, B1 => n1107, B2 => 
                           n1181, ZN => n1114);
   U1389 : AOI22_X1 port map( A1 => n1348, A2 => OP2(23), B1 => n1330, B2 => 
                           OP1(23), ZN => n1110);
   U1390 : OAI211_X1 port map( C1 => n1112, C2 => n1111, A => n1110, B => n1109
                           , ZN => n1113);
   U1391 : AOI211_X1 port map( C1 => n1115, C2 => N279, A => n1114, B => n1113,
                           ZN => n1116);
   U1392 : OAI211_X1 port map( C1 => n1284, C2 => n1118, A => n1117, B => n1116
                           , ZN => Y(23));
   U1393 : AOI22_X1 port map( A1 => n1242, A2 => n1269, B1 => n1230, B2 => 
                           n1119, ZN => n1152);
   U1394 : OAI22_X1 port map( A1 => n1193, A2 => n1369, B1 => n1129, B2 => 
                           n1372, ZN => n1120);
   U1395 : AOI211_X1 port map( C1 => n1122, C2 => n1268, A => n1121, B => n1120
                           , ZN => n1151);
   U1396 : OAI211_X1 port map( C1 => n1126, C2 => n1125, A => n1124, B => n1123
                           , ZN => n1127);
   U1397 : OAI21_X1 port map( B1 => OP_A_23_port, B2 => OP_B_23_port, A => 
                           n1127, ZN => n1192);
   U1398 : NOR2_X1 port map( A1 => n1192, A2 => n1129, ZN => n1128);
   U1399 : AOI211_X1 port map( C1 => n1192, C2 => n1129, A => n1398, B => n1128
                           , ZN => n1141);
   U1400 : NAND4_X1 port map( A1 => n1133, A2 => n1132, A3 => n1131, A4 => 
                           n1130, ZN => n1274);
   U1401 : AOI22_X1 port map( A1 => n1330, A2 => OP1(24), B1 => n1228, B2 => 
                           n1274, ZN => n1137);
   U1402 : AOI22_X1 port map( A1 => n1252, A2 => n1135, B1 => n1244, B2 => 
                           n1134, ZN => n1136);
   U1403 : OAI211_X1 port map( C1 => n1139, C2 => n1138, A => n1137, B => n1136
                           , ZN => n1140);
   U1404 : AOI211_X1 port map( C1 => n1367, C2 => n1142, A => n1141, B => n1140
                           , ZN => n1150);
   U1405 : AOI21_X1 port map( B1 => intadd_1_SUM_17_port, B2 => n1144, A => 
                           n1143, ZN => n1145);
   U1406 : NOR3_X1 port map( A1 => n1145, A2 => n57, A3 => n1380, ZN => n1153);
   U1407 : INV_X1 port map( A => n1153, ZN => n1146);
   U1408 : OAI21_X1 port map( B1 => n1380, B2 => n57, A => n1145, ZN => n1154);
   U1409 : NAND2_X1 port map( A1 => n1146, A2 => n1154, ZN => n1148);
   U1410 : AOI21_X1 port map( B1 => intadd_1_SUM_18_port, B2 => n1148, A => 
                           n1284, ZN => n1147);
   U1411 : OAI21_X1 port map( B1 => intadd_1_SUM_18_port, B2 => n1148, A => 
                           n1147, ZN => n1149);
   U1412 : NAND4_X1 port map( A1 => n1152, A2 => n1151, A3 => n1150, A4 => 
                           n1149, ZN => Y(24));
   U1413 : AOI21_X1 port map( B1 => intadd_1_SUM_18_port, B2 => n1154, A => 
                           n1153, ZN => n1155);
   U1414 : NOR3_X1 port map( A1 => n1155, A2 => n57, A3 => n1380, ZN => n1186);
   U1415 : INV_X1 port map( A => n1186, ZN => n1156);
   U1416 : OAI21_X1 port map( B1 => n1380, B2 => n57, A => n1155, ZN => n1187);
   U1417 : NAND2_X1 port map( A1 => n1156, A2 => n1187, ZN => n1157);
   U1418 : XNOR2_X1 port map( A => intadd_1_SUM_19_port, B => n1157, ZN => 
                           n1180);
   U1419 : AOI211_X1 port map( C1 => n1160, C2 => n1363, A => n1159, B => n1158
                           , ZN => n1236);
   U1420 : AOI22_X1 port map( A1 => n1244, A2 => n1161, B1 => n1242, B2 => 
                           n1286, ZN => n1162);
   U1421 : OAI21_X1 port map( B1 => n1194, B2 => n1369, A => n1162, ZN => n1163
                           );
   U1422 : AOI211_X1 port map( C1 => n1165, C2 => n1344, A => n1236, B => n1163
                           , ZN => n1179);
   U1423 : AOI21_X1 port map( B1 => n1192, B2 => n1193, A => n1195, ZN => n1164
                           );
   U1424 : XOR2_X1 port map( A => n1165, B => n1164, Z => n1177);
   U1425 : INV_X1 port map( A => n1285, ZN => n1173);
   U1426 : NAND4_X1 port map( A1 => n1169, A2 => n1168, A3 => n1167, A4 => 
                           n1166, ZN => n1291);
   U1427 : AOI22_X1 port map( A1 => n1230, A2 => n1170, B1 => n1228, B2 => 
                           n1291, ZN => n1172);
   U1428 : AOI22_X1 port map( A1 => n1348, A2 => OP2(25), B1 => n1330, B2 => 
                           OP1(25), ZN => n1171);
   U1429 : OAI211_X1 port map( C1 => n1173, C2 => n1233, A => n1172, B => n1171
                           , ZN => n1176);
   U1430 : OAI22_X1 port map( A1 => n1196, A2 => n1368, B1 => n1174, B2 => 
                           n1181, ZN => n1175);
   U1431 : AOI211_X1 port map( C1 => n1177, C2 => N279, A => n1176, B => n1175,
                           ZN => n1178);
   U1432 : OAI211_X1 port map( C1 => n1284, C2 => n1180, A => n1179, B => n1178
                           , ZN => Y(25));
   U1433 : INV_X1 port map( A => n1200, ZN => n1202);
   U1434 : OAI22_X1 port map( A1 => n1184, A2 => n1183, B1 => n1182, B2 => 
                           n1181, ZN => n1185);
   U1435 : AOI211_X1 port map( C1 => n1202, C2 => n1344, A => n1236, B => n1185
                           , ZN => n1218);
   U1436 : AOI21_X1 port map( B1 => intadd_1_SUM_19_port, B2 => n1187, A => 
                           n1186, ZN => n1188);
   U1437 : NOR3_X1 port map( A1 => n1188, A2 => n57, A3 => n1380, ZN => n1219);
   U1438 : INV_X1 port map( A => n1219, ZN => n1189);
   U1439 : OAI21_X1 port map( B1 => n1380, B2 => n57, A => n1188, ZN => n1220);
   U1440 : NAND2_X1 port map( A1 => n1189, A2 => n1220, ZN => n1191);
   U1441 : NOR2_X1 port map( A1 => intadd_1_SUM_20_port, A2 => n1191, ZN => 
                           n1190);
   U1442 : AOI211_X1 port map( C1 => intadd_1_SUM_20_port, C2 => n1191, A => 
                           n1284, B => n1190, ZN => n1216);
   U1443 : INV_X1 port map( A => n1192, ZN => n1199);
   U1444 : NAND2_X1 port map( A1 => n1194, A2 => n1193, ZN => n1198);
   U1445 : OAI21_X1 port map( B1 => n1196, B2 => n1195, A => n1194, ZN => n1197
                           );
   U1446 : OAI21_X1 port map( B1 => n1199, B2 => n1198, A => n1197, ZN => n1238
                           );
   U1447 : INV_X1 port map( A => n1238, ZN => n1201);
   U1448 : AOI221_X1 port map( B1 => n1202, B2 => n1201, C1 => n1200, C2 => 
                           n1238, A => n1398, ZN => n1215);
   U1449 : NAND4_X1 port map( A1 => n1206, A2 => n1205, A3 => n1204, A4 => 
                           n1203, ZN => n1322);
   U1450 : AOI22_X1 port map( A1 => n1230, A2 => n1207, B1 => n1228, B2 => 
                           n1322, ZN => n1209);
   U1451 : AOI22_X1 port map( A1 => n1348, A2 => OP2(26), B1 => n1330, B2 => 
                           OP1(26), ZN => n1208);
   U1452 : OAI211_X1 port map( C1 => n1210, C2 => n1233, A => n1209, B => n1208
                           , ZN => n1214);
   U1453 : NOR2_X1 port map( A1 => OP_A_26_port, A2 => OP_B_26_port, ZN => 
                           n1239);
   U1454 : OAI22_X1 port map( A1 => n1239, A2 => n1368, B1 => n1212, B2 => 
                           n1211, ZN => n1213);
   U1455 : NOR4_X1 port map( A1 => n1216, A2 => n1215, A3 => n1214, A4 => n1213
                           , ZN => n1217);
   U1456 : OAI211_X1 port map( C1 => n1237, C2 => n1369, A => n1218, B => n1217
                           , ZN => Y(26));
   U1457 : AOI21_X1 port map( B1 => intadd_1_SUM_20_port, B2 => n1220, A => 
                           n1219, ZN => n1221);
   U1458 : NOR3_X1 port map( A1 => n1221, A2 => n57, A3 => n1380, ZN => n1256);
   U1459 : INV_X1 port map( A => n1256, ZN => n1222);
   U1460 : OAI21_X1 port map( B1 => n1380, B2 => n57, A => n1221, ZN => n1257);
   U1461 : NAND2_X1 port map( A1 => n1222, A2 => n1257, ZN => n1223);
   U1462 : XNOR2_X1 port map( A => intadd_1_SUM_21_port, B => n1223, ZN => 
                           n1255);
   U1463 : INV_X1 port map( A => n1351, ZN => n1234);
   U1464 : NAND4_X1 port map( A1 => n1227, A2 => n1226, A3 => n1225, A4 => 
                           n1224, ZN => n1357);
   U1465 : AOI22_X1 port map( A1 => n1230, A2 => n1229, B1 => n1228, B2 => 
                           n1357, ZN => n1232);
   U1466 : AOI22_X1 port map( A1 => n1348, A2 => OP2(27), B1 => n1330, B2 => 
                           OP1(27), ZN => n1231);
   U1467 : OAI211_X1 port map( C1 => n1234, C2 => n1233, A => n1232, B => n1231
                           , ZN => n1235);
   U1468 : AOI211_X1 port map( C1 => n1344, C2 => n1241, A => n1236, B => n1235
                           , ZN => n1254);
   U1469 : OAI21_X1 port map( B1 => n1239, B2 => n1238, A => n1237, ZN => n1266
                           );
   U1470 : OAI21_X1 port map( B1 => n1241, B2 => n1266, A => N279, ZN => n1240)
                           ;
   U1471 : AOI21_X1 port map( B1 => n1241, B2 => n1266, A => n1240, ZN => n1250
                           );
   U1472 : AOI22_X1 port map( A1 => n1244, A2 => n1243, B1 => n1242, B2 => 
                           n1349, ZN => n1247);
   U1473 : OAI221_X1 port map( B1 => n1367, B2 => n1245, C1 => n1367, C2 => 
                           OP_A_27_port, A => OP_B_27_port, ZN => n1246);
   U1474 : OAI211_X1 port map( C1 => n1368, C2 => n1248, A => n1247, B => n1246
                           , ZN => n1249);
   U1475 : AOI211_X1 port map( C1 => n1252, C2 => n1251, A => n1250, B => n1249
                           , ZN => n1253);
   U1476 : OAI211_X1 port map( C1 => n1284, C2 => n1255, A => n1254, B => n1253
                           , ZN => Y(27));
   U1477 : AOI21_X1 port map( B1 => intadd_1_SUM_21_port, B2 => n1257, A => 
                           n1256, ZN => n1258);
   U1478 : NOR3_X1 port map( A1 => n1258, A2 => n57, A3 => n1380, ZN => n1303);
   U1479 : INV_X1 port map( A => n1303, ZN => n1259);
   U1480 : OAI21_X1 port map( B1 => n1380, B2 => n57, A => n1258, ZN => n1304);
   U1481 : NAND2_X1 port map( A1 => n1259, A2 => n1304, ZN => n1260);
   U1482 : XNOR2_X1 port map( A => intadd_1_SUM_22_port, B => n1260, ZN => 
                           n1283);
   U1483 : AOI22_X1 port map( A1 => n1348, A2 => OP2(28), B1 => n1330, B2 => 
                           OP1(28), ZN => n1262);
   U1484 : NAND3_X1 port map( A1 => OP_SHIFT, A2 => N284, A3 => n1261, ZN => 
                           n1402);
   U1485 : OAI211_X1 port map( C1 => n1299, C2 => n1368, A => n1262, B => n1402
                           , ZN => n1264);
   U1486 : OAI22_X1 port map( A1 => n1301, A2 => n1369, B1 => n1372, B2 => 
                           n1267, ZN => n1263);
   U1487 : AOI211_X1 port map( C1 => n1329, C2 => n1265, A => n1264, B => n1263
                           , ZN => n1282);
   U1488 : AOI222_X1 port map( A1 => OP_A_27_port, A2 => OP_B_27_port, B1 => 
                           OP_A_27_port, B2 => n1266, C1 => OP_B_27_port, C2 =>
                           n1266, ZN => n1300);
   U1489 : XOR2_X1 port map( A => n1267, B => n1300, Z => n1280);
   U1490 : AOI22_X1 port map( A1 => n1350, A2 => n1269, B1 => n1352, B2 => 
                           n1268, ZN => n1277);
   U1491 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n56, ZN => n1273);
   U1492 : NAND4_X1 port map( A1 => n1273, A2 => n1272, A3 => n1271, A4 => 
                           n1270, ZN => n1275);
   U1493 : AOI22_X1 port map( A1 => n1360, A2 => n1275, B1 => n1358, B2 => 
                           n1274, ZN => n1276);
   U1494 : OAI211_X1 port map( C1 => n1278, C2 => n1363, A => n1277, B => n1276
                           , ZN => n1279);
   U1495 : AOI22_X1 port map( A1 => n1280, A2 => N279, B1 => n1366, B2 => n1279
                           , ZN => n1281);
   U1496 : OAI211_X1 port map( C1 => n1284, C2 => n1283, A => n1282, B => n1281
                           , ZN => Y(28));
   U1497 : AOI22_X1 port map( A1 => n1348, A2 => OP2(29), B1 => n1330, B2 => 
                           OP1(29), ZN => n1315);
   U1498 : AOI22_X1 port map( A1 => n1350, A2 => n1286, B1 => n1352, B2 => 
                           n1285, ZN => n1294);
   U1499 : NAND4_X1 port map( A1 => n1290, A2 => n1289, A3 => n1288, A4 => 
                           n1287, ZN => n1292);
   U1500 : AOI22_X1 port map( A1 => n1360, A2 => n1292, B1 => n1358, B2 => 
                           n1291, ZN => n1293);
   U1501 : OAI211_X1 port map( C1 => n1295, C2 => n1363, A => n1294, B => n1293
                           , ZN => n1296);
   U1502 : AOI22_X1 port map( A1 => OP_A_29_port, A2 => n1367, B1 => n1366, B2 
                           => n1296, ZN => n1314);
   U1503 : OAI21_X1 port map( B1 => n1297, B2 => n1369, A => n1368, ZN => n1312
                           );
   U1504 : OAI22_X1 port map( A1 => n1302, A2 => n1372, B1 => n1298, B2 => 
                           n1373, ZN => n1311);
   U1505 : AOI21_X1 port map( B1 => n1301, B2 => n1300, A => n1299, ZN => n1332
                           );
   U1506 : XOR2_X1 port map( A => n1332, B => n1302, Z => n1309);
   U1507 : AOI21_X1 port map( B1 => intadd_1_SUM_22_port, B2 => n1304, A => 
                           n1303, ZN => n1305);
   U1508 : NOR3_X1 port map( A1 => n1305, A2 => n57, A3 => n1380, ZN => n1334);
   U1509 : INV_X1 port map( A => n1334, ZN => n1306);
   U1510 : OAI21_X1 port map( B1 => n1380, B2 => n57, A => n1305, ZN => n1335);
   U1511 : NAND2_X1 port map( A1 => n1306, A2 => n1335, ZN => n1307);
   U1512 : XNOR2_X1 port map( A => intadd_1_SUM_23_port, B => n1307, ZN => 
                           n1308);
   U1513 : OAI22_X1 port map( A1 => n1398, A2 => n1309, B1 => n1396, B2 => 
                           n1308, ZN => n1310);
   U1514 : AOI211_X1 port map( C1 => OP_B_29_port, C2 => n1312, A => n1311, B 
                           => n1310, ZN => n1313);
   U1515 : NAND4_X1 port map( A1 => n1315, A2 => n1314, A3 => n1313, A4 => 
                           n1402, ZN => Y(29));
   U1516 : AOI22_X1 port map( A1 => n1350, A2 => n1317, B1 => n1352, B2 => 
                           n1316, ZN => n1325);
   U1517 : NAND2_X1 port map( A1 => OP_A_30_port, A2 => n56, ZN => n1321);
   U1518 : NAND4_X1 port map( A1 => n1321, A2 => n1320, A3 => n1319, A4 => 
                           n1318, ZN => n1323);
   U1519 : AOI22_X1 port map( A1 => n1360, A2 => n1323, B1 => n1358, B2 => 
                           n1322, ZN => n1324);
   U1520 : OAI211_X1 port map( C1 => n1326, C2 => n1363, A => n1325, B => n1324
                           , ZN => n1327);
   U1521 : AOI22_X1 port map( A1 => n1329, A2 => n1328, B1 => n1366, B2 => 
                           n1327, ZN => n1346);
   U1522 : AOI22_X1 port map( A1 => n1348, A2 => OP2(30), B1 => n1330, B2 => 
                           OP1(30), ZN => n1331);
   U1523 : OAI211_X1 port map( C1 => n1375, C2 => n1368, A => n1331, B => n1402
                           , ZN => n1342);
   U1524 : AOI222_X1 port map( A1 => OP_B_29_port, A2 => OP_A_29_port, B1 => 
                           OP_B_29_port, B2 => n1332, C1 => OP_A_29_port, C2 =>
                           n1332, ZN => n1376);
   U1525 : XNOR2_X1 port map( A => n1376, B => n1333, ZN => n1340);
   U1526 : AOI21_X1 port map( B1 => intadd_1_SUM_23_port, B2 => n1335, A => 
                           n1334, ZN => n1336);
   U1527 : NOR3_X1 port map( A1 => n1336, A2 => n57, A3 => n1380, ZN => n1386);
   U1528 : INV_X1 port map( A => n1386, ZN => n1337);
   U1529 : OAI21_X1 port map( B1 => n1380, B2 => n57, A => n1336, ZN => n1387);
   U1530 : NAND2_X1 port map( A1 => n1337, A2 => n1387, ZN => n1338);
   U1531 : XNOR2_X1 port map( A => intadd_1_SUM_24_port, B => n1338, ZN => 
                           n1339);
   U1532 : OAI22_X1 port map( A1 => n1398, A2 => n1340, B1 => n1396, B2 => 
                           n1339, ZN => n1341);
   U1533 : AOI211_X1 port map( C1 => n1344, C2 => n1343, A => n1342, B => n1341
                           , ZN => n1345);
   U1534 : OAI211_X1 port map( C1 => n1377, C2 => n1369, A => n1346, B => n1345
                           , ZN => Y(30));
   U1535 : AOI22_X1 port map( A1 => n1348, A2 => OP2(31), B1 => OP1(31), B2 => 
                           n1347, ZN => n1405);
   U1536 : AOI22_X1 port map( A1 => n1352, A2 => n1351, B1 => n1350, B2 => 
                           n1349, ZN => n1362);
   U1537 : NAND2_X1 port map( A1 => OP_A_31_port, A2 => n56, ZN => n1356);
   U1538 : NAND4_X1 port map( A1 => n1356, A2 => n1355, A3 => n1354, A4 => 
                           n1353, ZN => n1359);
   U1539 : AOI22_X1 port map( A1 => n1360, A2 => n1359, B1 => n1358, B2 => 
                           n1357, ZN => n1361);
   U1540 : OAI211_X1 port map( C1 => n1364, C2 => n1363, A => n1362, B => n1361
                           , ZN => n1365);
   U1541 : AOI22_X1 port map( A1 => OP_A_31_port, A2 => n1367, B1 => n1366, B2 
                           => n1365, ZN => n1404);
   U1542 : OAI21_X1 port map( B1 => n1370, B2 => n1369, A => n1368, ZN => n1401
                           );
   U1543 : INV_X1 port map( A => n1371, ZN => n1378);
   U1544 : OAI22_X1 port map( A1 => n1374, A2 => n1373, B1 => n1378, B2 => 
                           n1372, ZN => n1400);
   U1545 : AOI21_X1 port map( B1 => n1377, B2 => n1376, A => n1375, ZN => n1379
                           );
   U1546 : XOR2_X1 port map( A => n1379, B => n1378, Z => n1397);
   U1547 : NOR2_X1 port map( A1 => n57, A2 => n1380, ZN => n1385);
   U1548 : INV_X1 port map( A => n1381, ZN => n1382);
   U1549 : AOI21_X1 port map( B1 => n1383, B2 => n1382, A => n1385, ZN => n1384
                           );
   U1550 : AOI21_X1 port map( B1 => n1385, B2 => intadd_1_B_18_port, A => n1384
                           , ZN => n1389);
   U1551 : AOI21_X1 port map( B1 => intadd_1_SUM_24_port, B2 => n1387, A => 
                           n1386, ZN => n1388);
   U1552 : XOR2_X1 port map( A => n1389, B => n1388, Z => n1390);
   U1553 : MUX2_X1 port map( A => n62, B => n58, S => n1390, Z => n1394);
   U1554 : INV_X1 port map( A => intadd_0_A_16_port, ZN => n1391);
   U1555 : MUX2_X1 port map( A => intadd_0_A_16_port, B => n1391, S => 
                           intadd_0_n1, Z => n1392);
   U1556 : XOR2_X1 port map( A => intadd_1_n1, B => n1392, Z => n1393);
   U1557 : XNOR2_X1 port map( A => n1394, B => n1393, ZN => n1395);
   U1558 : OAI22_X1 port map( A1 => n1398, A2 => n1397, B1 => n1396, B2 => 
                           n1395, ZN => n1399);
   U1559 : AOI211_X1 port map( C1 => OP_B_31_port, C2 => n1401, A => n1400, B 
                           => n1399, ZN => n1403);
   U1560 : NAND4_X1 port map( A1 => n1405, A2 => n1404, A3 => n1403, A4 => 
                           n1402, ZN => Y(31));
   U1561 : OAI22_X1 port map( A1 => OPC(6), A2 => n1407, B1 => n1406, B2 => 
                           n1411, ZN => N282);
   U1562 : OAI22_X1 port map( A1 => n1411, A2 => n1410, B1 => n1409, B2 => 
                           n1408, ZN => N283);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( CLK, RST : in std_logic);

end DLX;

architecture SYN_DLX_RTL of DLX is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component RF_N32_NA5
      port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
            ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component ALU_N32_NB8
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
            std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);
            Z : out std_logic);
   end component;
   
   component DLX_DRAM_N256_NW32
      port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector 
            (31 downto 0);  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component DLX_IRAM_RAM_DEPTH256_I_SIZE32
      port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  
            DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, 
      IR_26_port, IR_10_port, IR_9_port, IR_8_port, IR_7_port, IR_6_port, 
      IR_5_port, IR_4_port, IR_3_port, IR_2_port, IR_1_port, IR_0_port, 
      ALU_OPCODE_i_0_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_4_port, ALU_OPCODE_i_5_port, 
      ALU_OPCODE_i_6_port, IR_BUS_31_port, IR_BUS_30_port, IR_BUS_29_port, 
      IR_BUS_28_port, IR_BUS_27_port, IR_BUS_26_port, IR_BUS_25_port, 
      IR_BUS_24_port, IR_BUS_23_port, IR_BUS_22_port, IR_BUS_21_port, 
      IR_BUS_20_port, IR_BUS_19_port, IR_BUS_18_port, IR_BUS_17_port, 
      IR_BUS_16_port, IR_BUS_15_port, IR_BUS_14_port, IR_BUS_13_port, 
      IR_BUS_12_port, IR_BUS_11_port, IR_BUS_10_port, IR_BUS_9_port, 
      IR_BUS_8_port, IR_BUS_7_port, IR_BUS_6_port, IR_BUS_5_port, IR_BUS_4_port
      , IR_BUS_3_port, IR_BUS_2_port, IR_BUS_1_port, IR_BUS_0_port, 
      DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, DATA_OUT_28_port, 
      DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, DATA_OUT_24_port, 
      DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, 
      DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, 
      DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, 
      DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, 
      DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, 
      DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port, 
      DATA_ADDR_31_port, DATA_ADDR_30_port, DATA_ADDR_29_port, 
      DATA_ADDR_28_port, DATA_ADDR_27_port, DATA_ADDR_26_port, 
      DATA_ADDR_25_port, DATA_ADDR_24_port, DATA_ADDR_23_port, 
      DATA_ADDR_22_port, DATA_ADDR_21_port, DATA_ADDR_20_port, 
      DATA_ADDR_19_port, DATA_ADDR_18_port, DATA_ADDR_17_port, 
      DATA_ADDR_16_port, DATA_ADDR_15_port, DATA_ADDR_14_port, 
      DATA_ADDR_13_port, DATA_ADDR_12_port, DATA_ADDR_11_port, 
      DATA_ADDR_10_port, DATA_ADDR_9_port, DATA_ADDR_8_port, DATA_ADDR_7_port, 
      DATA_ADDR_6_port, DATA_ADDR_5_port, DATA_ADDR_4_port, DATA_ADDR_3_port, 
      DATA_ADDR_2_port, DATA_ADDR_1_port, DATA_ADDR_0_port, DATA_IN_31_port, 
      DATA_IN_30_port, DATA_IN_29_port, DATA_IN_28_port, DATA_IN_27_port, 
      DATA_IN_26_port, DATA_IN_25_port, DATA_IN_24_port, DATA_IN_23_port, 
      DATA_IN_22_port, DATA_IN_21_port, DATA_IN_20_port, DATA_IN_19_port, 
      DATA_IN_18_port, DATA_IN_17_port, DATA_IN_16_port, DATA_IN_15_port, 
      DATA_IN_14_port, DATA_IN_13_port, DATA_IN_12_port, DATA_IN_11_port, 
      DATA_IN_10_port, DATA_IN_9_port, DATA_IN_8_port, DATA_IN_7_port, 
      DATA_IN_6_port, DATA_IN_5_port, DATA_IN_4_port, DATA_IN_3_port, 
      DATA_IN_2_port, DATA_IN_1_port, DATA_IN_0_port, CU_I_aluOpcode2_0_port, 
      CU_I_aluOpcode2_1_port, CU_I_aluOpcode2_2_port, CU_I_aluOpcode2_3_port, 
      CU_I_aluOpcode2_4_port, CU_I_aluOpcode2_5_port, CU_I_aluOpcode2_6_port, 
      CU_I_aluOpcode1_0_port, CU_I_aluOpcode1_1_port, CU_I_aluOpcode1_2_port, 
      CU_I_aluOpcode1_3_port, CU_I_aluOpcode1_4_port, CU_I_aluOpcode1_5_port, 
      CU_I_aluOpcode1_6_port, DATAPATH_I_ALU_OUTPUT_0_port, 
      DATAPATH_I_ALU_OUTPUT_1_port, DATAPATH_I_ALU_OUTPUT_2_port, 
      DATAPATH_I_ALU_OUTPUT_3_port, DATAPATH_I_ALU_OUTPUT_4_port, 
      DATAPATH_I_ALU_OUTPUT_5_port, DATAPATH_I_ALU_OUTPUT_6_port, 
      DATAPATH_I_ALU_OUTPUT_7_port, DATAPATH_I_ALU_OUTPUT_8_port, 
      DATAPATH_I_ALU_OUTPUT_9_port, DATAPATH_I_ALU_OUTPUT_10_port, 
      DATAPATH_I_ALU_OUTPUT_11_port, DATAPATH_I_ALU_OUTPUT_12_port, 
      DATAPATH_I_ALU_OUTPUT_13_port, DATAPATH_I_ALU_OUTPUT_14_port, 
      DATAPATH_I_ALU_OUTPUT_15_port, DATAPATH_I_ALU_OUTPUT_16_port, 
      DATAPATH_I_ALU_OUTPUT_17_port, DATAPATH_I_ALU_OUTPUT_18_port, 
      DATAPATH_I_ALU_OUTPUT_19_port, DATAPATH_I_ALU_OUTPUT_20_port, 
      DATAPATH_I_ALU_OUTPUT_21_port, DATAPATH_I_ALU_OUTPUT_22_port, 
      DATAPATH_I_ALU_OUTPUT_23_port, DATAPATH_I_ALU_OUTPUT_24_port, 
      DATAPATH_I_ALU_OUTPUT_25_port, DATAPATH_I_ALU_OUTPUT_26_port, 
      DATAPATH_I_ALU_OUTPUT_27_port, DATAPATH_I_ALU_OUTPUT_28_port, 
      DATAPATH_I_ALU_OUTPUT_29_port, DATAPATH_I_ALU_OUTPUT_30_port, 
      DATAPATH_I_ALU_OUTPUT_31_port, DATAPATH_I_RF_OUT2_0_port, 
      DATAPATH_I_RF_OUT2_1_port, DATAPATH_I_RF_OUT2_2_port, 
      DATAPATH_I_RF_OUT2_3_port, DATAPATH_I_RF_OUT2_4_port, 
      DATAPATH_I_RF_OUT2_5_port, DATAPATH_I_RF_OUT2_6_port, 
      DATAPATH_I_RF_OUT2_7_port, DATAPATH_I_RF_OUT2_8_port, 
      DATAPATH_I_RF_OUT2_9_port, DATAPATH_I_RF_OUT2_10_port, 
      DATAPATH_I_RF_OUT2_11_port, DATAPATH_I_RF_OUT2_12_port, 
      DATAPATH_I_RF_OUT2_13_port, DATAPATH_I_RF_OUT2_14_port, 
      DATAPATH_I_RF_OUT2_15_port, DATAPATH_I_RF_OUT2_16_port, 
      DATAPATH_I_RF_OUT2_17_port, DATAPATH_I_RF_OUT2_18_port, 
      DATAPATH_I_RF_OUT2_19_port, DATAPATH_I_RF_OUT2_20_port, 
      DATAPATH_I_RF_OUT2_21_port, DATAPATH_I_RF_OUT2_22_port, 
      DATAPATH_I_RF_OUT2_23_port, DATAPATH_I_RF_OUT2_24_port, 
      DATAPATH_I_RF_OUT2_25_port, DATAPATH_I_RF_OUT2_26_port, 
      DATAPATH_I_RF_OUT2_27_port, DATAPATH_I_RF_OUT2_28_port, 
      DATAPATH_I_RF_OUT2_29_port, DATAPATH_I_RF_OUT2_30_port, 
      DATAPATH_I_RF_OUT2_31_port, DATAPATH_I_RF_OUT1_0_port, 
      DATAPATH_I_RF_OUT1_1_port, DATAPATH_I_RF_OUT1_2_port, 
      DATAPATH_I_RF_OUT1_3_port, DATAPATH_I_RF_OUT1_4_port, 
      DATAPATH_I_RF_OUT1_5_port, DATAPATH_I_RF_OUT1_6_port, 
      DATAPATH_I_RF_OUT1_7_port, DATAPATH_I_RF_OUT1_8_port, 
      DATAPATH_I_RF_OUT1_9_port, DATAPATH_I_RF_OUT1_10_port, 
      DATAPATH_I_RF_OUT1_11_port, DATAPATH_I_RF_OUT1_12_port, 
      DATAPATH_I_RF_OUT1_13_port, DATAPATH_I_RF_OUT1_14_port, 
      DATAPATH_I_RF_OUT1_15_port, DATAPATH_I_RF_OUT1_16_port, 
      DATAPATH_I_RF_OUT1_17_port, DATAPATH_I_RF_OUT1_18_port, 
      DATAPATH_I_RF_OUT1_19_port, DATAPATH_I_RF_OUT1_20_port, 
      DATAPATH_I_RF_OUT1_21_port, DATAPATH_I_RF_OUT1_22_port, 
      DATAPATH_I_RF_OUT1_23_port, DATAPATH_I_RF_OUT1_24_port, 
      DATAPATH_I_RF_OUT1_25_port, DATAPATH_I_RF_OUT1_26_port, 
      DATAPATH_I_RF_OUT1_27_port, DATAPATH_I_RF_OUT1_28_port, 
      DATAPATH_I_RF_OUT1_29_port, DATAPATH_I_RF_OUT1_30_port, 
      DATAPATH_I_RF_OUT1_31_port, DATAPATH_I_N414, DATAPATH_I_N413, 
      DATAPATH_I_N412, DATAPATH_I_N411, DATAPATH_I_N410, DATAPATH_I_N409, 
      DATAPATH_I_N408, DATAPATH_I_N407, DATAPATH_I_N406, DATAPATH_I_N405, 
      DATAPATH_I_N404, DATAPATH_I_N403, DATAPATH_I_N402, DATAPATH_I_N401, 
      DATAPATH_I_N400, DATAPATH_I_N399, DATAPATH_I_N398, DATAPATH_I_N397, 
      DATAPATH_I_N396, DATAPATH_I_N395, DATAPATH_I_N394, DATAPATH_I_N393, 
      DATAPATH_I_N392, DATAPATH_I_N391, DATAPATH_I_N390, DATAPATH_I_N389, 
      DATAPATH_I_N388, DATAPATH_I_N387, DATAPATH_I_N386, DATAPATH_I_N385, 
      DATAPATH_I_N384, DATAPATH_I_N383, DATAPATH_I_N382, DATAPATH_I_N381, 
      DATAPATH_I_N380, DATAPATH_I_N379, DATAPATH_I_N378, DATAPATH_I_N312, 
      DATAPATH_I_N311, DATAPATH_I_N310, DATAPATH_I_N309, DATAPATH_I_N308, 
      DATAPATH_I_N306, DATAPATH_I_N305, DATAPATH_I_N304, DATAPATH_I_N303, 
      DATAPATH_I_N302, DATAPATH_I_N301, DATAPATH_I_N300, DATAPATH_I_N299, 
      DATAPATH_I_N298, DATAPATH_I_N297, DATAPATH_I_N296, DATAPATH_I_N295, 
      DATAPATH_I_N294, DATAPATH_I_N293, DATAPATH_I_N292, DATAPATH_I_N291, 
      DATAPATH_I_N290, DATAPATH_I_N289, DATAPATH_I_N288, DATAPATH_I_N287, 
      DATAPATH_I_N286, DATAPATH_I_N285, DATAPATH_I_N284, DATAPATH_I_N283, 
      DATAPATH_I_N282, DATAPATH_I_N281, DATAPATH_I_N280, DATAPATH_I_N279, 
      DATAPATH_I_N278, DATAPATH_I_N277, DATAPATH_I_N276, DATAPATH_I_N275, 
      DATAPATH_I_N274, DATAPATH_I_N273, DATAPATH_I_N272, DATAPATH_I_N271, 
      DATAPATH_I_N270, DATAPATH_I_N269, DATAPATH_I_N268, DATAPATH_I_N267, 
      DATAPATH_I_N266, DATAPATH_I_N265, DATAPATH_I_N264, DATAPATH_I_N263, 
      DATAPATH_I_N262, DATAPATH_I_N261, DATAPATH_I_N260, DATAPATH_I_N259, 
      DATAPATH_I_N258, DATAPATH_I_N257, DATAPATH_I_N256, DATAPATH_I_N255, 
      DATAPATH_I_N254, DATAPATH_I_N253, DATAPATH_I_N252, DATAPATH_I_N251, 
      DATAPATH_I_N250, DATAPATH_I_N249, DATAPATH_I_N248, DATAPATH_I_N247, 
      DATAPATH_I_N246, DATAPATH_I_N245, DATAPATH_I_N244, DATAPATH_I_N243, 
      DATAPATH_I_N177, DATAPATH_I_N176, DATAPATH_I_N175, DATAPATH_I_N174, 
      DATAPATH_I_N173, DATAPATH_I_N172, DATAPATH_I_N171, DATAPATH_I_N170, 
      DATAPATH_I_N169, DATAPATH_I_N168, DATAPATH_I_N167, DATAPATH_I_N166, 
      DATAPATH_I_N165, DATAPATH_I_N164, DATAPATH_I_N163, DATAPATH_I_N162, 
      DATAPATH_I_N161, DATAPATH_I_N160, DATAPATH_I_N159, DATAPATH_I_N158, 
      DATAPATH_I_N157, DATAPATH_I_N156, DATAPATH_I_N155, DATAPATH_I_N154, 
      DATAPATH_I_N153, DATAPATH_I_N152, DATAPATH_I_N151, DATAPATH_I_N150, 
      DATAPATH_I_N149, DATAPATH_I_N148, DATAPATH_I_N147, DATAPATH_I_N146, 
      DATAPATH_I_N145, DATAPATH_I_N144, DATAPATH_I_N143, DATAPATH_I_N142, 
      DATAPATH_I_N141, DATAPATH_I_N140, DATAPATH_I_N139, DATAPATH_I_N138, 
      DATAPATH_I_N137, DATAPATH_I_N136, DATAPATH_I_N135, DATAPATH_I_N134, 
      DATAPATH_I_N133, DATAPATH_I_N132, DATAPATH_I_N131, DATAPATH_I_N130, 
      DATAPATH_I_N129, DATAPATH_I_N128, DATAPATH_I_N127, DATAPATH_I_N126, 
      DATAPATH_I_N125, DATAPATH_I_N124, DATAPATH_I_N123, DATAPATH_I_N122, 
      DATAPATH_I_N121, DATAPATH_I_N120, DATAPATH_I_N119, DATAPATH_I_N118, 
      DATAPATH_I_N117, DATAPATH_I_N116, DATAPATH_I_N115, DATAPATH_I_N114, 
      DATAPATH_I_N113, DATAPATH_I_N112, DATAPATH_I_N111, DATAPATH_I_N110, 
      DATAPATH_I_N109, DATAPATH_I_N65, DATAPATH_I_N64, DATAPATH_I_N63, 
      DATAPATH_I_N62, DATAPATH_I_N61, DATAPATH_I_N60, DATAPATH_I_N59, 
      DATAPATH_I_N58, DATAPATH_I_N57, DATAPATH_I_N56, DATAPATH_I_N55, 
      DATAPATH_I_N54, DATAPATH_I_N53, DATAPATH_I_N52, DATAPATH_I_N51, 
      DATAPATH_I_N50, DATAPATH_I_N49, DATAPATH_I_N48, DATAPATH_I_N47, 
      DATAPATH_I_N46, DATAPATH_I_N45, DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_0_port
      , DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_1_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_2_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_3_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_4_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_5_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_6_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_7_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_8_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_9_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_10_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_11_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_12_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_13_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_14_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_15_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_16_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_17_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_18_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_19_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_20_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_21_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_22_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_23_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_24_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_25_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_26_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_27_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_28_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_29_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_30_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_31_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_0_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_1_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_2_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_3_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_4_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_5_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_6_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_7_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_8_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_9_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_10_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_11_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_12_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_13_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_14_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_15_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_16_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_17_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_18_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_19_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_20_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_21_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_22_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_23_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_24_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_25_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_26_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_27_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_28_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_29_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_30_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_31_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_0_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_1_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_2_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_3_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_4_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_5_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_6_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_7_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_8_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_9_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_10_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_11_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_12_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_13_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_14_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_15_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_16_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_17_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_18_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_19_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_20_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_21_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_22_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_23_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_24_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_25_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_26_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_27_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_28_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_29_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_30_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_31_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_0_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_1_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_2_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_3_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_4_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_5_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_6_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_7_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_8_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_9_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_10_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_11_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_12_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_13_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_14_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_15_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_16_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_17_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_18_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_19_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_20_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_21_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_22_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_23_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_24_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_25_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_26_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_27_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_28_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_29_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_30_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_31_port, DATAPATH_I_ID_EX_RS2_NEXT_0_port, 
      DATAPATH_I_ID_EX_RS2_NEXT_1_port, DATAPATH_I_ID_EX_RS2_NEXT_2_port, 
      DATAPATH_I_ID_EX_RS2_NEXT_3_port, DATAPATH_I_ID_EX_RS2_NEXT_4_port, 
      DATAPATH_I_ID_EX_RS1_NEXT_0_port, DATAPATH_I_ID_EX_RS1_NEXT_1_port, 
      DATAPATH_I_ID_EX_RS1_NEXT_2_port, DATAPATH_I_ID_EX_RS1_NEXT_3_port, 
      DATAPATH_I_ID_EX_RS1_NEXT_4_port, DATAPATH_I_MEM_WB_RD_0_port, 
      DATAPATH_I_MEM_WB_RD_1_port, DATAPATH_I_MEM_WB_RD_2_port, 
      DATAPATH_I_MEM_WB_RD_3_port, DATAPATH_I_MEM_WB_RD_4_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_0_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_1_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_2_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_3_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_4_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_5_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_6_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_7_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_8_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_9_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_10_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_11_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_12_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_13_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_14_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_15_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_16_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_17_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_18_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_19_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_20_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_21_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_22_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_23_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_24_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_25_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_26_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_27_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_28_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_29_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_30_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_31_port, DATAPATH_I_MEM_WB_RF_WE, 
      DATAPATH_I_EX_MEM_RD_0_port, DATAPATH_I_EX_MEM_RD_1_port, 
      DATAPATH_I_EX_MEM_RD_2_port, DATAPATH_I_EX_MEM_RD_3_port, 
      DATAPATH_I_EX_MEM_RD_4_port, DATAPATH_I_ID_EX_RF_OUT2_0_port, 
      DATAPATH_I_ID_EX_RF_OUT2_1_port, DATAPATH_I_ID_EX_RF_OUT2_2_port, 
      DATAPATH_I_ID_EX_RF_OUT2_3_port, DATAPATH_I_ID_EX_RF_OUT2_4_port, 
      DATAPATH_I_ID_EX_RF_OUT2_5_port, DATAPATH_I_ID_EX_RF_OUT2_6_port, 
      DATAPATH_I_ID_EX_RF_OUT2_7_port, DATAPATH_I_ID_EX_RF_OUT2_8_port, 
      DATAPATH_I_ID_EX_RF_OUT2_9_port, DATAPATH_I_ID_EX_RF_OUT2_10_port, 
      DATAPATH_I_ID_EX_RF_OUT2_11_port, DATAPATH_I_ID_EX_RF_OUT2_12_port, 
      DATAPATH_I_ID_EX_RF_OUT2_13_port, DATAPATH_I_ID_EX_RF_OUT2_14_port, 
      DATAPATH_I_ID_EX_RF_OUT2_15_port, DATAPATH_I_ID_EX_RF_OUT2_16_port, 
      DATAPATH_I_ID_EX_RF_OUT2_17_port, DATAPATH_I_ID_EX_RF_OUT2_18_port, 
      DATAPATH_I_ID_EX_RF_OUT2_19_port, DATAPATH_I_ID_EX_RF_OUT2_20_port, 
      DATAPATH_I_ID_EX_RF_OUT2_21_port, DATAPATH_I_ID_EX_RF_OUT2_22_port, 
      DATAPATH_I_ID_EX_RF_OUT2_23_port, DATAPATH_I_ID_EX_RF_OUT2_24_port, 
      DATAPATH_I_ID_EX_RF_OUT2_25_port, DATAPATH_I_ID_EX_RF_OUT2_26_port, 
      DATAPATH_I_ID_EX_RF_OUT2_27_port, DATAPATH_I_ID_EX_RF_OUT2_28_port, 
      DATAPATH_I_ID_EX_RF_OUT2_29_port, DATAPATH_I_ID_EX_RF_OUT2_30_port, 
      DATAPATH_I_ID_EX_RF_OUT2_31_port, DATAPATH_I_ID_EX_RF_OUT1_0_port, 
      DATAPATH_I_ID_EX_RF_OUT1_1_port, DATAPATH_I_ID_EX_RF_OUT1_2_port, 
      DATAPATH_I_ID_EX_RF_OUT1_3_port, DATAPATH_I_ID_EX_RF_OUT1_4_port, 
      DATAPATH_I_ID_EX_RF_OUT1_5_port, DATAPATH_I_ID_EX_RF_OUT1_6_port, 
      DATAPATH_I_ID_EX_RF_OUT1_7_port, DATAPATH_I_ID_EX_RF_OUT1_8_port, 
      DATAPATH_I_ID_EX_RF_OUT1_9_port, DATAPATH_I_ID_EX_RF_OUT1_10_port, 
      DATAPATH_I_ID_EX_RF_OUT1_11_port, DATAPATH_I_ID_EX_RF_OUT1_12_port, 
      DATAPATH_I_ID_EX_RF_OUT1_13_port, DATAPATH_I_ID_EX_RF_OUT1_14_port, 
      DATAPATH_I_ID_EX_RF_OUT1_15_port, DATAPATH_I_ID_EX_RF_OUT1_16_port, 
      DATAPATH_I_ID_EX_RF_OUT1_17_port, DATAPATH_I_ID_EX_RF_OUT1_18_port, 
      DATAPATH_I_ID_EX_RF_OUT1_19_port, DATAPATH_I_ID_EX_RF_OUT1_20_port, 
      DATAPATH_I_ID_EX_RF_OUT1_21_port, DATAPATH_I_ID_EX_RF_OUT1_22_port, 
      DATAPATH_I_ID_EX_RF_OUT1_23_port, DATAPATH_I_ID_EX_RF_OUT1_24_port, 
      DATAPATH_I_ID_EX_RF_OUT1_25_port, DATAPATH_I_ID_EX_RF_OUT1_26_port, 
      DATAPATH_I_ID_EX_RF_OUT1_27_port, DATAPATH_I_ID_EX_RF_OUT1_28_port, 
      DATAPATH_I_ID_EX_RF_OUT1_29_port, DATAPATH_I_ID_EX_RF_OUT1_30_port, 
      DATAPATH_I_ID_EX_RF_OUT1_31_port, DATAPATH_I_ID_EX_RD_0_port, 
      DATAPATH_I_ID_EX_RD_1_port, DATAPATH_I_ID_EX_RD_2_port, 
      DATAPATH_I_ID_EX_RD_3_port, DATAPATH_I_ID_EX_RD_4_port, 
      DATAPATH_I_IF_ID_IR_11_port, DATAPATH_I_IF_ID_IR_12_port, 
      DATAPATH_I_IF_ID_IR_13_port, DATAPATH_I_IF_ID_IR_14_port, 
      DATAPATH_I_IF_ID_IR_15_port, DATAPATH_I_IF_ID_IR_16_port, 
      DATAPATH_I_IF_ID_IR_17_port, DATAPATH_I_IF_ID_IR_18_port, 
      DATAPATH_I_IF_ID_IR_19_port, DATAPATH_I_IF_ID_IR_20_port, 
      DATAPATH_I_IF_ID_IR_21_port, DATAPATH_I_IF_ID_IR_22_port, 
      DATAPATH_I_IF_ID_IR_23_port, DATAPATH_I_IF_ID_IR_24_port, 
      DATAPATH_I_IF_ID_IR_25_port, DATAPATH_I_IF_ID_IR_26_port, 
      DATAPATH_I_IF_ID_IR_27_port, DATAPATH_I_IF_ID_IR_28_port, 
      DATAPATH_I_IF_ID_IR_29_port, DATAPATH_I_IF_ID_IR_30_port, 
      DATAPATH_I_IF_ID_IR_31_port, DATAPATH_I_n29, DATAPATH_I_n28, 
      DATAPATH_I_n27, DATAPATH_I_n26, DATAPATH_I_n25, DATAPATH_I_n24, 
      DATAPATH_I_n23, DATAPATH_I_n22, DATAPATH_I_n21, DATAPATH_I_n20, 
      DATAPATH_I_n19, DATAPATH_I_n18, DATAPATH_I_n17, DATAPATH_I_n16, 
      DATAPATH_I_n15, DATAPATH_I_LATCH_LMD_LDI_0_N3, 
      DATAPATH_I_LATCH_LMD_LDI_1_N3, DATAPATH_I_LATCH_LMD_LDI_2_N3, 
      DATAPATH_I_LATCH_LMD_LDI_3_N3, DATAPATH_I_LATCH_LMD_LDI_4_N3, 
      DATAPATH_I_LATCH_LMD_LDI_5_N3, DATAPATH_I_LATCH_LMD_LDI_6_N3, 
      DATAPATH_I_LATCH_LMD_LDI_7_N3, DATAPATH_I_LATCH_LMD_LDI_8_N3, 
      DATAPATH_I_LATCH_LMD_LDI_9_N3, DATAPATH_I_LATCH_LMD_LDI_10_N3, 
      DATAPATH_I_LATCH_LMD_LDI_11_N3, DATAPATH_I_LATCH_LMD_LDI_12_N3, 
      DATAPATH_I_LATCH_LMD_LDI_13_N3, DATAPATH_I_LATCH_LMD_LDI_14_N3, 
      DATAPATH_I_LATCH_LMD_LDI_15_N3, DATAPATH_I_LATCH_LMD_LDI_16_N3, 
      DATAPATH_I_LATCH_LMD_LDI_17_N3, DATAPATH_I_LATCH_LMD_LDI_18_N3, 
      DATAPATH_I_LATCH_LMD_LDI_19_N3, DATAPATH_I_LATCH_LMD_LDI_20_N3, 
      DATAPATH_I_LATCH_LMD_LDI_21_N3, DATAPATH_I_LATCH_LMD_LDI_22_N3, 
      DATAPATH_I_LATCH_LMD_LDI_23_N3, DATAPATH_I_LATCH_LMD_LDI_24_N3, 
      DATAPATH_I_LATCH_LMD_LDI_25_N3, DATAPATH_I_LATCH_LMD_LDI_26_N3, 
      DATAPATH_I_LATCH_LMD_LDI_27_N3, DATAPATH_I_LATCH_LMD_LDI_28_N3, 
      DATAPATH_I_LATCH_LMD_LDI_29_N3, DATAPATH_I_LATCH_LMD_LDI_30_N3, 
      DATAPATH_I_LATCH_LMD_LDI_31_N3, DATAPATH_I_LATCH_ALUOUT_LDI_0_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_1_N3, DATAPATH_I_LATCH_ALUOUT_LDI_2_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_3_N3, DATAPATH_I_LATCH_ALUOUT_LDI_4_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_5_N3, DATAPATH_I_LATCH_ALUOUT_LDI_6_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_7_N3, DATAPATH_I_LATCH_ALUOUT_LDI_8_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_9_N3, DATAPATH_I_LATCH_ALUOUT_LDI_10_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_11_N3, DATAPATH_I_LATCH_ALUOUT_LDI_12_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_13_N3, DATAPATH_I_LATCH_ALUOUT_LDI_14_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_15_N3, DATAPATH_I_LATCH_ALUOUT_LDI_16_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_17_N3, DATAPATH_I_LATCH_ALUOUT_LDI_18_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_19_N3, DATAPATH_I_LATCH_ALUOUT_LDI_20_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_21_N3, DATAPATH_I_LATCH_ALUOUT_LDI_22_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_23_N3, DATAPATH_I_LATCH_ALUOUT_LDI_24_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_25_N3, DATAPATH_I_LATCH_ALUOUT_LDI_26_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_27_N3, DATAPATH_I_LATCH_ALUOUT_LDI_28_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_29_N3, DATAPATH_I_LATCH_ALUOUT_LDI_30_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_31_N3, DATAPATH_I_LATCH_RF2_LDI_0_N3, 
      DATAPATH_I_LATCH_RF2_LDI_1_N3, DATAPATH_I_LATCH_RF2_LDI_2_N3, 
      DATAPATH_I_LATCH_RF2_LDI_3_N3, DATAPATH_I_LATCH_RF2_LDI_4_N3, 
      DATAPATH_I_LATCH_RF2_LDI_5_N3, DATAPATH_I_LATCH_RF2_LDI_6_N3, 
      DATAPATH_I_LATCH_RF2_LDI_7_N3, DATAPATH_I_LATCH_RF2_LDI_8_N3, 
      DATAPATH_I_LATCH_RF2_LDI_9_N3, DATAPATH_I_LATCH_RF2_LDI_10_N3, 
      DATAPATH_I_LATCH_RF2_LDI_11_N3, DATAPATH_I_LATCH_RF2_LDI_12_N3, 
      DATAPATH_I_LATCH_RF2_LDI_13_N3, DATAPATH_I_LATCH_RF2_LDI_14_N3, 
      DATAPATH_I_LATCH_RF2_LDI_15_N3, DATAPATH_I_LATCH_RF2_LDI_16_N3, 
      DATAPATH_I_LATCH_RF2_LDI_17_N3, DATAPATH_I_LATCH_RF2_LDI_18_N3, 
      DATAPATH_I_LATCH_RF2_LDI_19_N3, DATAPATH_I_LATCH_RF2_LDI_20_N3, 
      DATAPATH_I_LATCH_RF2_LDI_21_N3, DATAPATH_I_LATCH_RF2_LDI_22_N3, 
      DATAPATH_I_LATCH_RF2_LDI_23_N3, DATAPATH_I_LATCH_RF2_LDI_24_N3, 
      DATAPATH_I_LATCH_RF2_LDI_25_N3, DATAPATH_I_LATCH_RF2_LDI_26_N3, 
      DATAPATH_I_LATCH_RF2_LDI_27_N3, DATAPATH_I_LATCH_RF2_LDI_28_N3, 
      DATAPATH_I_LATCH_RF2_LDI_29_N3, DATAPATH_I_LATCH_RF2_LDI_30_N3, 
      DATAPATH_I_LATCH_RF2_LDI_31_N3, DATAPATH_I_LATCH_RF1_LDI_0_N3, 
      DATAPATH_I_LATCH_RF1_LDI_1_N3, DATAPATH_I_LATCH_RF1_LDI_2_N3, 
      DATAPATH_I_LATCH_RF1_LDI_3_N3, DATAPATH_I_LATCH_RF1_LDI_4_N3, 
      DATAPATH_I_LATCH_RF1_LDI_5_N3, DATAPATH_I_LATCH_RF1_LDI_6_N3, 
      DATAPATH_I_LATCH_RF1_LDI_7_N3, DATAPATH_I_LATCH_RF1_LDI_8_N3, 
      DATAPATH_I_LATCH_RF1_LDI_9_N3, DATAPATH_I_LATCH_RF1_LDI_10_N3, 
      DATAPATH_I_LATCH_RF1_LDI_11_N3, DATAPATH_I_LATCH_RF1_LDI_12_N3, 
      DATAPATH_I_LATCH_RF1_LDI_13_N3, DATAPATH_I_LATCH_RF1_LDI_14_N3, 
      DATAPATH_I_LATCH_RF1_LDI_15_N3, DATAPATH_I_LATCH_RF1_LDI_16_N3, 
      DATAPATH_I_LATCH_RF1_LDI_17_N3, DATAPATH_I_LATCH_RF1_LDI_18_N3, 
      DATAPATH_I_LATCH_RF1_LDI_19_N3, DATAPATH_I_LATCH_RF1_LDI_20_N3, 
      DATAPATH_I_LATCH_RF1_LDI_21_N3, DATAPATH_I_LATCH_RF1_LDI_22_N3, 
      DATAPATH_I_LATCH_RF1_LDI_23_N3, DATAPATH_I_LATCH_RF1_LDI_24_N3, 
      DATAPATH_I_LATCH_RF1_LDI_25_N3, DATAPATH_I_LATCH_RF1_LDI_26_N3, 
      DATAPATH_I_LATCH_RF1_LDI_27_N3, DATAPATH_I_LATCH_RF1_LDI_28_N3, 
      DATAPATH_I_LATCH_RF1_LDI_29_N3, DATAPATH_I_LATCH_RF1_LDI_30_N3, 
      DATAPATH_I_LATCH_RF1_LDI_31_N3, DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_N3,
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_N3, n285, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, 
      n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, 
      n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
      n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, 
      n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, 
      n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, 
      n441, n442, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378 : std_logic;

begin
   
   IRAM_I : DLX_IRAM_RAM_DEPTH256_I_SIZE32 port map( RST => RST, ADDR(31) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(30) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(29) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(28) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(27) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(26) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(25) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(24) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(23) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(22) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(21) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(20) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(19) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(18) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(17) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(16) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(15) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(14) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(13) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(12) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(11) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(10) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(9) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(8) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(7) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(6) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(5) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(4) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(3) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(2) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(1) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(0) => 
                           DATAPATH_I_MEM_WB_RF_WE, DOUT(31) => IR_BUS_31_port,
                           DOUT(30) => IR_BUS_30_port, DOUT(29) => 
                           IR_BUS_29_port, DOUT(28) => IR_BUS_28_port, DOUT(27)
                           => IR_BUS_27_port, DOUT(26) => IR_BUS_26_port, 
                           DOUT(25) => IR_BUS_25_port, DOUT(24) => 
                           IR_BUS_24_port, DOUT(23) => IR_BUS_23_port, DOUT(22)
                           => IR_BUS_22_port, DOUT(21) => IR_BUS_21_port, 
                           DOUT(20) => IR_BUS_20_port, DOUT(19) => 
                           IR_BUS_19_port, DOUT(18) => IR_BUS_18_port, DOUT(17)
                           => IR_BUS_17_port, DOUT(16) => IR_BUS_16_port, 
                           DOUT(15) => IR_BUS_15_port, DOUT(14) => 
                           IR_BUS_14_port, DOUT(13) => IR_BUS_13_port, DOUT(12)
                           => IR_BUS_12_port, DOUT(11) => IR_BUS_11_port, 
                           DOUT(10) => IR_BUS_10_port, DOUT(9) => IR_BUS_9_port
                           , DOUT(8) => IR_BUS_8_port, DOUT(7) => IR_BUS_7_port
                           , DOUT(6) => IR_BUS_6_port, DOUT(5) => IR_BUS_5_port
                           , DOUT(4) => IR_BUS_4_port, DOUT(3) => IR_BUS_3_port
                           , DOUT(2) => IR_BUS_2_port, DOUT(1) => IR_BUS_1_port
                           , DOUT(0) => IR_BUS_0_port);
   DRAM_I : DLX_DRAM_N256_NW32 port map( CLK => CLK, RST => RST, RE => 
                           DATAPATH_I_MEM_WB_RF_WE, WE => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(31) => 
                           DATA_ADDR_31_port, ADDR(30) => DATA_ADDR_30_port, 
                           ADDR(29) => DATA_ADDR_29_port, ADDR(28) => 
                           DATA_ADDR_28_port, ADDR(27) => DATA_ADDR_27_port, 
                           ADDR(26) => DATA_ADDR_26_port, ADDR(25) => 
                           DATA_ADDR_25_port, ADDR(24) => DATA_ADDR_24_port, 
                           ADDR(23) => DATA_ADDR_23_port, ADDR(22) => 
                           DATA_ADDR_22_port, ADDR(21) => DATA_ADDR_21_port, 
                           ADDR(20) => DATA_ADDR_20_port, ADDR(19) => 
                           DATA_ADDR_19_port, ADDR(18) => DATA_ADDR_18_port, 
                           ADDR(17) => DATA_ADDR_17_port, ADDR(16) => 
                           DATA_ADDR_16_port, ADDR(15) => DATA_ADDR_15_port, 
                           ADDR(14) => DATA_ADDR_14_port, ADDR(13) => 
                           DATA_ADDR_13_port, ADDR(12) => DATA_ADDR_12_port, 
                           ADDR(11) => DATA_ADDR_11_port, ADDR(10) => 
                           DATA_ADDR_10_port, ADDR(9) => DATA_ADDR_9_port, 
                           ADDR(8) => DATA_ADDR_8_port, ADDR(7) => 
                           DATA_ADDR_7_port, ADDR(6) => DATA_ADDR_6_port, 
                           ADDR(5) => DATA_ADDR_5_port, ADDR(4) => 
                           DATA_ADDR_4_port, ADDR(3) => DATA_ADDR_3_port, 
                           ADDR(2) => DATA_ADDR_2_port, ADDR(1) => 
                           DATA_ADDR_1_port, ADDR(0) => DATA_ADDR_0_port, 
                           DIN(31) => DATA_IN_31_port, DIN(30) => 
                           DATA_IN_30_port, DIN(29) => DATA_IN_29_port, DIN(28)
                           => DATA_IN_28_port, DIN(27) => DATA_IN_27_port, 
                           DIN(26) => DATA_IN_26_port, DIN(25) => 
                           DATA_IN_25_port, DIN(24) => DATA_IN_24_port, DIN(23)
                           => DATA_IN_23_port, DIN(22) => DATA_IN_22_port, 
                           DIN(21) => DATA_IN_21_port, DIN(20) => 
                           DATA_IN_20_port, DIN(19) => DATA_IN_19_port, DIN(18)
                           => DATA_IN_18_port, DIN(17) => DATA_IN_17_port, 
                           DIN(16) => DATA_IN_16_port, DIN(15) => 
                           DATA_IN_15_port, DIN(14) => DATA_IN_14_port, DIN(13)
                           => DATA_IN_13_port, DIN(12) => DATA_IN_12_port, 
                           DIN(11) => DATA_IN_11_port, DIN(10) => 
                           DATA_IN_10_port, DIN(9) => DATA_IN_9_port, DIN(8) =>
                           DATA_IN_8_port, DIN(7) => DATA_IN_7_port, DIN(6) => 
                           DATA_IN_6_port, DIN(5) => DATA_IN_5_port, DIN(4) => 
                           DATA_IN_4_port, DIN(3) => DATA_IN_3_port, DIN(2) => 
                           DATA_IN_2_port, DIN(1) => DATA_IN_1_port, DIN(0) => 
                           DATA_IN_0_port, DOUT(31) => DATA_OUT_31_port, 
                           DOUT(30) => DATA_OUT_30_port, DOUT(29) => 
                           DATA_OUT_29_port, DOUT(28) => DATA_OUT_28_port, 
                           DOUT(27) => DATA_OUT_27_port, DOUT(26) => 
                           DATA_OUT_26_port, DOUT(25) => DATA_OUT_25_port, 
                           DOUT(24) => DATA_OUT_24_port, DOUT(23) => 
                           DATA_OUT_23_port, DOUT(22) => DATA_OUT_22_port, 
                           DOUT(21) => DATA_OUT_21_port, DOUT(20) => 
                           DATA_OUT_20_port, DOUT(19) => DATA_OUT_19_port, 
                           DOUT(18) => DATA_OUT_18_port, DOUT(17) => 
                           DATA_OUT_17_port, DOUT(16) => DATA_OUT_16_port, 
                           DOUT(15) => DATA_OUT_15_port, DOUT(14) => 
                           DATA_OUT_14_port, DOUT(13) => DATA_OUT_13_port, 
                           DOUT(12) => DATA_OUT_12_port, DOUT(11) => 
                           DATA_OUT_11_port, DOUT(10) => DATA_OUT_10_port, 
                           DOUT(9) => DATA_OUT_9_port, DOUT(8) => 
                           DATA_OUT_8_port, DOUT(7) => DATA_OUT_7_port, DOUT(6)
                           => DATA_OUT_6_port, DOUT(5) => DATA_OUT_5_port, 
                           DOUT(4) => DATA_OUT_4_port, DOUT(3) => 
                           DATA_OUT_3_port, DOUT(2) => DATA_OUT_2_port, DOUT(1)
                           => DATA_OUT_1_port, DOUT(0) => DATA_OUT_0_port);
   DATAPATH_I_ARITHMETIC_LOGIC_UNIT : ALU_N32_NB8 port map( OP1(31) => 
                           DATAPATH_I_ID_EX_RF_OUT1_31_port, OP1(30) => 
                           DATAPATH_I_ID_EX_RF_OUT1_30_port, OP1(29) => 
                           DATAPATH_I_ID_EX_RF_OUT1_29_port, OP1(28) => 
                           DATAPATH_I_ID_EX_RF_OUT1_28_port, OP1(27) => 
                           DATAPATH_I_ID_EX_RF_OUT1_27_port, OP1(26) => 
                           DATAPATH_I_ID_EX_RF_OUT1_26_port, OP1(25) => 
                           DATAPATH_I_ID_EX_RF_OUT1_25_port, OP1(24) => 
                           DATAPATH_I_ID_EX_RF_OUT1_24_port, OP1(23) => 
                           DATAPATH_I_ID_EX_RF_OUT1_23_port, OP1(22) => 
                           DATAPATH_I_ID_EX_RF_OUT1_22_port, OP1(21) => 
                           DATAPATH_I_ID_EX_RF_OUT1_21_port, OP1(20) => 
                           DATAPATH_I_ID_EX_RF_OUT1_20_port, OP1(19) => 
                           DATAPATH_I_ID_EX_RF_OUT1_19_port, OP1(18) => 
                           DATAPATH_I_ID_EX_RF_OUT1_18_port, OP1(17) => 
                           DATAPATH_I_ID_EX_RF_OUT1_17_port, OP1(16) => 
                           DATAPATH_I_ID_EX_RF_OUT1_16_port, OP1(15) => 
                           DATAPATH_I_ID_EX_RF_OUT1_15_port, OP1(14) => 
                           DATAPATH_I_ID_EX_RF_OUT1_14_port, OP1(13) => 
                           DATAPATH_I_ID_EX_RF_OUT1_13_port, OP1(12) => 
                           DATAPATH_I_ID_EX_RF_OUT1_12_port, OP1(11) => 
                           DATAPATH_I_ID_EX_RF_OUT1_11_port, OP1(10) => 
                           DATAPATH_I_ID_EX_RF_OUT1_10_port, OP1(9) => 
                           DATAPATH_I_ID_EX_RF_OUT1_9_port, OP1(8) => 
                           DATAPATH_I_ID_EX_RF_OUT1_8_port, OP1(7) => 
                           DATAPATH_I_ID_EX_RF_OUT1_7_port, OP1(6) => 
                           DATAPATH_I_ID_EX_RF_OUT1_6_port, OP1(5) => 
                           DATAPATH_I_ID_EX_RF_OUT1_5_port, OP1(4) => 
                           DATAPATH_I_ID_EX_RF_OUT1_4_port, OP1(3) => 
                           DATAPATH_I_ID_EX_RF_OUT1_3_port, OP1(2) => 
                           DATAPATH_I_ID_EX_RF_OUT1_2_port, OP1(1) => 
                           DATAPATH_I_ID_EX_RF_OUT1_1_port, OP1(0) => 
                           DATAPATH_I_ID_EX_RF_OUT1_0_port, OP2(31) => 
                           DATAPATH_I_ID_EX_RF_OUT2_31_port, OP2(30) => 
                           DATAPATH_I_ID_EX_RF_OUT2_30_port, OP2(29) => 
                           DATAPATH_I_ID_EX_RF_OUT2_29_port, OP2(28) => 
                           DATAPATH_I_ID_EX_RF_OUT2_28_port, OP2(27) => 
                           DATAPATH_I_ID_EX_RF_OUT2_27_port, OP2(26) => 
                           DATAPATH_I_ID_EX_RF_OUT2_26_port, OP2(25) => 
                           DATAPATH_I_ID_EX_RF_OUT2_25_port, OP2(24) => 
                           DATAPATH_I_ID_EX_RF_OUT2_24_port, OP2(23) => 
                           DATAPATH_I_ID_EX_RF_OUT2_23_port, OP2(22) => 
                           DATAPATH_I_ID_EX_RF_OUT2_22_port, OP2(21) => 
                           DATAPATH_I_ID_EX_RF_OUT2_21_port, OP2(20) => 
                           DATAPATH_I_ID_EX_RF_OUT2_20_port, OP2(19) => 
                           DATAPATH_I_ID_EX_RF_OUT2_19_port, OP2(18) => 
                           DATAPATH_I_ID_EX_RF_OUT2_18_port, OP2(17) => 
                           DATAPATH_I_ID_EX_RF_OUT2_17_port, OP2(16) => 
                           DATAPATH_I_ID_EX_RF_OUT2_16_port, OP2(15) => 
                           DATAPATH_I_ID_EX_RF_OUT2_15_port, OP2(14) => 
                           DATAPATH_I_ID_EX_RF_OUT2_14_port, OP2(13) => 
                           DATAPATH_I_ID_EX_RF_OUT2_13_port, OP2(12) => 
                           DATAPATH_I_ID_EX_RF_OUT2_12_port, OP2(11) => 
                           DATAPATH_I_ID_EX_RF_OUT2_11_port, OP2(10) => 
                           DATAPATH_I_ID_EX_RF_OUT2_10_port, OP2(9) => 
                           DATAPATH_I_ID_EX_RF_OUT2_9_port, OP2(8) => 
                           DATAPATH_I_ID_EX_RF_OUT2_8_port, OP2(7) => 
                           DATAPATH_I_ID_EX_RF_OUT2_7_port, OP2(6) => 
                           DATAPATH_I_ID_EX_RF_OUT2_6_port, OP2(5) => 
                           DATAPATH_I_ID_EX_RF_OUT2_5_port, OP2(4) => 
                           DATAPATH_I_ID_EX_RF_OUT2_4_port, OP2(3) => 
                           DATAPATH_I_ID_EX_RF_OUT2_3_port, OP2(2) => 
                           DATAPATH_I_ID_EX_RF_OUT2_2_port, OP2(1) => 
                           DATAPATH_I_ID_EX_RF_OUT2_1_port, OP2(0) => 
                           DATAPATH_I_ID_EX_RF_OUT2_0_port, OPC(0) => 
                           ALU_OPCODE_i_0_port, OPC(1) => ALU_OPCODE_i_1_port, 
                           OPC(2) => ALU_OPCODE_i_2_port, OPC(3) => 
                           ALU_OPCODE_i_3_port, OPC(4) => ALU_OPCODE_i_4_port, 
                           OPC(5) => ALU_OPCODE_i_5_port, OPC(6) => 
                           ALU_OPCODE_i_6_port, Y(31) => 
                           DATAPATH_I_ALU_OUTPUT_31_port, Y(30) => 
                           DATAPATH_I_ALU_OUTPUT_30_port, Y(29) => 
                           DATAPATH_I_ALU_OUTPUT_29_port, Y(28) => 
                           DATAPATH_I_ALU_OUTPUT_28_port, Y(27) => 
                           DATAPATH_I_ALU_OUTPUT_27_port, Y(26) => 
                           DATAPATH_I_ALU_OUTPUT_26_port, Y(25) => 
                           DATAPATH_I_ALU_OUTPUT_25_port, Y(24) => 
                           DATAPATH_I_ALU_OUTPUT_24_port, Y(23) => 
                           DATAPATH_I_ALU_OUTPUT_23_port, Y(22) => 
                           DATAPATH_I_ALU_OUTPUT_22_port, Y(21) => 
                           DATAPATH_I_ALU_OUTPUT_21_port, Y(20) => 
                           DATAPATH_I_ALU_OUTPUT_20_port, Y(19) => 
                           DATAPATH_I_ALU_OUTPUT_19_port, Y(18) => 
                           DATAPATH_I_ALU_OUTPUT_18_port, Y(17) => 
                           DATAPATH_I_ALU_OUTPUT_17_port, Y(16) => 
                           DATAPATH_I_ALU_OUTPUT_16_port, Y(15) => 
                           DATAPATH_I_ALU_OUTPUT_15_port, Y(14) => 
                           DATAPATH_I_ALU_OUTPUT_14_port, Y(13) => 
                           DATAPATH_I_ALU_OUTPUT_13_port, Y(12) => 
                           DATAPATH_I_ALU_OUTPUT_12_port, Y(11) => 
                           DATAPATH_I_ALU_OUTPUT_11_port, Y(10) => 
                           DATAPATH_I_ALU_OUTPUT_10_port, Y(9) => 
                           DATAPATH_I_ALU_OUTPUT_9_port, Y(8) => 
                           DATAPATH_I_ALU_OUTPUT_8_port, Y(7) => 
                           DATAPATH_I_ALU_OUTPUT_7_port, Y(6) => 
                           DATAPATH_I_ALU_OUTPUT_6_port, Y(5) => 
                           DATAPATH_I_ALU_OUTPUT_5_port, Y(4) => 
                           DATAPATH_I_ALU_OUTPUT_4_port, Y(3) => 
                           DATAPATH_I_ALU_OUTPUT_3_port, Y(2) => 
                           DATAPATH_I_ALU_OUTPUT_2_port, Y(1) => 
                           DATAPATH_I_ALU_OUTPUT_1_port, Y(0) => 
                           DATAPATH_I_ALU_OUTPUT_0_port, Z => n_1171);
   DATAPATH_I_REGISTER_FILE : RF_N32_NA5 port map( RST => RST, EN => n285, 
                           EN_RD1 => n285, EN_RD2 => n285, EN_WR => 
                           DATAPATH_I_MEM_WB_RF_WE, ADD_RD1(4) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_4_port, ADD_RD1(3) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_3_port, ADD_RD1(2) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_2_port, ADD_RD1(1) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_1_port, ADD_RD1(0) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_0_port, ADD_RD2(4) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_4_port, ADD_RD2(3) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_3_port, ADD_RD2(2) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_2_port, ADD_RD2(1) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_1_port, ADD_RD2(0) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_0_port, ADD_WR(4) => 
                           DATAPATH_I_MEM_WB_RD_4_port, ADD_WR(3) => 
                           DATAPATH_I_MEM_WB_RD_3_port, ADD_WR(2) => 
                           DATAPATH_I_MEM_WB_RD_2_port, ADD_WR(1) => 
                           DATAPATH_I_MEM_WB_RD_1_port, ADD_WR(0) => 
                           DATAPATH_I_MEM_WB_RD_0_port, DATAIN(31) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_31_port, DATAIN(30) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_30_port, DATAIN(29) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_29_port, DATAIN(28) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_28_port, DATAIN(27) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_27_port, DATAIN(26) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_26_port, DATAIN(25) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_25_port, DATAIN(24) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_24_port, DATAIN(23) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_23_port, DATAIN(22) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_22_port, DATAIN(21) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_21_port, DATAIN(20) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_20_port, DATAIN(19) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_19_port, DATAIN(18) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_18_port, DATAIN(17) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_17_port, DATAIN(16) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_16_port, DATAIN(15) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_15_port, DATAIN(14) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_14_port, DATAIN(13) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_13_port, DATAIN(12) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_12_port, DATAIN(11) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_11_port, DATAIN(10) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_10_port, DATAIN(9) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_9_port, DATAIN(8) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_8_port, DATAIN(7) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_7_port, DATAIN(6) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_6_port, DATAIN(5) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_5_port, DATAIN(4) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_4_port, DATAIN(3) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_3_port, DATAIN(2) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_2_port, DATAIN(1) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_1_port, DATAIN(0) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_0_port, OUT1(31) => 
                           DATAPATH_I_RF_OUT1_31_port, OUT1(30) => 
                           DATAPATH_I_RF_OUT1_30_port, OUT1(29) => 
                           DATAPATH_I_RF_OUT1_29_port, OUT1(28) => 
                           DATAPATH_I_RF_OUT1_28_port, OUT1(27) => 
                           DATAPATH_I_RF_OUT1_27_port, OUT1(26) => 
                           DATAPATH_I_RF_OUT1_26_port, OUT1(25) => 
                           DATAPATH_I_RF_OUT1_25_port, OUT1(24) => 
                           DATAPATH_I_RF_OUT1_24_port, OUT1(23) => 
                           DATAPATH_I_RF_OUT1_23_port, OUT1(22) => 
                           DATAPATH_I_RF_OUT1_22_port, OUT1(21) => 
                           DATAPATH_I_RF_OUT1_21_port, OUT1(20) => 
                           DATAPATH_I_RF_OUT1_20_port, OUT1(19) => 
                           DATAPATH_I_RF_OUT1_19_port, OUT1(18) => 
                           DATAPATH_I_RF_OUT1_18_port, OUT1(17) => 
                           DATAPATH_I_RF_OUT1_17_port, OUT1(16) => 
                           DATAPATH_I_RF_OUT1_16_port, OUT1(15) => 
                           DATAPATH_I_RF_OUT1_15_port, OUT1(14) => 
                           DATAPATH_I_RF_OUT1_14_port, OUT1(13) => 
                           DATAPATH_I_RF_OUT1_13_port, OUT1(12) => 
                           DATAPATH_I_RF_OUT1_12_port, OUT1(11) => 
                           DATAPATH_I_RF_OUT1_11_port, OUT1(10) => 
                           DATAPATH_I_RF_OUT1_10_port, OUT1(9) => 
                           DATAPATH_I_RF_OUT1_9_port, OUT1(8) => 
                           DATAPATH_I_RF_OUT1_8_port, OUT1(7) => 
                           DATAPATH_I_RF_OUT1_7_port, OUT1(6) => 
                           DATAPATH_I_RF_OUT1_6_port, OUT1(5) => 
                           DATAPATH_I_RF_OUT1_5_port, OUT1(4) => 
                           DATAPATH_I_RF_OUT1_4_port, OUT1(3) => 
                           DATAPATH_I_RF_OUT1_3_port, OUT1(2) => 
                           DATAPATH_I_RF_OUT1_2_port, OUT1(1) => 
                           DATAPATH_I_RF_OUT1_1_port, OUT1(0) => 
                           DATAPATH_I_RF_OUT1_0_port, OUT2(31) => 
                           DATAPATH_I_RF_OUT2_31_port, OUT2(30) => 
                           DATAPATH_I_RF_OUT2_30_port, OUT2(29) => 
                           DATAPATH_I_RF_OUT2_29_port, OUT2(28) => 
                           DATAPATH_I_RF_OUT2_28_port, OUT2(27) => 
                           DATAPATH_I_RF_OUT2_27_port, OUT2(26) => 
                           DATAPATH_I_RF_OUT2_26_port, OUT2(25) => 
                           DATAPATH_I_RF_OUT2_25_port, OUT2(24) => 
                           DATAPATH_I_RF_OUT2_24_port, OUT2(23) => 
                           DATAPATH_I_RF_OUT2_23_port, OUT2(22) => 
                           DATAPATH_I_RF_OUT2_22_port, OUT2(21) => 
                           DATAPATH_I_RF_OUT2_21_port, OUT2(20) => 
                           DATAPATH_I_RF_OUT2_20_port, OUT2(19) => 
                           DATAPATH_I_RF_OUT2_19_port, OUT2(18) => 
                           DATAPATH_I_RF_OUT2_18_port, OUT2(17) => 
                           DATAPATH_I_RF_OUT2_17_port, OUT2(16) => 
                           DATAPATH_I_RF_OUT2_16_port, OUT2(15) => 
                           DATAPATH_I_RF_OUT2_15_port, OUT2(14) => 
                           DATAPATH_I_RF_OUT2_14_port, OUT2(13) => 
                           DATAPATH_I_RF_OUT2_13_port, OUT2(12) => 
                           DATAPATH_I_RF_OUT2_12_port, OUT2(11) => 
                           DATAPATH_I_RF_OUT2_11_port, OUT2(10) => 
                           DATAPATH_I_RF_OUT2_10_port, OUT2(9) => 
                           DATAPATH_I_RF_OUT2_9_port, OUT2(8) => 
                           DATAPATH_I_RF_OUT2_8_port, OUT2(7) => 
                           DATAPATH_I_RF_OUT2_7_port, OUT2(6) => 
                           DATAPATH_I_RF_OUT2_6_port, OUT2(5) => 
                           DATAPATH_I_RF_OUT2_5_port, OUT2(4) => 
                           DATAPATH_I_RF_OUT2_4_port, OUT2(3) => 
                           DATAPATH_I_RF_OUT2_3_port, OUT2(2) => 
                           DATAPATH_I_RF_OUT2_2_port, OUT2(1) => 
                           DATAPATH_I_RF_OUT2_1_port, OUT2(0) => 
                           DATAPATH_I_RF_OUT2_0_port);
   DATAPATH_I_IF_ID_IR_reg_11_inst : DFF_X1 port map( D => DATAPATH_I_N45, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_11_port, QN => 
                           n_1172);
   DATAPATH_I_IF_ID_IR_reg_12_inst : DFF_X1 port map( D => DATAPATH_I_N46, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_12_port, QN => 
                           n_1173);
   DATAPATH_I_IF_ID_IR_reg_13_inst : DFF_X1 port map( D => DATAPATH_I_N47, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_13_port, QN => 
                           n_1174);
   DATAPATH_I_IF_ID_IR_reg_14_inst : DFF_X1 port map( D => DATAPATH_I_N48, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_14_port, QN => 
                           n_1175);
   DATAPATH_I_IF_ID_IR_reg_15_inst : DFF_X1 port map( D => DATAPATH_I_N49, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_15_port, QN => 
                           n_1176);
   DATAPATH_I_IF_ID_IR_reg_16_inst : DFF_X1 port map( D => DATAPATH_I_N50, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_16_port, QN => 
                           n_1177);
   DATAPATH_I_IF_ID_IR_reg_17_inst : DFF_X1 port map( D => DATAPATH_I_N51, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_17_port, QN => 
                           n_1178);
   DATAPATH_I_IF_ID_IR_reg_18_inst : DFF_X1 port map( D => DATAPATH_I_N52, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_18_port, QN => 
                           n_1179);
   DATAPATH_I_IF_ID_IR_reg_19_inst : DFF_X1 port map( D => DATAPATH_I_N53, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_19_port, QN => 
                           n_1180);
   DATAPATH_I_IF_ID_IR_reg_20_inst : DFF_X1 port map( D => DATAPATH_I_N54, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_20_port, QN => 
                           n_1181);
   DATAPATH_I_IF_ID_IR_reg_21_inst : DFF_X1 port map( D => DATAPATH_I_N55, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_21_port, QN => 
                           n_1182);
   DATAPATH_I_IF_ID_IR_reg_22_inst : DFF_X1 port map( D => DATAPATH_I_N56, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_22_port, QN => 
                           n_1183);
   DATAPATH_I_IF_ID_IR_reg_23_inst : DFF_X1 port map( D => DATAPATH_I_N57, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_23_port, QN => 
                           n_1184);
   DATAPATH_I_IF_ID_IR_reg_24_inst : DFF_X1 port map( D => DATAPATH_I_N58, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_24_port, QN => 
                           n_1185);
   DATAPATH_I_IF_ID_IR_reg_25_inst : DFF_X1 port map( D => DATAPATH_I_N59, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_25_port, QN => 
                           n_1186);
   DATAPATH_I_IF_ID_IR_reg_26_inst : DFF_X1 port map( D => DATAPATH_I_N60, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_26_port, QN => n440
                           );
   DATAPATH_I_IF_ID_IR_reg_27_inst : DFF_X1 port map( D => DATAPATH_I_N61, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_27_port, QN => n441
                           );
   DATAPATH_I_IF_ID_IR_reg_28_inst : DFF_X1 port map( D => DATAPATH_I_N62, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_28_port, QN => 
                           n_1187);
   DATAPATH_I_IF_ID_IR_reg_29_inst : DFF_X1 port map( D => DATAPATH_I_N63, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_29_port, QN => 
                           n_1188);
   DATAPATH_I_IF_ID_IR_reg_30_inst : DFF_X1 port map( D => DATAPATH_I_N64, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_30_port, QN => n442
                           );
   DATAPATH_I_IF_ID_IR_reg_31_inst : DFF_X1 port map( D => DATAPATH_I_N65, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_31_port, QN => 
                           n_1189);
   DATAPATH_I_EX_MEM_RD_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N308, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_0_port, QN => 
                           n_1190);
   DATAPATH_I_MEM_WB_RD_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N410, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_0_port, QN => 
                           n_1191);
   DATAPATH_I_EX_MEM_RD_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N309, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_1_port, QN => 
                           n_1192);
   DATAPATH_I_MEM_WB_RD_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N411, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_1_port, QN => 
                           n_1193);
   DATAPATH_I_EX_MEM_RD_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N310, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_2_port, QN => 
                           n_1194);
   DATAPATH_I_MEM_WB_RD_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N412, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_2_port, QN => 
                           n_1195);
   DATAPATH_I_ID_EX_RD_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N112, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_3_port, QN => 
                           n_1196);
   DATAPATH_I_EX_MEM_RD_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N311, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_3_port, QN => 
                           n_1197);
   DATAPATH_I_MEM_WB_RD_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N413, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_3_port, QN => 
                           n_1198);
   DATAPATH_I_ID_EX_RD_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N113, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_4_port, QN => 
                           n_1199);
   DATAPATH_I_EX_MEM_RD_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N312, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_4_port, QN => 
                           n_1200);
   DATAPATH_I_MEM_WB_RD_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N414, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_4_port, QN => 
                           n_1201);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_0_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N275, CK => CLK, Q => DATA_ADDR_0_port, 
                           QN => n_1202);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_1_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N276, CK => CLK, Q => DATA_ADDR_1_port, 
                           QN => n_1203);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_2_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N277, CK => CLK, Q => DATA_ADDR_2_port, 
                           QN => n_1204);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_3_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N278, CK => CLK, Q => DATA_ADDR_3_port, 
                           QN => n_1205);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_4_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N279, CK => CLK, Q => DATA_ADDR_4_port, 
                           QN => n_1206);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_5_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N280, CK => CLK, Q => DATA_ADDR_5_port, 
                           QN => n_1207);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_6_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N281, CK => CLK, Q => DATA_ADDR_6_port, 
                           QN => n_1208);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_7_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N282, CK => CLK, Q => DATA_ADDR_7_port, 
                           QN => n_1209);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_8_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N283, CK => CLK, Q => DATA_ADDR_8_port, 
                           QN => n_1210);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_9_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N284, CK => CLK, Q => DATA_ADDR_9_port, 
                           QN => n_1211);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_10_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N285, CK => CLK, Q => DATA_ADDR_10_port, 
                           QN => n_1212);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_11_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N286, CK => CLK, Q => DATA_ADDR_11_port, 
                           QN => n_1213);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_12_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N287, CK => CLK, Q => DATA_ADDR_12_port, 
                           QN => n_1214);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_13_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N288, CK => CLK, Q => DATA_ADDR_13_port, 
                           QN => n_1215);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_14_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N289, CK => CLK, Q => DATA_ADDR_14_port, 
                           QN => n_1216);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_15_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N290, CK => CLK, Q => DATA_ADDR_15_port, 
                           QN => n_1217);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_16_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N291, CK => CLK, Q => DATA_ADDR_16_port, 
                           QN => n_1218);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_17_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N292, CK => CLK, Q => DATA_ADDR_17_port, 
                           QN => n_1219);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_18_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N293, CK => CLK, Q => DATA_ADDR_18_port, 
                           QN => n_1220);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_19_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N294, CK => CLK, Q => DATA_ADDR_19_port, 
                           QN => n_1221);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_20_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N295, CK => CLK, Q => DATA_ADDR_20_port, 
                           QN => n_1222);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_21_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N296, CK => CLK, Q => DATA_ADDR_21_port, 
                           QN => n_1223);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_22_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N297, CK => CLK, Q => DATA_ADDR_22_port, 
                           QN => n_1224);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_23_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N298, CK => CLK, Q => DATA_ADDR_23_port, 
                           QN => n_1225);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_24_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N299, CK => CLK, Q => DATA_ADDR_24_port, 
                           QN => n_1226);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_25_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N300, CK => CLK, Q => DATA_ADDR_25_port, 
                           QN => n_1227);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_26_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N301, CK => CLK, Q => DATA_ADDR_26_port, 
                           QN => n_1228);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_27_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N302, CK => CLK, Q => DATA_ADDR_27_port, 
                           QN => n_1229);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_28_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N303, CK => CLK, Q => DATA_ADDR_28_port, 
                           QN => n_1230);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_29_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N304, CK => CLK, Q => DATA_ADDR_29_port, 
                           QN => n_1231);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_30_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N305, CK => CLK, Q => DATA_ADDR_30_port, 
                           QN => n_1232);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_31_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N306, CK => CLK, Q => DATA_ADDR_31_port, 
                           QN => n_1233);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_0_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N378, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_0_port, QN => n_1234);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_1_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N379, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_1_port, QN => n_1235);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_2_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N380, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_2_port, QN => n_1236);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_3_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N381, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_3_port, QN => n_1237);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_4_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N382, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_4_port, QN => n_1238);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_5_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N383, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_5_port, QN => n_1239);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_6_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N384, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_6_port, QN => n_1240);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_7_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N385, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_7_port, QN => n_1241);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_8_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N386, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_8_port, QN => n_1242);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_9_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N387, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_9_port, QN => n_1243);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_10_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N388, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_10_port, QN => n_1244)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_11_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N389, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_11_port, QN => n_1245)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_12_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N390, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_12_port, QN => n_1246)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_13_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N391, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_13_port, QN => n_1247)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_14_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N392, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_14_port, QN => n_1248)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_15_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N393, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_15_port, QN => n_1249)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_16_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N394, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_16_port, QN => n_1250)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_17_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N395, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_17_port, QN => n_1251)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_18_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N396, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_18_port, QN => n_1252)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_19_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N397, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_19_port, QN => n_1253)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_20_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N398, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_20_port, QN => n_1254)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_21_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N399, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_21_port, QN => n_1255)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_22_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N400, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_22_port, QN => n_1256)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_23_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N401, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_23_port, QN => n_1257)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_24_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N402, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_24_port, QN => n_1258)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_25_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N403, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_25_port, QN => n_1259)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_26_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N404, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_26_port, QN => n_1260)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_27_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N405, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_27_port, QN => n_1261)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_28_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N406, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_28_port, QN => n_1262)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_29_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N407, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_29_port, QN => n_1263)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_30_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N408, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_30_port, QN => n_1264)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_31_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N409, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_31_port, QN => n_1265)
                           ;
   DATAPATH_I_ID_EX_RF_OUT2_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N146,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_0_port, QN 
                           => n_1266);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N243
                           , CK => CLK, Q => DATA_IN_0_port, QN => n_1267);
   DATAPATH_I_ID_EX_RF_OUT2_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N147,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_1_port, QN 
                           => n_1268);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N244
                           , CK => CLK, Q => DATA_IN_1_port, QN => n_1269);
   DATAPATH_I_ID_EX_RF_OUT2_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N148,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_2_port, QN 
                           => n_1270);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N245
                           , CK => CLK, Q => DATA_IN_2_port, QN => n_1271);
   DATAPATH_I_ID_EX_RF_OUT2_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N149,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_3_port, QN 
                           => n_1272);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N246
                           , CK => CLK, Q => DATA_IN_3_port, QN => n_1273);
   DATAPATH_I_ID_EX_RF_OUT2_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N150,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_4_port, QN 
                           => n_1274);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N247
                           , CK => CLK, Q => DATA_IN_4_port, QN => n_1275);
   DATAPATH_I_ID_EX_RF_OUT2_reg_5_inst : DFF_X1 port map( D => DATAPATH_I_N151,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_5_port, QN 
                           => n_1276);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_5_inst : DFF_X1 port map( D => DATAPATH_I_N248
                           , CK => CLK, Q => DATA_IN_5_port, QN => n_1277);
   DATAPATH_I_ID_EX_RF_OUT2_reg_6_inst : DFF_X1 port map( D => DATAPATH_I_N152,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_6_port, QN 
                           => n_1278);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_6_inst : DFF_X1 port map( D => DATAPATH_I_N249
                           , CK => CLK, Q => DATA_IN_6_port, QN => n_1279);
   DATAPATH_I_ID_EX_RF_OUT2_reg_7_inst : DFF_X1 port map( D => DATAPATH_I_N153,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_7_port, QN 
                           => n_1280);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_7_inst : DFF_X1 port map( D => DATAPATH_I_N250
                           , CK => CLK, Q => DATA_IN_7_port, QN => n_1281);
   DATAPATH_I_ID_EX_RF_OUT2_reg_8_inst : DFF_X1 port map( D => DATAPATH_I_N154,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_8_port, QN 
                           => n_1282);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_8_inst : DFF_X1 port map( D => DATAPATH_I_N251
                           , CK => CLK, Q => DATA_IN_8_port, QN => n_1283);
   DATAPATH_I_ID_EX_RF_OUT2_reg_9_inst : DFF_X1 port map( D => DATAPATH_I_N155,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_9_port, QN 
                           => n_1284);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_9_inst : DFF_X1 port map( D => DATAPATH_I_N252
                           , CK => CLK, Q => DATA_IN_9_port, QN => n_1285);
   DATAPATH_I_ID_EX_RF_OUT2_reg_10_inst : DFF_X1 port map( D => DATAPATH_I_N156
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_10_port, 
                           QN => n_1286);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_10_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N253, CK => CLK, Q => DATA_IN_10_port, QN
                           => n_1287);
   DATAPATH_I_ID_EX_RF_OUT2_reg_11_inst : DFF_X1 port map( D => DATAPATH_I_N157
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_11_port, 
                           QN => n_1288);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_11_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N254, CK => CLK, Q => DATA_IN_11_port, QN
                           => n_1289);
   DATAPATH_I_ID_EX_RF_OUT2_reg_12_inst : DFF_X1 port map( D => DATAPATH_I_N158
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_12_port, 
                           QN => n_1290);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_12_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N255, CK => CLK, Q => DATA_IN_12_port, QN
                           => n_1291);
   DATAPATH_I_ID_EX_RF_OUT2_reg_13_inst : DFF_X1 port map( D => DATAPATH_I_N159
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_13_port, 
                           QN => n_1292);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_13_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N256, CK => CLK, Q => DATA_IN_13_port, QN
                           => n_1293);
   DATAPATH_I_ID_EX_RF_OUT2_reg_14_inst : DFF_X1 port map( D => DATAPATH_I_N160
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_14_port, 
                           QN => n_1294);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_14_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N257, CK => CLK, Q => DATA_IN_14_port, QN
                           => n_1295);
   DATAPATH_I_ID_EX_RF_OUT2_reg_15_inst : DFF_X1 port map( D => DATAPATH_I_N161
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_15_port, 
                           QN => n_1296);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_15_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N258, CK => CLK, Q => DATA_IN_15_port, QN
                           => n_1297);
   DATAPATH_I_ID_EX_RF_OUT2_reg_16_inst : DFF_X1 port map( D => DATAPATH_I_N162
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_16_port, 
                           QN => n_1298);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_16_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N259, CK => CLK, Q => DATA_IN_16_port, QN
                           => n_1299);
   DATAPATH_I_ID_EX_RF_OUT2_reg_17_inst : DFF_X1 port map( D => DATAPATH_I_N163
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_17_port, 
                           QN => n_1300);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_17_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N260, CK => CLK, Q => DATA_IN_17_port, QN
                           => n_1301);
   DATAPATH_I_ID_EX_RF_OUT2_reg_18_inst : DFF_X1 port map( D => DATAPATH_I_N164
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_18_port, 
                           QN => n_1302);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_18_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N261, CK => CLK, Q => DATA_IN_18_port, QN
                           => n_1303);
   DATAPATH_I_ID_EX_RF_OUT2_reg_19_inst : DFF_X1 port map( D => DATAPATH_I_N165
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_19_port, 
                           QN => n_1304);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_19_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N262, CK => CLK, Q => DATA_IN_19_port, QN
                           => n_1305);
   DATAPATH_I_ID_EX_RF_OUT2_reg_20_inst : DFF_X1 port map( D => DATAPATH_I_N166
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_20_port, 
                           QN => n_1306);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_20_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N263, CK => CLK, Q => DATA_IN_20_port, QN
                           => n_1307);
   DATAPATH_I_ID_EX_RF_OUT2_reg_21_inst : DFF_X1 port map( D => DATAPATH_I_N167
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_21_port, 
                           QN => n_1308);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_21_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N264, CK => CLK, Q => DATA_IN_21_port, QN
                           => n_1309);
   DATAPATH_I_ID_EX_RF_OUT2_reg_22_inst : DFF_X1 port map( D => DATAPATH_I_N168
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_22_port, 
                           QN => n_1310);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_22_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N265, CK => CLK, Q => DATA_IN_22_port, QN
                           => n_1311);
   DATAPATH_I_ID_EX_RF_OUT2_reg_23_inst : DFF_X1 port map( D => DATAPATH_I_N169
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_23_port, 
                           QN => n_1312);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_23_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N266, CK => CLK, Q => DATA_IN_23_port, QN
                           => n_1313);
   DATAPATH_I_ID_EX_RF_OUT2_reg_24_inst : DFF_X1 port map( D => DATAPATH_I_N170
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_24_port, 
                           QN => n_1314);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_24_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N267, CK => CLK, Q => DATA_IN_24_port, QN
                           => n_1315);
   DATAPATH_I_ID_EX_RF_OUT2_reg_25_inst : DFF_X1 port map( D => DATAPATH_I_N171
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_25_port, 
                           QN => n_1316);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_25_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N268, CK => CLK, Q => DATA_IN_25_port, QN
                           => n_1317);
   DATAPATH_I_ID_EX_RF_OUT2_reg_26_inst : DFF_X1 port map( D => DATAPATH_I_N172
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_26_port, 
                           QN => n_1318);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_26_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N269, CK => CLK, Q => DATA_IN_26_port, QN
                           => n_1319);
   DATAPATH_I_ID_EX_RF_OUT2_reg_27_inst : DFF_X1 port map( D => DATAPATH_I_N173
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_27_port, 
                           QN => n_1320);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_27_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N270, CK => CLK, Q => DATA_IN_27_port, QN
                           => n_1321);
   DATAPATH_I_ID_EX_RF_OUT2_reg_28_inst : DFF_X1 port map( D => DATAPATH_I_N174
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_28_port, 
                           QN => n_1322);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_28_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N271, CK => CLK, Q => DATA_IN_28_port, QN
                           => n_1323);
   DATAPATH_I_ID_EX_RF_OUT2_reg_29_inst : DFF_X1 port map( D => DATAPATH_I_N175
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_29_port, 
                           QN => n_1324);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_29_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N272, CK => CLK, Q => DATA_IN_29_port, QN
                           => n_1325);
   DATAPATH_I_ID_EX_RF_OUT2_reg_30_inst : DFF_X1 port map( D => DATAPATH_I_N176
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_30_port, 
                           QN => n_1326);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_30_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N273, CK => CLK, Q => DATA_IN_30_port, QN
                           => n_1327);
   DATAPATH_I_ID_EX_RF_OUT2_reg_31_inst : DFF_X1 port map( D => DATAPATH_I_N177
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_31_port, 
                           QN => n_1328);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_31_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N274, CK => CLK, Q => DATA_IN_31_port, QN
                           => n_1329);
   DATAPATH_I_ID_EX_RF_OUT1_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N114,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_0_port, QN 
                           => n_1330);
   DATAPATH_I_ID_EX_RF_OUT1_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N115,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_1_port, QN 
                           => n_1331);
   DATAPATH_I_ID_EX_RF_OUT1_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N116,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_2_port, QN 
                           => n_1332);
   DATAPATH_I_ID_EX_RF_OUT1_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N117,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_3_port, QN 
                           => n_1333);
   DATAPATH_I_ID_EX_RF_OUT1_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N118,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_4_port, QN 
                           => n_1334);
   DATAPATH_I_ID_EX_RF_OUT1_reg_5_inst : DFF_X1 port map( D => DATAPATH_I_N119,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_5_port, QN 
                           => n_1335);
   DATAPATH_I_ID_EX_RF_OUT1_reg_6_inst : DFF_X1 port map( D => DATAPATH_I_N120,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_6_port, QN 
                           => n_1336);
   DATAPATH_I_ID_EX_RF_OUT1_reg_7_inst : DFF_X1 port map( D => DATAPATH_I_N121,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_7_port, QN 
                           => n_1337);
   DATAPATH_I_ID_EX_RF_OUT1_reg_8_inst : DFF_X1 port map( D => DATAPATH_I_N122,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_8_port, QN 
                           => n_1338);
   DATAPATH_I_ID_EX_RF_OUT1_reg_9_inst : DFF_X1 port map( D => DATAPATH_I_N123,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_9_port, QN 
                           => n_1339);
   DATAPATH_I_ID_EX_RF_OUT1_reg_10_inst : DFF_X1 port map( D => DATAPATH_I_N124
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_10_port, 
                           QN => n_1340);
   DATAPATH_I_ID_EX_RF_OUT1_reg_11_inst : DFF_X1 port map( D => DATAPATH_I_N125
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_11_port, 
                           QN => n_1341);
   DATAPATH_I_ID_EX_RF_OUT1_reg_12_inst : DFF_X1 port map( D => DATAPATH_I_N126
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_12_port, 
                           QN => n_1342);
   DATAPATH_I_ID_EX_RF_OUT1_reg_13_inst : DFF_X1 port map( D => DATAPATH_I_N127
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_13_port, 
                           QN => n_1343);
   DATAPATH_I_ID_EX_RF_OUT1_reg_14_inst : DFF_X1 port map( D => DATAPATH_I_N128
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_14_port, 
                           QN => n_1344);
   DATAPATH_I_ID_EX_RF_OUT1_reg_15_inst : DFF_X1 port map( D => DATAPATH_I_N129
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_15_port, 
                           QN => n_1345);
   DATAPATH_I_ID_EX_RF_OUT1_reg_16_inst : DFF_X1 port map( D => DATAPATH_I_N130
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_16_port, 
                           QN => n_1346);
   DATAPATH_I_ID_EX_RF_OUT1_reg_17_inst : DFF_X1 port map( D => DATAPATH_I_N131
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_17_port, 
                           QN => n_1347);
   DATAPATH_I_ID_EX_RF_OUT1_reg_18_inst : DFF_X1 port map( D => DATAPATH_I_N132
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_18_port, 
                           QN => n_1348);
   DATAPATH_I_ID_EX_RF_OUT1_reg_19_inst : DFF_X1 port map( D => DATAPATH_I_N133
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_19_port, 
                           QN => n_1349);
   DATAPATH_I_ID_EX_RF_OUT1_reg_20_inst : DFF_X1 port map( D => DATAPATH_I_N134
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_20_port, 
                           QN => n_1350);
   DATAPATH_I_ID_EX_RF_OUT1_reg_21_inst : DFF_X1 port map( D => DATAPATH_I_N135
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_21_port, 
                           QN => n_1351);
   DATAPATH_I_ID_EX_RF_OUT1_reg_22_inst : DFF_X1 port map( D => DATAPATH_I_N136
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_22_port, 
                           QN => n_1352);
   DATAPATH_I_ID_EX_RF_OUT1_reg_23_inst : DFF_X1 port map( D => DATAPATH_I_N137
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_23_port, 
                           QN => n_1353);
   DATAPATH_I_ID_EX_RF_OUT1_reg_24_inst : DFF_X1 port map( D => DATAPATH_I_N138
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_24_port, 
                           QN => n_1354);
   DATAPATH_I_ID_EX_RF_OUT1_reg_25_inst : DFF_X1 port map( D => DATAPATH_I_N139
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_25_port, 
                           QN => n_1355);
   DATAPATH_I_ID_EX_RF_OUT1_reg_26_inst : DFF_X1 port map( D => DATAPATH_I_N140
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_26_port, 
                           QN => n_1356);
   DATAPATH_I_ID_EX_RF_OUT1_reg_27_inst : DFF_X1 port map( D => DATAPATH_I_N141
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_27_port, 
                           QN => n_1357);
   DATAPATH_I_ID_EX_RF_OUT1_reg_28_inst : DFF_X1 port map( D => DATAPATH_I_N142
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_28_port, 
                           QN => n_1358);
   DATAPATH_I_ID_EX_RF_OUT1_reg_29_inst : DFF_X1 port map( D => DATAPATH_I_N143
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_29_port, 
                           QN => n_1359);
   DATAPATH_I_ID_EX_RF_OUT1_reg_30_inst : DFF_X1 port map( D => DATAPATH_I_N144
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_30_port, 
                           QN => n_1360);
   DATAPATH_I_ID_EX_RF_OUT1_reg_31_inst : DFF_X1 port map( D => DATAPATH_I_N145
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_31_port, 
                           QN => n_1361);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_N3, GN => RST,
                           Q => IR_0_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_N3, GN => RST,
                           Q => IR_1_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_N3, GN => RST,
                           Q => IR_2_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_N3, GN => RST,
                           Q => IR_3_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_N3, GN => RST,
                           Q => IR_4_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_N3, GN => RST,
                           Q => IR_5_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_N3, GN => RST,
                           Q => IR_6_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_N3, GN => RST,
                           Q => IR_7_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_N3, GN => RST,
                           Q => IR_8_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_N3, GN => RST,
                           Q => IR_9_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_N3, GN => RST
                           , Q => IR_10_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_N3, GN => RST
                           , Q => DATAPATH_I_n29);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_N3, GN => RST
                           , Q => DATAPATH_I_n28);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_N3, GN => RST
                           , Q => DATAPATH_I_n27);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_N3, GN => RST
                           , Q => DATAPATH_I_n26);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_N3, GN => RST
                           , Q => DATAPATH_I_n25);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_N3, GN => RST
                           , Q => DATAPATH_I_n24);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_N3, GN => RST
                           , Q => DATAPATH_I_n23);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_N3, GN => RST
                           , Q => DATAPATH_I_n22);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_N3, GN => RST
                           , Q => DATAPATH_I_n21);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_N3, GN => RST
                           , Q => DATAPATH_I_n20);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_N3, GN => RST
                           , Q => DATAPATH_I_n19);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_N3, GN => RST
                           , Q => DATAPATH_I_n18);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_N3, GN => RST
                           , Q => DATAPATH_I_n17);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_N3, GN => RST
                           , Q => DATAPATH_I_n16);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_N3, GN => RST
                           , Q => DATAPATH_I_n15);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_N3, GN => RST
                           , Q => IR_26_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_N3, GN => RST
                           , Q => IR_27_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_N3, GN => RST
                           , Q => IR_28_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_N3, GN => RST
                           , Q => IR_29_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_N3, GN => RST
                           , Q => IR_30_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_N3, GN => RST
                           , Q => IR_31_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_0_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_0_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_1_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_1_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_2_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_2_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_3_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_3_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_4_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_4_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_5_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_5_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_6_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_6_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_7_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_7_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_8_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_8_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_9_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_9_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_10_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_10_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_11_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_11_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_12_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_12_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_13_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_13_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_14_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_14_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_15_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_15_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_16_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_16_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_17_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_17_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_18_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_18_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_19_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_19_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_20_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_20_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_21_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_21_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_22_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_22_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_23_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_23_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_24_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_24_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_25_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_25_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_26_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_26_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_27_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_27_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_28_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_28_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_29_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_29_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_30_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_30_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_31_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_31_port);
   DATAPATH_I_LATCH_LMD_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_0_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_0_port);
   DATAPATH_I_LATCH_LMD_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_1_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_1_port);
   DATAPATH_I_LATCH_LMD_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_2_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_2_port);
   DATAPATH_I_LATCH_LMD_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_3_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_3_port);
   DATAPATH_I_LATCH_LMD_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_4_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_4_port);
   DATAPATH_I_LATCH_LMD_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_5_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_5_port);
   DATAPATH_I_LATCH_LMD_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_6_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_6_port);
   DATAPATH_I_LATCH_LMD_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_7_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_7_port);
   DATAPATH_I_LATCH_LMD_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_8_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_8_port);
   DATAPATH_I_LATCH_LMD_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_9_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_9_port);
   DATAPATH_I_LATCH_LMD_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_10_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_10_port);
   DATAPATH_I_LATCH_LMD_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_11_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_11_port);
   DATAPATH_I_LATCH_LMD_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_12_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_12_port);
   DATAPATH_I_LATCH_LMD_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_13_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_13_port);
   DATAPATH_I_LATCH_LMD_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_14_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_14_port);
   DATAPATH_I_LATCH_LMD_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_15_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_15_port);
   DATAPATH_I_LATCH_LMD_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_16_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_16_port);
   DATAPATH_I_LATCH_LMD_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_17_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_17_port);
   DATAPATH_I_LATCH_LMD_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_18_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_18_port);
   DATAPATH_I_LATCH_LMD_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_19_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_19_port);
   DATAPATH_I_LATCH_LMD_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_20_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_20_port);
   DATAPATH_I_LATCH_LMD_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_21_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_21_port);
   DATAPATH_I_LATCH_LMD_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_22_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_22_port);
   DATAPATH_I_LATCH_LMD_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_23_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_23_port);
   DATAPATH_I_LATCH_LMD_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_24_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_24_port);
   DATAPATH_I_LATCH_LMD_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_25_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_25_port);
   DATAPATH_I_LATCH_LMD_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_26_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_26_port);
   DATAPATH_I_LATCH_LMD_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_27_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_27_port);
   DATAPATH_I_LATCH_LMD_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_28_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_28_port);
   DATAPATH_I_LATCH_LMD_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_29_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_29_port);
   DATAPATH_I_LATCH_LMD_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_30_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_30_port);
   DATAPATH_I_LATCH_LMD_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_31_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_31_port);
   DATAPATH_I_LATCH_RF2_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_0_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_0_port);
   DATAPATH_I_LATCH_RF2_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_1_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_1_port);
   DATAPATH_I_LATCH_RF2_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_2_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_2_port);
   DATAPATH_I_LATCH_RF2_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_3_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_3_port);
   DATAPATH_I_LATCH_RF2_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_4_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_4_port);
   DATAPATH_I_LATCH_RF2_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_5_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_5_port);
   DATAPATH_I_LATCH_RF2_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_6_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_6_port);
   DATAPATH_I_LATCH_RF2_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_7_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_7_port);
   DATAPATH_I_LATCH_RF2_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_8_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_8_port);
   DATAPATH_I_LATCH_RF2_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_9_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_9_port);
   DATAPATH_I_LATCH_RF2_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_10_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_10_port);
   DATAPATH_I_LATCH_RF2_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_11_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_11_port);
   DATAPATH_I_LATCH_RF2_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_12_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_12_port);
   DATAPATH_I_LATCH_RF2_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_13_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_13_port);
   DATAPATH_I_LATCH_RF2_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_14_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_14_port);
   DATAPATH_I_LATCH_RF2_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_15_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_15_port);
   DATAPATH_I_LATCH_RF2_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_16_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_16_port);
   DATAPATH_I_LATCH_RF2_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_17_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_17_port);
   DATAPATH_I_LATCH_RF2_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_18_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_18_port);
   DATAPATH_I_LATCH_RF2_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_19_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_19_port);
   DATAPATH_I_LATCH_RF2_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_20_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_20_port);
   DATAPATH_I_LATCH_RF2_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_21_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_21_port);
   DATAPATH_I_LATCH_RF2_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_22_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_22_port);
   DATAPATH_I_LATCH_RF2_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_23_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_23_port);
   DATAPATH_I_LATCH_RF2_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_24_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_24_port);
   DATAPATH_I_LATCH_RF2_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_25_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_25_port);
   DATAPATH_I_LATCH_RF2_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_26_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_26_port);
   DATAPATH_I_LATCH_RF2_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_27_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_27_port);
   DATAPATH_I_LATCH_RF2_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_28_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_28_port);
   DATAPATH_I_LATCH_RF2_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_29_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_29_port);
   DATAPATH_I_LATCH_RF2_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_30_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_30_port);
   DATAPATH_I_LATCH_RF2_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_31_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_31_port);
   DATAPATH_I_LATCH_RF1_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_0_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_0_port);
   DATAPATH_I_LATCH_RF1_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_1_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_1_port);
   DATAPATH_I_LATCH_RF1_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_2_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_2_port);
   DATAPATH_I_LATCH_RF1_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_3_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_3_port);
   DATAPATH_I_LATCH_RF1_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_4_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_4_port);
   DATAPATH_I_LATCH_RF1_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_5_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_5_port);
   DATAPATH_I_LATCH_RF1_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_6_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_6_port);
   DATAPATH_I_LATCH_RF1_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_7_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_7_port);
   DATAPATH_I_LATCH_RF1_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_8_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_8_port);
   DATAPATH_I_LATCH_RF1_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_9_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_9_port);
   DATAPATH_I_LATCH_RF1_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_10_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_10_port);
   DATAPATH_I_LATCH_RF1_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_11_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_11_port);
   DATAPATH_I_LATCH_RF1_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_12_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_12_port);
   DATAPATH_I_LATCH_RF1_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_13_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_13_port);
   DATAPATH_I_LATCH_RF1_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_14_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_14_port);
   DATAPATH_I_LATCH_RF1_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_15_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_15_port);
   DATAPATH_I_LATCH_RF1_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_16_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_16_port);
   DATAPATH_I_LATCH_RF1_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_17_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_17_port);
   DATAPATH_I_LATCH_RF1_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_18_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_18_port);
   DATAPATH_I_LATCH_RF1_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_19_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_19_port);
   DATAPATH_I_LATCH_RF1_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_20_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_20_port);
   DATAPATH_I_LATCH_RF1_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_21_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_21_port);
   DATAPATH_I_LATCH_RF1_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_22_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_22_port);
   DATAPATH_I_LATCH_RF1_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_23_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_23_port);
   DATAPATH_I_LATCH_RF1_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_24_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_24_port);
   DATAPATH_I_LATCH_RF1_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_25_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_25_port);
   DATAPATH_I_LATCH_RF1_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_26_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_26_port);
   DATAPATH_I_LATCH_RF1_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_27_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_27_port);
   DATAPATH_I_LATCH_RF1_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_28_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_28_port);
   DATAPATH_I_LATCH_RF1_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_29_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_29_port);
   DATAPATH_I_LATCH_RF1_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_30_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_30_port);
   DATAPATH_I_LATCH_RF1_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_31_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_31_port);
   CU_I_aluOpcode2_reg_0_inst : DFFR_X1 port map( D => CU_I_aluOpcode1_0_port, 
                           CK => CLK, RN => RST, Q => CU_I_aluOpcode2_0_port, 
                           QN => n_1362);
   CU_I_aluOpcode3_reg_0_inst : DFFR_X1 port map( D => CU_I_aluOpcode2_0_port, 
                           CK => CLK, RN => RST, Q => ALU_OPCODE_i_6_port, QN 
                           => n_1363);
   CU_I_aluOpcode2_reg_3_inst : DFFR_X1 port map( D => CU_I_aluOpcode1_3_port, 
                           CK => CLK, RN => RST, Q => CU_I_aluOpcode2_3_port, 
                           QN => n_1364);
   CU_I_aluOpcode3_reg_3_inst : DFFR_X1 port map( D => CU_I_aluOpcode2_3_port, 
                           CK => CLK, RN => RST, Q => ALU_OPCODE_i_3_port, QN 
                           => n_1365);
   CU_I_aluOpcode2_reg_4_inst : DFFR_X1 port map( D => CU_I_aluOpcode1_4_port, 
                           CK => CLK, RN => RST, Q => CU_I_aluOpcode2_4_port, 
                           QN => n_1366);
   CU_I_aluOpcode3_reg_4_inst : DFFR_X1 port map( D => CU_I_aluOpcode2_4_port, 
                           CK => CLK, RN => RST, Q => ALU_OPCODE_i_2_port, QN 
                           => n_1367);
   CU_I_aluOpcode2_reg_2_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_2_port, 
                           CK => CLK, SN => RST, Q => CU_I_aluOpcode2_2_port, 
                           QN => n_1368);
   CU_I_aluOpcode3_reg_2_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_2_port, 
                           CK => CLK, SN => RST, Q => ALU_OPCODE_i_4_port, QN 
                           => n_1369);
   CU_I_aluOpcode2_reg_1_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_1_port, 
                           CK => CLK, SN => RST, Q => CU_I_aluOpcode2_1_port, 
                           QN => n_1370);
   CU_I_aluOpcode3_reg_1_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_1_port, 
                           CK => CLK, SN => RST, Q => ALU_OPCODE_i_5_port, QN 
                           => n_1371);
   CU_I_aluOpcode2_reg_5_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_5_port, 
                           CK => CLK, SN => RST, Q => CU_I_aluOpcode2_5_port, 
                           QN => n_1372);
   CU_I_aluOpcode3_reg_5_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_5_port, 
                           CK => CLK, SN => RST, Q => ALU_OPCODE_i_1_port, QN 
                           => n_1373);
   CU_I_aluOpcode2_reg_6_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_6_port, 
                           CK => CLK, SN => RST, Q => CU_I_aluOpcode2_6_port, 
                           QN => n_1374);
   CU_I_aluOpcode3_reg_6_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_6_port, 
                           CK => CLK, SN => RST, Q => ALU_OPCODE_i_0_port, QN 
                           => n_1375);
   DATAPATH_I_ID_EX_RD_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N111, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_2_port, QN => 
                           n_1376);
   DATAPATH_I_ID_EX_RD_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N109, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_0_port, QN => 
                           n_1377);
   DATAPATH_I_ID_EX_RD_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N110, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_1_port, QN => 
                           n_1378);
   U751 : INV_X1 port map( A => RST, ZN => n317);
   U752 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_0_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_N3);
   U753 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_1_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_N3);
   U754 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_2_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_N3);
   U755 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_3_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_N3);
   U756 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_4_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_N3);
   U757 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_5_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_N3);
   U758 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_6_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_N3);
   U759 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_7_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_N3);
   U760 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_8_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_N3);
   U761 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_9_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_N3);
   U762 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_10_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_N3);
   U763 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_11_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_N3);
   U764 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_12_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_N3);
   U765 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_13_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_N3);
   U766 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_14_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_N3);
   U767 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_15_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_N3);
   U768 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_16_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_N3);
   U769 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_17_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_N3);
   U770 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_18_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_N3);
   U771 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_19_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_N3);
   U772 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_20_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_N3);
   U773 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_21_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_N3);
   U774 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_22_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_N3);
   U775 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_23_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_N3);
   U776 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_24_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_N3);
   U777 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_25_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_N3);
   U778 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_26_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_N3);
   U779 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_27_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_N3);
   U780 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_28_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_N3);
   U781 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_29_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_N3);
   U782 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_30_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_N3);
   U783 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_31_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_N3);
   U784 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_0_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_0_N3);
   U785 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_1_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_1_N3);
   U786 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_2_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_2_N3);
   U787 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_3_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_3_N3);
   U788 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_4_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_4_N3);
   U789 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_5_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_5_N3);
   U790 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_6_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_6_N3);
   U791 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_7_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_7_N3);
   U792 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_8_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_8_N3);
   U793 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_9_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_9_N3);
   U794 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_10_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_10_N3);
   U795 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_11_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_11_N3);
   U796 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_12_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_12_N3);
   U797 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_13_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_13_N3);
   U798 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_14_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_14_N3);
   U799 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_15_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_15_N3);
   U800 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_16_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_16_N3);
   U801 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_17_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_17_N3);
   U802 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_18_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_18_N3);
   U803 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_19_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_19_N3);
   U804 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_20_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_20_N3);
   U805 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_21_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_21_N3);
   U806 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_22_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_22_N3);
   U807 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_23_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_23_N3);
   U808 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_24_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_24_N3);
   U809 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_25_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_25_N3);
   U810 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_26_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_26_N3);
   U811 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_27_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_27_N3);
   U812 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_28_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_28_N3);
   U813 : INV_X1 port map( A => IR_28_port, ZN => n407);
   U814 : NOR2_X1 port map( A1 => n317, A2 => n407, ZN => DATAPATH_I_N62);
   U815 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_29_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_29_N3);
   U816 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_30_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_30_N3);
   U817 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_31_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_31_N3);
   U818 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_0_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_0_N3);
   U819 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_1_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_1_N3);
   U820 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_2_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_2_N3);
   U821 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_3_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_3_N3);
   U822 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_4_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_4_N3);
   U823 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_5_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_5_N3);
   U824 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_6_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_6_N3);
   U825 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_7_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_7_N3);
   U826 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_8_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_8_N3);
   U827 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_9_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_9_N3);
   U828 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_10_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_10_N3);
   U829 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_11_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_11_N3);
   U830 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_12_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_12_N3);
   U831 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_13_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_13_N3);
   U832 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_15_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_15_N3);
   U833 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_16_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_16_N3);
   U834 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_17_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_17_N3);
   U835 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_18_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_18_N3);
   U836 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_19_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_19_N3);
   U837 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_20_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_20_N3);
   U838 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_21_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_21_N3);
   U839 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_22_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_22_N3);
   U840 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_23_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_23_N3);
   U841 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_24_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_24_N3);
   U842 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_25_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_25_N3);
   U843 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_26_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_26_N3);
   U844 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_27_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_27_N3);
   U845 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_28_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_28_N3);
   U846 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_29_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_29_N3);
   U847 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_30_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_30_N3);
   U848 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_31_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_31_N3);
   U849 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_0_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_0_N3);
   U850 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_1_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_1_N3);
   U851 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_2_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_2_N3);
   U852 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_3_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_3_N3);
   U853 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_4_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_4_N3);
   U854 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_5_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_5_N3);
   U855 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_6_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_6_N3);
   U856 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_7_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_7_N3);
   U857 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_8_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_8_N3);
   U858 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_9_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_9_N3);
   U859 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_10_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_10_N3);
   U860 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_11_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_11_N3);
   U861 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_12_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_12_N3);
   U862 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_13_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_13_N3);
   U863 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_14_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_14_N3);
   U864 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_15_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_15_N3);
   U865 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_16_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_16_N3);
   U866 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_17_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_17_N3);
   U867 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_18_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_18_N3);
   U868 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_19_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_19_N3);
   U869 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_20_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_20_N3);
   U870 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_21_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_21_N3);
   U871 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_22_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_22_N3);
   U872 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_23_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_23_N3);
   U873 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_24_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_24_N3);
   U874 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_25_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_25_N3);
   U875 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_26_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_26_N3);
   U876 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_27_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_27_N3);
   U877 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_28_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_28_N3);
   U878 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_29_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_29_N3);
   U879 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_30_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_30_N3);
   U880 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_14_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_14_N3);
   U881 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_31_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_31_N3);
   U882 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_0_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_0_N3);
   U883 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_1_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_1_N3);
   U884 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_2_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_2_N3);
   U885 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_3_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_3_N3);
   U886 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_4_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_4_N3);
   U887 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_5_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_5_N3);
   U888 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_6_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_6_N3);
   U889 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_7_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_7_N3);
   U890 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_8_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_8_N3);
   U891 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_9_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_9_N3);
   U892 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_10_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_10_N3);
   U893 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_11_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_11_N3);
   U894 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_12_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_12_N3);
   U895 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_13_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_13_N3);
   U896 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_14_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_14_N3);
   U897 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_15_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_15_N3);
   U898 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_16_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_16_N3);
   U899 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_17_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_17_N3);
   U900 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_18_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_18_N3);
   U901 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_30_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_30_N3);
   U902 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_19_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_19_N3);
   U903 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_23_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_23_N3);
   U904 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_20_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_20_N3);
   U905 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_27_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_27_N3);
   U906 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_21_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_21_N3);
   U907 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_24_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_24_N3);
   U908 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_22_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_22_N3);
   U909 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_28_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_28_N3);
   U910 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_29_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_29_N3);
   U911 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_25_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_25_N3);
   U912 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_26_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_26_N3);
   U913 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_31_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_31_N3);
   U914 : NOR4_X1 port map( A1 => DATAPATH_I_IF_ID_IR_28_port, A2 => 
                           DATAPATH_I_IF_ID_IR_29_port, A3 => 
                           DATAPATH_I_IF_ID_IR_31_port, A4 => n441, ZN => n347)
                           ;
   U915 : NAND2_X1 port map( A1 => n347, A2 => n442, ZN => n318);
   U916 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_25_port, A2 => n318, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_4_port);
   U917 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_23_port, A2 => n318, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_2_port);
   U918 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_22_port, A2 => n318, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_1_port);
   U919 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_21_port, A2 => n318, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_0_port);
   U920 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_0_port, ZN => 
                           DATAPATH_I_N308);
   U921 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_3_port, ZN => 
                           DATAPATH_I_N311);
   U922 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_2_port, ZN =>
                           DATAPATH_I_N412);
   U923 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_4_port, ZN =>
                           DATAPATH_I_N414);
   U924 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_3_port, ZN =>
                           DATAPATH_I_N413);
   U925 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_1_port, ZN =>
                           DATAPATH_I_N411);
   U926 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_0_port, ZN =>
                           DATAPATH_I_N410);
   U927 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_1_port, ZN => 
                           DATAPATH_I_N309);
   U928 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_2_port, ZN => 
                           DATAPATH_I_N310);
   U929 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_4_port, ZN => 
                           DATAPATH_I_N312);
   U930 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_12_port, ZN => 
                           DATAPATH_I_N126);
   U931 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_9_port, ZN => 
                           DATAPATH_I_N123);
   U932 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_11_port, ZN => 
                           DATAPATH_I_N125);
   U933 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_14_port, ZN => 
                           DATAPATH_I_N128);
   U934 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_18_port, ZN => 
                           DATAPATH_I_N132);
   U935 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_10_port, ZN => 
                           DATAPATH_I_N124);
   U936 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_17_port, ZN => 
                           DATAPATH_I_N131);
   U937 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_3_port, ZN => 
                           DATAPATH_I_N117);
   U938 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_4_port, ZN => 
                           DATAPATH_I_N118);
   U939 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_13_port, ZN => 
                           DATAPATH_I_N127);
   U940 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_2_port, ZN => 
                           DATAPATH_I_N116);
   U941 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_5_port, ZN => 
                           DATAPATH_I_N119);
   U942 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_20_port, ZN => 
                           DATAPATH_I_N134);
   U943 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_1_port, ZN => 
                           DATAPATH_I_N115);
   U944 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_7_port, ZN => 
                           DATAPATH_I_N121);
   U945 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_0_port, ZN => 
                           DATAPATH_I_N114);
   U946 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_21_port, ZN => 
                           DATAPATH_I_N135);
   U947 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_6_port, ZN => 
                           DATAPATH_I_N120);
   U948 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_31_port, ZN => 
                           DATAPATH_I_N177);
   U949 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_15_port, ZN => 
                           DATAPATH_I_N129);
   U950 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_22_port, ZN => 
                           DATAPATH_I_N136);
   U951 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_30_port, ZN => 
                           DATAPATH_I_N176);
   U952 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_8_port, ZN => 
                           DATAPATH_I_N122);
   U953 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_29_port, ZN => 
                           DATAPATH_I_N175);
   U954 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_23_port, ZN => 
                           DATAPATH_I_N137);
   U955 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_16_port, ZN => 
                           DATAPATH_I_N130);
   U956 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_28_port, ZN => 
                           DATAPATH_I_N174);
   U957 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_19_port, ZN => 
                           DATAPATH_I_N133);
   U958 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_24_port, ZN => 
                           DATAPATH_I_N138);
   U959 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_27_port, ZN => 
                           DATAPATH_I_N173);
   U960 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_25_port, ZN => 
                           DATAPATH_I_N139);
   U961 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_26_port, ZN => 
                           DATAPATH_I_N140);
   U962 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_27_port, ZN => 
                           DATAPATH_I_N141);
   U963 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_28_port, ZN => 
                           DATAPATH_I_N142);
   U964 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_29_port, ZN => 
                           DATAPATH_I_N143);
   U965 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_30_port, ZN => 
                           DATAPATH_I_N144);
   U966 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_31_port, ZN => 
                           DATAPATH_I_N145);
   U967 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n28, ZN => 
                           DATAPATH_I_N46);
   U968 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n27, ZN => 
                           DATAPATH_I_N47);
   U969 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n26, ZN => 
                           DATAPATH_I_N48);
   U970 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n25, ZN => 
                           DATAPATH_I_N49);
   U971 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n24, ZN => 
                           DATAPATH_I_N50);
   U972 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n23, ZN => 
                           DATAPATH_I_N51);
   U973 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n22, ZN => 
                           DATAPATH_I_N52);
   U974 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n21, ZN => 
                           DATAPATH_I_N53);
   U975 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n20, ZN => 
                           DATAPATH_I_N54);
   U976 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n19, ZN => 
                           DATAPATH_I_N55);
   U977 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n18, ZN => 
                           DATAPATH_I_N56);
   U978 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n17, ZN => 
                           DATAPATH_I_N57);
   U979 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n16, ZN => 
                           DATAPATH_I_N58);
   U980 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n15, ZN => 
                           DATAPATH_I_N59);
   U981 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_0_port, ZN => 
                           DATAPATH_I_N275);
   U982 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_1_port, ZN => 
                           DATAPATH_I_N276);
   U983 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_2_port, ZN => 
                           DATAPATH_I_N277);
   U984 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_3_port, ZN => 
                           DATAPATH_I_N278);
   U985 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_4_port, ZN => 
                           DATAPATH_I_N279);
   U986 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_5_port, ZN => 
                           DATAPATH_I_N280);
   U987 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_6_port, ZN => 
                           DATAPATH_I_N281);
   U988 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_7_port, ZN => 
                           DATAPATH_I_N282);
   U989 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_8_port, ZN => 
                           DATAPATH_I_N283);
   U990 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_9_port, ZN => 
                           DATAPATH_I_N284);
   U991 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_10_port, ZN => 
                           DATAPATH_I_N285);
   U992 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_11_port, ZN => 
                           DATAPATH_I_N286);
   U993 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_12_port, ZN => 
                           DATAPATH_I_N287);
   U994 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_13_port, ZN => 
                           DATAPATH_I_N288);
   U995 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_14_port, ZN => 
                           DATAPATH_I_N289);
   U996 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_15_port, ZN => 
                           DATAPATH_I_N290);
   U997 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_16_port, ZN => 
                           DATAPATH_I_N291);
   U998 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_17_port, ZN => 
                           DATAPATH_I_N292);
   U999 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_18_port, ZN => 
                           DATAPATH_I_N293);
   U1000 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_19_port, ZN => 
                           DATAPATH_I_N294);
   U1001 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_20_port, ZN => 
                           DATAPATH_I_N295);
   U1002 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_21_port, ZN => 
                           DATAPATH_I_N296);
   U1003 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_22_port, ZN => 
                           DATAPATH_I_N297);
   U1004 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_23_port, ZN => 
                           DATAPATH_I_N298);
   U1005 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_24_port, ZN => 
                           DATAPATH_I_N299);
   U1006 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_25_port, ZN => 
                           DATAPATH_I_N300);
   U1007 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_26_port, ZN => 
                           DATAPATH_I_N301);
   U1008 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_27_port, ZN => 
                           DATAPATH_I_N302);
   U1009 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_28_port, ZN => 
                           DATAPATH_I_N303);
   U1010 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_29_port, ZN => 
                           DATAPATH_I_N304);
   U1011 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_30_port, ZN => 
                           DATAPATH_I_N305);
   U1012 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_31_port, ZN => 
                           DATAPATH_I_N306);
   U1013 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_0_port, ZN => 
                           DATAPATH_I_N378);
   U1014 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_1_port, ZN => 
                           DATAPATH_I_N379);
   U1015 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_2_port, ZN => 
                           DATAPATH_I_N380);
   U1016 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n29, ZN => 
                           DATAPATH_I_N45);
   U1017 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_3_port, ZN => 
                           DATAPATH_I_N381);
   U1018 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_4_port, ZN => 
                           DATAPATH_I_N382);
   U1019 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_5_port, ZN => 
                           DATAPATH_I_N383);
   U1020 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_6_port, ZN => 
                           DATAPATH_I_N384);
   U1021 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_7_port, ZN => 
                           DATAPATH_I_N385);
   U1022 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_9_port, ZN => 
                           DATAPATH_I_N387);
   U1023 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_10_port, ZN => 
                           DATAPATH_I_N388);
   U1024 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_11_port, ZN => 
                           DATAPATH_I_N389);
   U1025 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_12_port, ZN => 
                           DATAPATH_I_N390);
   U1026 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_13_port, ZN => 
                           DATAPATH_I_N391);
   U1027 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_14_port, ZN => 
                           DATAPATH_I_N392);
   U1028 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_15_port, ZN => 
                           DATAPATH_I_N393);
   U1029 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_16_port, ZN => 
                           DATAPATH_I_N394);
   U1030 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_17_port, ZN => 
                           DATAPATH_I_N395);
   U1031 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_18_port, ZN => 
                           DATAPATH_I_N396);
   U1032 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_19_port, ZN => 
                           DATAPATH_I_N397);
   U1033 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_20_port, ZN => 
                           DATAPATH_I_N398);
   U1034 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_21_port, ZN => 
                           DATAPATH_I_N399);
   U1035 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_22_port, ZN => 
                           DATAPATH_I_N400);
   U1036 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_23_port, ZN => 
                           DATAPATH_I_N401);
   U1037 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_24_port, ZN => 
                           DATAPATH_I_N402);
   U1038 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_25_port, ZN => 
                           DATAPATH_I_N403);
   U1039 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_26_port, ZN => 
                           DATAPATH_I_N404);
   U1040 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_27_port, ZN => 
                           DATAPATH_I_N405);
   U1041 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_28_port, ZN => 
                           DATAPATH_I_N406);
   U1042 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_29_port, ZN => 
                           DATAPATH_I_N407);
   U1043 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_30_port, ZN => 
                           DATAPATH_I_N408);
   U1044 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_31_port, ZN => 
                           DATAPATH_I_N409);
   U1045 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_0_port, ZN => 
                           DATAPATH_I_N146);
   U1046 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_1_port, ZN => 
                           DATAPATH_I_N147);
   U1047 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_2_port, ZN => 
                           DATAPATH_I_N148);
   U1048 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_3_port, ZN => 
                           DATAPATH_I_N149);
   U1049 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_4_port, ZN => 
                           DATAPATH_I_N150);
   U1050 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_5_port, ZN => 
                           DATAPATH_I_N151);
   U1051 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_6_port, ZN => 
                           DATAPATH_I_N152);
   U1052 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_7_port, ZN => 
                           DATAPATH_I_N153);
   U1053 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_8_port, ZN => 
                           DATAPATH_I_N154);
   U1054 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_9_port, ZN => 
                           DATAPATH_I_N155);
   U1055 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_10_port, ZN => 
                           DATAPATH_I_N156);
   U1056 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_11_port, ZN => 
                           DATAPATH_I_N157);
   U1057 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_12_port, ZN => 
                           DATAPATH_I_N158);
   U1058 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_13_port, ZN => 
                           DATAPATH_I_N159);
   U1059 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_14_port, ZN => 
                           DATAPATH_I_N160);
   U1060 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_15_port, ZN => 
                           DATAPATH_I_N161);
   U1061 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_16_port, ZN => 
                           DATAPATH_I_N162);
   U1062 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_17_port, ZN => 
                           DATAPATH_I_N163);
   U1063 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_18_port, ZN => 
                           DATAPATH_I_N164);
   U1064 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_19_port, ZN => 
                           DATAPATH_I_N165);
   U1065 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_20_port, ZN => 
                           DATAPATH_I_N166);
   U1066 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_21_port, ZN => 
                           DATAPATH_I_N167);
   U1067 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_22_port, ZN => 
                           DATAPATH_I_N168);
   U1068 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_23_port, ZN => 
                           DATAPATH_I_N169);
   U1069 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_24_port, ZN => 
                           DATAPATH_I_N170);
   U1070 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_25_port, ZN => 
                           DATAPATH_I_N171);
   U1071 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_26_port, ZN => 
                           DATAPATH_I_N172);
   U1072 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_8_port, ZN => 
                           DATAPATH_I_N386);
   U1073 : AND2_X1 port map( A1 => RST, A2 => IR_30_port, ZN => DATAPATH_I_N64)
                           ;
   U1074 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_0_port, 
                           ZN => DATAPATH_I_N243);
   U1075 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_24_port,
                           ZN => DATAPATH_I_N267);
   U1076 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_9_port, 
                           ZN => DATAPATH_I_N252);
   U1077 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_1_port, 
                           ZN => DATAPATH_I_N244);
   U1078 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_7_port, 
                           ZN => DATAPATH_I_N250);
   U1079 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_15_port,
                           ZN => DATAPATH_I_N258);
   U1080 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_13_port,
                           ZN => DATAPATH_I_N256);
   U1081 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_5_port, 
                           ZN => DATAPATH_I_N248);
   U1082 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_12_port,
                           ZN => DATAPATH_I_N255);
   U1083 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_11_port,
                           ZN => DATAPATH_I_N254);
   U1084 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_4_port, 
                           ZN => DATAPATH_I_N247);
   U1085 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_25_port,
                           ZN => DATAPATH_I_N268);
   U1086 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_29_port,
                           ZN => DATAPATH_I_N272);
   U1087 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_31_port,
                           ZN => DATAPATH_I_N274);
   U1088 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_19_port,
                           ZN => DATAPATH_I_N262);
   U1089 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_16_port,
                           ZN => DATAPATH_I_N259);
   U1090 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_30_port,
                           ZN => DATAPATH_I_N273);
   U1091 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_2_port, 
                           ZN => DATAPATH_I_N245);
   U1092 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_21_port,
                           ZN => DATAPATH_I_N264);
   U1093 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_27_port,
                           ZN => DATAPATH_I_N270);
   U1094 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_14_port,
                           ZN => DATAPATH_I_N257);
   U1095 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_18_port,
                           ZN => DATAPATH_I_N261);
   U1096 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_3_port, 
                           ZN => DATAPATH_I_N246);
   U1097 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_26_port,
                           ZN => DATAPATH_I_N269);
   U1098 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_28_port,
                           ZN => DATAPATH_I_N271);
   U1099 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_6_port, 
                           ZN => DATAPATH_I_N249);
   U1100 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_17_port,
                           ZN => DATAPATH_I_N260);
   U1101 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_10_port,
                           ZN => DATAPATH_I_N253);
   U1102 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_23_port,
                           ZN => DATAPATH_I_N266);
   U1103 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_8_port, 
                           ZN => DATAPATH_I_N251);
   U1104 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_22_port,
                           ZN => DATAPATH_I_N265);
   U1105 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_20_port,
                           ZN => DATAPATH_I_N263);
   U1106 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_24_port, A2 => n318, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_3_port);
   U1107 : NOR2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_28_port, A2 => 
                           DATAPATH_I_IF_ID_IR_30_port, ZN => n322);
   U1108 : AND4_X1 port map( A1 => DATAPATH_I_IF_ID_IR_29_port, A2 => 
                           DATAPATH_I_IF_ID_IR_31_port, A3 => 
                           DATAPATH_I_IF_ID_IR_27_port, A4 => 
                           DATAPATH_I_IF_ID_IR_26_port, ZN => n321);
   U1109 : NOR3_X1 port map( A1 => DATAPATH_I_IF_ID_IR_28_port, A2 => 
                           DATAPATH_I_IF_ID_IR_29_port, A3 => 
                           DATAPATH_I_IF_ID_IR_31_port, ZN => n319);
   U1110 : NAND4_X1 port map( A1 => n440, A2 => n441, A3 => n442, A4 => n319, 
                           ZN => n346);
   U1111 : INV_X1 port map( A => n346, ZN => n320);
   U1112 : AOI21_X1 port map( B1 => n322, B2 => n321, A => n320, ZN => n323);
   U1113 : INV_X1 port map( A => n323, ZN => n345);
   U1114 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_20_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_4_port);
   U1115 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_18_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_2_port);
   U1116 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_17_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_1_port);
   U1117 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_16_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_0_port);
   U1118 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_19_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_3_port);
   U1119 : INV_X1 port map( A => IR_26_port, ZN => n387);
   U1120 : NOR2_X1 port map( A1 => n317, A2 => n387, ZN => DATAPATH_I_N60);
   U1121 : INV_X1 port map( A => IR_5_port, ZN => n384);
   U1122 : OR4_X1 port map( A1 => IR_6_port, A2 => IR_9_port, A3 => IR_7_port, 
                           A4 => IR_8_port, ZN => n324);
   U1123 : NOR2_X1 port map( A1 => IR_10_port, A2 => n324, ZN => n325);
   U1124 : INV_X1 port map( A => IR_4_port, ZN => n327);
   U1125 : NAND2_X1 port map( A1 => n325, A2 => n327, ZN => n329);
   U1126 : NOR2_X1 port map( A1 => n384, A2 => n329, ZN => n332);
   U1127 : INV_X1 port map( A => n332, ZN => n328);
   U1128 : NOR2_X1 port map( A1 => IR_1_port, A2 => n328, ZN => n367);
   U1129 : INV_X1 port map( A => IR_1_port, ZN => n370);
   U1130 : INV_X1 port map( A => IR_2_port, ZN => n330);
   U1131 : NAND2_X1 port map( A1 => n325, A2 => IR_3_port, ZN => n326);
   U1132 : NOR2_X1 port map( A1 => n327, A2 => n326, ZN => n385);
   U1133 : NAND2_X1 port map( A1 => IR_5_port, A2 => n385, ZN => n375);
   U1134 : AOI221_X1 port map( B1 => IR_1_port, B2 => IR_2_port, C1 => n370, C2
                           => n330, A => n375, ZN => n383);
   U1135 : AOI21_X1 port map( B1 => IR_3_port, B2 => n367, A => n383, ZN => 
                           n405);
   U1136 : NOR2_X1 port map( A1 => IR_31_port, A2 => IR_30_port, ZN => n362);
   U1137 : INV_X1 port map( A => IR_29_port, ZN => n357);
   U1138 : NAND2_X1 port map( A1 => n362, A2 => n357, ZN => n408);
   U1139 : NOR4_X1 port map( A1 => IR_28_port, A2 => IR_27_port, A3 => 
                           IR_26_port, A4 => n408, ZN => n439);
   U1140 : INV_X1 port map( A => IR_3_port, ZN => n366);
   U1141 : NAND2_X1 port map( A1 => n330, A2 => IR_1_port, ZN => n376);
   U1142 : NOR2_X1 port map( A1 => n376, A2 => n328, ZN => n371);
   U1143 : OR4_X1 port map( A1 => IR_5_port, A2 => IR_3_port, A3 => n330, A4 =>
                           n329, ZN => n372);
   U1144 : NOR2_X1 port map( A1 => n370, A2 => n372, ZN => n380);
   U1145 : AOI21_X1 port map( B1 => n366, B2 => n371, A => n380, ZN => n331);
   U1146 : INV_X1 port map( A => n331, ZN => n404);
   U1147 : INV_X1 port map( A => n367, ZN => n418);
   U1148 : NOR2_X1 port map( A1 => IR_2_port, A2 => n418, ZN => n382);
   U1149 : INV_X1 port map( A => IR_0_port, ZN => n421);
   U1150 : OAI211_X1 port map( C1 => n404, C2 => n382, A => n366, B => n421, ZN
                           => n334);
   U1151 : NAND3_X1 port map( A1 => IR_3_port, A2 => n371, A3 => IR_0_port, ZN 
                           => n333);
   U1152 : NAND4_X1 port map( A1 => IR_2_port, A2 => n332, A3 => n366, A4 => 
                           n421, ZN => n369);
   U1153 : AND4_X1 port map( A1 => n439, A2 => n334, A3 => n333, A4 => n369, ZN
                           => n344);
   U1154 : NAND2_X1 port map( A1 => IR_29_port, A2 => n362, ZN => n406);
   U1155 : INV_X1 port map( A => n406, ZN => n430);
   U1156 : INV_X1 port map( A => DATAPATH_I_N62, ZN => n398);
   U1157 : NOR4_X1 port map( A1 => IR_27_port, A2 => n408, A3 => n387, A4 => 
                           n398, ZN => n342);
   U1158 : INV_X1 port map( A => IR_27_port, ZN => n356);
   U1159 : NAND2_X1 port map( A1 => IR_28_port, A2 => n356, ZN => n427);
   U1160 : NAND3_X1 port map( A1 => IR_29_port, A2 => IR_31_port, A3 => 
                           IR_30_port, ZN => n389);
   U1161 : NOR2_X1 port map( A1 => n427, A2 => n389, ZN => n336);
   U1162 : INV_X1 port map( A => IR_31_port, ZN => n358);
   U1163 : NAND3_X1 port map( A1 => IR_29_port, A2 => IR_30_port, A3 => n358, 
                           ZN => n400);
   U1164 : NAND2_X1 port map( A1 => IR_27_port, A2 => n407, ZN => n411);
   U1165 : NOR2_X1 port map( A1 => n400, A2 => n411, ZN => n359);
   U1166 : NAND2_X1 port map( A1 => n356, A2 => n387, ZN => n399);
   U1167 : INV_X1 port map( A => n439, ZN => n335);
   U1168 : OAI21_X1 port map( B1 => n399, B2 => n400, A => n335, ZN => n379);
   U1169 : AOI221_X1 port map( B1 => n336, B2 => IR_26_port, C1 => n359, C2 => 
                           n387, A => n379, ZN => n340);
   U1170 : INV_X1 port map( A => n411, ZN => n360);
   U1171 : NAND2_X1 port map( A1 => IR_26_port, A2 => n360, ZN => n390);
   U1172 : NOR3_X1 port map( A1 => IR_30_port, A2 => n358, A3 => n390, ZN => 
                           n417);
   U1173 : AOI21_X1 port map( B1 => n408, B2 => n389, A => n390, ZN => n338);
   U1174 : NAND3_X1 port map( A1 => IR_30_port, A2 => n357, A3 => n358, ZN => 
                           n412);
   U1175 : NOR3_X1 port map( A1 => n407, A2 => n356, A3 => n412, ZN => n402);
   U1176 : INV_X1 port map( A => n402, ZN => n337);
   U1177 : OAI22_X1 port map( A1 => IR_26_port, A2 => n337, B1 => n412, B2 => 
                           n390, ZN => n391);
   U1178 : AOI211_X1 port map( C1 => n417, C2 => n357, A => n338, B => n391, ZN
                           => n339);
   U1179 : AOI21_X1 port map( B1 => n340, B2 => n339, A => n317, ZN => n341);
   U1180 : AOI211_X1 port map( C1 => n430, C2 => DATAPATH_I_N60, A => n342, B 
                           => n341, ZN => n343);
   U1181 : AOI221_X1 port map( B1 => n405, B2 => n344, C1 => n421, C2 => n344, 
                           A => n343, ZN => CU_I_aluOpcode1_0_port);
   DATAPATH_I_MEM_WB_RF_WE <= '0';
   U1183 : NOR3_X2 port map( A1 => n345, A2 => n317, A3 => n347, ZN => n353);
   U1184 : NOR2_X1 port map( A1 => n317, A2 => n346, ZN => n352);
   U1185 : AOI22_X1 port map( A1 => n353, A2 => DATAPATH_I_IF_ID_IR_16_port, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_11_port, ZN => 
                           n348);
   U1186 : NAND3_X1 port map( A1 => RST, A2 => n347, A3 => 
                           DATAPATH_I_IF_ID_IR_26_port, ZN => n354);
   U1187 : NAND2_X1 port map( A1 => n348, A2 => n354, ZN => DATAPATH_I_N109);
   U1188 : AOI22_X1 port map( A1 => n353, A2 => DATAPATH_I_IF_ID_IR_17_port, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_12_port, ZN => 
                           n349);
   U1189 : NAND2_X1 port map( A1 => n349, A2 => n354, ZN => DATAPATH_I_N110);
   U1190 : AOI22_X1 port map( A1 => n353, A2 => DATAPATH_I_IF_ID_IR_18_port, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_13_port, ZN => 
                           n350);
   U1191 : NAND2_X1 port map( A1 => n350, A2 => n354, ZN => DATAPATH_I_N111);
   U1192 : AOI22_X1 port map( A1 => n353, A2 => DATAPATH_I_IF_ID_IR_19_port, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_14_port, ZN => 
                           n351);
   U1193 : NAND2_X1 port map( A1 => n351, A2 => n354, ZN => DATAPATH_I_N112);
   U1194 : AOI22_X1 port map( A1 => n353, A2 => DATAPATH_I_IF_ID_IR_20_port, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_15_port, ZN => 
                           n355);
   U1195 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => DATAPATH_I_N113);
   U1196 : NOR2_X1 port map( A1 => n317, A2 => n356, ZN => DATAPATH_I_N61);
   U1197 : NOR2_X1 port map( A1 => n317, A2 => n357, ZN => DATAPATH_I_N63);
   U1198 : NOR2_X1 port map( A1 => n317, A2 => n358, ZN => DATAPATH_I_N65);
   U1199 : INV_X1 port map( A => n417, ZN => n365);
   U1200 : INV_X1 port map( A => n412, ZN => n388);
   U1201 : OAI221_X1 port map( B1 => IR_28_port, B2 => n388, C1 => n407, C2 => 
                           n430, A => IR_27_port, ZN => n424);
   U1202 : OAI21_X1 port map( B1 => n402, B2 => n359, A => IR_26_port, ZN => 
                           n364);
   U1203 : INV_X1 port map( A => n389, ZN => n361);
   U1204 : OAI21_X1 port map( B1 => n362, B2 => n361, A => n360, ZN => n363);
   U1205 : NAND4_X1 port map( A1 => n365, A2 => n424, A3 => n364, A4 => n363, 
                           ZN => n378);
   U1206 : NAND2_X1 port map( A1 => IR_0_port, A2 => n366, ZN => n381);
   U1207 : INV_X1 port map( A => n381, ZN => n373);
   U1208 : NAND3_X1 port map( A1 => IR_2_port, A2 => n373, A3 => n367, ZN => 
                           n368);
   U1209 : OAI21_X1 port map( B1 => n370, B2 => n369, A => n368, ZN => n397);
   U1210 : AOI21_X1 port map( B1 => n371, B2 => n381, A => n397, ZN => n419);
   U1211 : OAI21_X1 port map( B1 => IR_0_port, B2 => n372, A => n439, ZN => 
                           n403);
   U1212 : AOI21_X1 port map( B1 => n373, B2 => n382, A => n403, ZN => n374);
   U1213 : OAI211_X1 port map( C1 => n376, C2 => n375, A => n419, B => n374, ZN
                           => n377);
   U1214 : OAI211_X1 port map( C1 => n379, C2 => n378, A => RST, B => n377, ZN 
                           => CU_I_aluOpcode1_1_port);
   U1215 : AOI211_X1 port map( C1 => n382, C2 => n381, A => n380, B => n403, ZN
                           => n386);
   U1216 : INV_X1 port map( A => n383, ZN => n435);
   U1217 : NAND4_X1 port map( A1 => IR_1_port, A2 => IR_2_port, A3 => n385, A4 
                           => n384, ZN => n434);
   U1218 : NAND3_X1 port map( A1 => n386, A2 => n435, A3 => n434, ZN => n396);
   U1219 : OR2_X1 port map( A1 => n408, A2 => IR_27_port, ZN => n394);
   U1220 : NAND2_X1 port map( A1 => n427, A2 => n411, ZN => n429);
   U1221 : NAND2_X1 port map( A1 => n388, A2 => n387, ZN => n426);
   U1222 : NAND3_X1 port map( A1 => n406, A2 => n426, A3 => n389, ZN => n392);
   U1223 : AOI21_X1 port map( B1 => n427, B2 => n390, A => n400, ZN => n416);
   U1224 : AOI211_X1 port map( C1 => n429, C2 => n392, A => n416, B => n391, ZN
                           => n393);
   U1225 : OAI221_X1 port map( B1 => n394, B2 => IR_26_port, C1 => n394, C2 => 
                           n407, A => n393, ZN => n395);
   U1226 : OAI211_X1 port map( C1 => n397, C2 => n396, A => RST, B => n395, ZN 
                           => CU_I_aluOpcode1_2_port);
   U1227 : OR3_X1 port map( A1 => n399, A2 => n398, A3 => n412, ZN => n415);
   U1228 : AOI211_X1 port map( C1 => IR_27_port, C2 => IR_26_port, A => 
                           IR_28_port, B => n400, ZN => n401);
   U1229 : NOR2_X1 port map( A1 => n402, A2 => n401, ZN => n425);
   U1230 : NOR2_X1 port map( A1 => n404, A2 => n403, ZN => n420);
   U1231 : OAI211_X1 port map( C1 => IR_0_port, C2 => n434, A => n419, B => 
                           n405, ZN => n409);
   U1232 : AOI221_X1 port map( B1 => IR_28_port, B2 => n408, C1 => n407, C2 => 
                           n406, A => IR_27_port, ZN => n438);
   U1233 : AOI21_X1 port map( B1 => n420, B2 => n409, A => n438, ZN => n410);
   U1234 : OAI211_X1 port map( C1 => n412, C2 => n411, A => n425, B => n410, ZN
                           => n413);
   U1235 : AOI22_X1 port map( A1 => RST, A2 => n413, B1 => n417, B2 => 
                           DATAPATH_I_N63, ZN => n414);
   U1236 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => 
                           CU_I_aluOpcode1_3_port);
   U1237 : NOR2_X1 port map( A1 => n417, A2 => n416, ZN => n431);
   U1238 : AND3_X1 port map( A1 => n420, A2 => n419, A3 => n418, ZN => n436);
   U1239 : OAI21_X1 port map( B1 => n421, B2 => n434, A => n435, ZN => n422);
   U1240 : AOI21_X1 port map( B1 => n436, B2 => n422, A => n438, ZN => n423);
   U1241 : AOI21_X1 port map( B1 => n431, B2 => n423, A => n317, ZN => 
                           CU_I_aluOpcode1_4_port);
   U1242 : OAI211_X1 port map( C1 => n427, C2 => n426, A => n425, B => n424, ZN
                           => n428);
   U1243 : AOI211_X1 port map( C1 => n430, C2 => n429, A => n439, B => n428, ZN
                           => n432);
   U1244 : AOI22_X1 port map( A1 => n432, A2 => n431, B1 => n436, B2 => n435, 
                           ZN => n433);
   U1245 : NAND2_X1 port map( A1 => RST, A2 => n433, ZN => 
                           CU_I_aluOpcode1_5_port);
   U1246 : NAND3_X1 port map( A1 => n436, A2 => n435, A3 => n434, ZN => n437);
   U1247 : OAI211_X1 port map( C1 => n439, C2 => n438, A => RST, B => n437, ZN 
                           => CU_I_aluOpcode1_6_port);
   n285 <= '1';

end SYN_DLX_RTL;

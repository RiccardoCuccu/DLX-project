
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (OP_SLL, OP_SRL, OP_SRA, OP_ADD, OP_ADDU, OP_SUB, OP_SUBU, 
   OP_AND, OP_OR, OP_XOR, OP_SEQ, OP_SNE, OP_SLT, OP_SGT, OP_SLE, OP_SGE, 
   OP_MOVI2S, OP_MOVS2I, OP_MOVF, OP_MOVD, OP_MOVFP2I, OP_MOVI2FP, OP_MOVI2T, 
   OP_MOVT2I, OP_SLTU, OP_SGTU, OP_SLEU, OP_SGEU, OP_ADDF, OP_SUBF, OP_MULTF, 
   OP_DIVF, OP_ADDD, OP_SUBD, OP_MULTD, OP_DIVD, OP_CVTF2D, OP_CVTF2I, 
   OP_CVTD2F, OP_CVTD2I, OP_CVTI2F, OP_CVTI2D, OP_MULT, OP_DIV, OP_EQF, OP_NEF,
   OP_LTF, OP_GTF, OP_LEF, OP_GEF, OP_MULTU, OP_DIVU, OP_EQD, OP_NED, OP_LTD, 
   OP_GTD, OP_LED, OP_GED, OP_BEQZ, OP_BNEZ, OP_BFPT, OP_BFPF, OP_ADDI, 
   OP_ADDUI, OP_SUBI, OP_SUBUI, OP_ANDI, OP_ORI, OP_XORI, OP_LHI, OP_RFE, 
   OP_TRAP, OP_JR, OP_JALR, OP_SLLI, OP_SRLI, OP_SRAI, OP_SEQI, OP_SNEI, 
   OP_SLTI, OP_SGTI, OP_SLEI, OP_SGEI, OP_LB, OP_LH, OP_LW, OP_LBU, OP_LHU, 
   OP_LF, OP_LD, OP_SB, OP_SH, OP_SW, OP_SF, OP_SD, OP_ITLB, OP_SLTUI, 
   OP_SGTUI, OP_SLEUI, OP_SGEUI, OP_J, OP_JAL, OP_NOP);
attribute ENUM_ENCODING of aluOp : type is 
   "0000000 0000001 0000010 0000011 0000100 0000101 0000110 0000111 0001000 0001001 0001010 0001011 0001100 0001101 0001110 0001111 0010000 0010001 0010010 0010011 0010100 0010101 0010110 0010111 0011000 0011001 0011010 0011011 0011100 0011101 0011110 0011111 0100000 0100001 0100010 0100011 0100100 0100101 0100110 0100111 0101000 0101001 0101010 0101011 0101100 0101101 0101110 0101111 0110000 0110001 0110010 0110011 0110100 0110101 0110110 0110111 0111000 0111001 0111010 0111011 0111100 0111101 0111110 0111111 1000000 1000001 1000010 1000011 1000100 1000101 1000110 1000111 1001000 1001001 1001010 1001011 1001100 1001101 1001110 1001111 1010000 1010001 1010010 1010011 1010100 1010101 1010110 1010111 1011000 1011001 1011010 1011011 1011100 1011101 1011110 1011111 1100000 1100001 1100010 1100011 1100100 1100101 1100110";
   
   -- Declarations for conversion functions.
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when OP_SLL => return "0000000";
         when OP_SRL => return "0000001";
         when OP_SRA => return "0000010";
         when OP_ADD => return "0000011";
         when OP_ADDU => return "0000100";
         when OP_SUB => return "0000101";
         when OP_SUBU => return "0000110";
         when OP_AND => return "0000111";
         when OP_OR => return "0001000";
         when OP_XOR => return "0001001";
         when OP_SEQ => return "0001010";
         when OP_SNE => return "0001011";
         when OP_SLT => return "0001100";
         when OP_SGT => return "0001101";
         when OP_SLE => return "0001110";
         when OP_SGE => return "0001111";
         when OP_MOVI2S => return "0010000";
         when OP_MOVS2I => return "0010001";
         when OP_MOVF => return "0010010";
         when OP_MOVD => return "0010011";
         when OP_MOVFP2I => return "0010100";
         when OP_MOVI2FP => return "0010101";
         when OP_MOVI2T => return "0010110";
         when OP_MOVT2I => return "0010111";
         when OP_SLTU => return "0011000";
         when OP_SGTU => return "0011001";
         when OP_SLEU => return "0011010";
         when OP_SGEU => return "0011011";
         when OP_ADDF => return "0011100";
         when OP_SUBF => return "0011101";
         when OP_MULTF => return "0011110";
         when OP_DIVF => return "0011111";
         when OP_ADDD => return "0100000";
         when OP_SUBD => return "0100001";
         when OP_MULTD => return "0100010";
         when OP_DIVD => return "0100011";
         when OP_CVTF2D => return "0100100";
         when OP_CVTF2I => return "0100101";
         when OP_CVTD2F => return "0100110";
         when OP_CVTD2I => return "0100111";
         when OP_CVTI2F => return "0101000";
         when OP_CVTI2D => return "0101001";
         when OP_MULT => return "0101010";
         when OP_DIV => return "0101011";
         when OP_EQF => return "0101100";
         when OP_NEF => return "0101101";
         when OP_LTF => return "0101110";
         when OP_GTF => return "0101111";
         when OP_LEF => return "0110000";
         when OP_GEF => return "0110001";
         when OP_MULTU => return "0110010";
         when OP_DIVU => return "0110011";
         when OP_EQD => return "0110100";
         when OP_NED => return "0110101";
         when OP_LTD => return "0110110";
         when OP_GTD => return "0110111";
         when OP_LED => return "0111000";
         when OP_GED => return "0111001";
         when OP_BEQZ => return "0111010";
         when OP_BNEZ => return "0111011";
         when OP_BFPT => return "0111100";
         when OP_BFPF => return "0111101";
         when OP_ADDI => return "0111110";
         when OP_ADDUI => return "0111111";
         when OP_SUBI => return "1000000";
         when OP_SUBUI => return "1000001";
         when OP_ANDI => return "1000010";
         when OP_ORI => return "1000011";
         when OP_XORI => return "1000100";
         when OP_LHI => return "1000101";
         when OP_RFE => return "1000110";
         when OP_TRAP => return "1000111";
         when OP_JR => return "1001000";
         when OP_JALR => return "1001001";
         when OP_SLLI => return "1001010";
         when OP_SRLI => return "1001011";
         when OP_SRAI => return "1001100";
         when OP_SEQI => return "1001101";
         when OP_SNEI => return "1001110";
         when OP_SLTI => return "1001111";
         when OP_SGTI => return "1010000";
         when OP_SLEI => return "1010001";
         when OP_SGEI => return "1010010";
         when OP_LB => return "1010011";
         when OP_LH => return "1010100";
         when OP_LW => return "1010101";
         when OP_LBU => return "1010110";
         when OP_LHU => return "1010111";
         when OP_LF => return "1011000";
         when OP_LD => return "1011001";
         when OP_SB => return "1011010";
         when OP_SH => return "1011011";
         when OP_SW => return "1011100";
         when OP_SF => return "1011101";
         when OP_SD => return "1011110";
         when OP_ITLB => return "1011111";
         when OP_SLTUI => return "1100000";
         when OP_SGTUI => return "1100001";
         when OP_SLEUI => return "1100010";
         when OP_SGEUI => return "1100011";
         when OP_J => return "1100100";
         when OP_JAL => return "1100101";
         when OP_NOP => return "1100110";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

   port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  DOUT :
         out std_logic_vector (31 downto 0));

end DLX_IRAM_RAM_DEPTH256_I_SIZE32;

architecture SYN_BEHAVIORAL of DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_DRAM_N256_NW32 is

   port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector (31 
         downto 0);  DOUT : out std_logic_vector (31 downto 0));

end DLX_DRAM_N256_NW32;

architecture SYN_BEHAVIORAL of DLX_DRAM_N256_NW32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5;

architecture SYN_rpl of COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal GT_port, GE_port, NE_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, LE_port, n20, n21, n22, n23, n24, n25, n26,
      n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41
      , n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, 
      n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70
      , n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, 
      n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202 : std_logic;

begin
   GT <= GT_port;
   LE <= LE_port;
   GE <= GE_port;
   NE <= NE_port;
   
   U1 : INV_X1 port map( A => n154, ZN => n62);
   U2 : INV_X1 port map( A => NE_port, ZN => EQ);
   U3 : INV_X1 port map( A => n142, ZN => n58);
   U4 : INV_X1 port map( A => n130, ZN => n54);
   U5 : INV_X1 port map( A => n118, ZN => n50);
   U6 : INV_X1 port map( A => n106, ZN => n43);
   U7 : INV_X1 port map( A => n94, ZN => n35);
   U8 : INV_X1 port map( A => A(0), ZN => n2);
   U9 : INV_X1 port map( A => A(3), ZN => n4);
   U10 : INV_X1 port map( A => A(5), ZN => n6);
   U11 : INV_X1 port map( A => A(7), ZN => n8);
   U12 : INV_X1 port map( A => A(9), ZN => n10);
   U13 : INV_X1 port map( A => A(11), ZN => n12);
   U14 : INV_X1 port map( A => A(13), ZN => n14);
   U15 : INV_X1 port map( A => A(15), ZN => n16);
   U16 : INV_X1 port map( A => B(1), ZN => n1);
   U17 : INV_X1 port map( A => A(4), ZN => n5);
   U18 : INV_X1 port map( A => A(8), ZN => n9);
   U19 : INV_X1 port map( A => A(12), ZN => n13);
   U20 : INV_X1 port map( A => A(2), ZN => n3);
   U21 : INV_X1 port map( A => A(6), ZN => n7);
   U22 : INV_X1 port map( A => A(10), ZN => n11);
   U23 : INV_X1 port map( A => A(14), ZN => n15);
   U24 : INV_X1 port map( A => n82, ZN => n27);
   U25 : INV_X1 port map( A => n139, ZN => n57);
   U26 : INV_X1 port map( A => n127, ZN => n53);
   U27 : INV_X1 port map( A => n115, ZN => n49);
   U28 : INV_X1 port map( A => n103, ZN => n41);
   U29 : INV_X1 port map( A => n91, ZN => n33);
   U30 : INV_X1 port map( A => n79, ZN => n25);
   U31 : INV_X1 port map( A => n151, ZN => n61);
   U32 : INV_X1 port map( A => GT_port, ZN => LE_port);
   U33 : INV_X1 port map( A => n144, ZN => n60);
   U34 : INV_X1 port map( A => n132, ZN => n56);
   U35 : INV_X1 port map( A => n120, ZN => n52);
   U36 : INV_X1 port map( A => n141, ZN => n59);
   U37 : INV_X1 port map( A => n129, ZN => n55);
   U38 : INV_X1 port map( A => n117, ZN => n51);
   U39 : INV_X1 port map( A => n108, ZN => n46);
   U40 : INV_X1 port map( A => n96, ZN => n38);
   U41 : INV_X1 port map( A => n84, ZN => n30);
   U42 : INV_X1 port map( A => n105, ZN => n44);
   U43 : INV_X1 port map( A => n93, ZN => n36);
   U44 : INV_X1 port map( A => n81, ZN => n28);
   U45 : INV_X1 port map( A => n202, ZN => n63);
   U46 : INV_X1 port map( A => n68, ZN => n20);
   U47 : INV_X1 port map( A => n72, ZN => n22);
   U48 : INV_X1 port map( A => GE_port, ZN => LT);
   U49 : INV_X1 port map( A => A(30), ZN => n21);
   U50 : INV_X1 port map( A => A(17), ZN => n47);
   U51 : INV_X1 port map( A => A(21), ZN => n39);
   U52 : INV_X1 port map( A => A(25), ZN => n31);
   U53 : INV_X1 port map( A => A(29), ZN => n23);
   U54 : INV_X1 port map( A => A(16), ZN => n48);
   U55 : INV_X1 port map( A => A(20), ZN => n40);
   U56 : INV_X1 port map( A => A(24), ZN => n32);
   U57 : INV_X1 port map( A => A(28), ZN => n24);
   U58 : INV_X1 port map( A => A(18), ZN => n45);
   U59 : INV_X1 port map( A => A(22), ZN => n37);
   U60 : INV_X1 port map( A => A(26), ZN => n29);
   U61 : INV_X1 port map( A => A(19), ZN => n42);
   U62 : INV_X1 port map( A => A(23), ZN => n34);
   U63 : INV_X1 port map( A => A(27), ZN => n26);
   U64 : INV_X1 port map( A => B(30), ZN => n65);
   U65 : INV_X1 port map( A => B(31), ZN => n64);
   U66 : NAND2_X1 port map( A1 => LE_port, A2 => GE_port, ZN => NE_port);
   U67 : AOI21_X1 port map( B1 => n66, B2 => n20, A => n67, ZN => GE_port);
   U68 : AOI22_X1 port map( A1 => B(30), A2 => n21, B1 => n69, B2 => n70, ZN =>
                           n68);
   U69 : AOI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n69);
   U70 : AOI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n71);
   U71 : AOI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n74);
   U72 : AOI21_X1 port map( B1 => n80, B2 => n27, A => n28, ZN => n77);
   U73 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n80);
   U74 : AOI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n83);
   U75 : AOI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n86);
   U76 : AOI21_X1 port map( B1 => n92, B2 => n35, A => n36, ZN => n89);
   U77 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n92);
   U78 : AOI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n95);
   U79 : AOI21_X1 port map( B1 => n101, B2 => n102, A => n103, ZN => n98);
   U80 : AOI21_X1 port map( B1 => n104, B2 => n43, A => n44, ZN => n101);
   U81 : AOI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n104);
   U82 : AOI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n107);
   U83 : AOI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n110);
   U84 : AOI21_X1 port map( B1 => n116, B2 => n50, A => n51, ZN => n113);
   U85 : AOI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n116);
   U86 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n119);
   U87 : AOI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n122);
   U88 : AOI21_X1 port map( B1 => n128, B2 => n54, A => n55, ZN => n125);
   U89 : AOI21_X1 port map( B1 => n131, B2 => n132, A => n133, ZN => n128);
   U90 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n131);
   U91 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n134);
   U92 : AOI21_X1 port map( B1 => n140, B2 => n58, A => n59, ZN => n137);
   U93 : AOI21_X1 port map( B1 => n143, B2 => n144, A => n145, ZN => n140);
   U94 : AOI21_X1 port map( B1 => n146, B2 => n147, A => n148, ZN => n143);
   U95 : AOI21_X1 port map( B1 => n149, B2 => n150, A => n151, ZN => n146);
   U96 : AOI21_X1 port map( B1 => n152, B2 => n153, A => n62, ZN => n149);
   U97 : AOI22_X1 port map( A1 => n155, A2 => n1, B1 => A(1), B2 => n156, ZN =>
                           n152);
   U98 : OR2_X1 port map( A1 => n156, A2 => A(1), ZN => n155);
   U99 : NAND2_X1 port map( A1 => B(0), A2 => n2, ZN => n156);
   U100 : OAI21_X1 port map( B1 => n67, B2 => n157, A => n66, ZN => GT_port);
   U101 : NAND2_X1 port map( A1 => A(31), A2 => n64, ZN => n66);
   U102 : AOI22_X1 port map( A1 => A(30), A2 => n65, B1 => n158, B2 => n70, ZN 
                           => n157);
   U103 : XOR2_X1 port map( A => A(30), B => n65, Z => n70);
   U104 : AOI21_X1 port map( B1 => n159, B2 => n160, A => n22, ZN => n158);
   U105 : NAND2_X1 port map( A1 => B(29), A2 => n23, ZN => n72);
   U106 : OAI211_X1 port map( C1 => n161, C2 => n162, A => n78, B => n75, ZN =>
                           n160);
   U107 : NOR2_X1 port map( A1 => n163, A2 => n76, ZN => n75);
   U108 : AND2_X1 port map( A1 => B(28), A2 => n24, ZN => n76);
   U109 : NAND2_X1 port map( A1 => B(27), A2 => n26, ZN => n78);
   U110 : NAND2_X1 port map( A1 => n25, A2 => n164, ZN => n162);
   U111 : NOR2_X1 port map( A1 => n26, A2 => B(27), ZN => n79);
   U112 : AOI211_X1 port map( C1 => n165, C2 => n166, A => n82, B => n30, ZN =>
                           n161);
   U113 : NAND2_X1 port map( A1 => B(25), A2 => n31, ZN => n84);
   U114 : NAND2_X1 port map( A1 => n164, A2 => n81, ZN => n82);
   U115 : NAND2_X1 port map( A1 => B(26), A2 => n29, ZN => n81);
   U116 : OR2_X1 port map( A1 => n29, A2 => B(26), ZN => n164);
   U117 : OAI211_X1 port map( C1 => n167, C2 => n168, A => n90, B => n87, ZN =>
                           n166);
   U118 : NOR2_X1 port map( A1 => n169, A2 => n88, ZN => n87);
   U119 : AND2_X1 port map( A1 => B(24), A2 => n32, ZN => n88);
   U120 : NAND2_X1 port map( A1 => B(23), A2 => n34, ZN => n90);
   U121 : NAND2_X1 port map( A1 => n33, A2 => n170, ZN => n168);
   U122 : NOR2_X1 port map( A1 => n34, A2 => B(23), ZN => n91);
   U123 : AOI211_X1 port map( C1 => n171, C2 => n172, A => n94, B => n38, ZN =>
                           n167);
   U124 : NAND2_X1 port map( A1 => B(21), A2 => n39, ZN => n96);
   U125 : NAND2_X1 port map( A1 => n170, A2 => n93, ZN => n94);
   U126 : NAND2_X1 port map( A1 => B(22), A2 => n37, ZN => n93);
   U127 : OR2_X1 port map( A1 => n37, A2 => B(22), ZN => n170);
   U128 : OAI211_X1 port map( C1 => n173, C2 => n174, A => n102, B => n99, ZN 
                           => n172);
   U129 : NOR2_X1 port map( A1 => n175, A2 => n100, ZN => n99);
   U130 : AND2_X1 port map( A1 => B(20), A2 => n40, ZN => n100);
   U131 : NAND2_X1 port map( A1 => B(19), A2 => n42, ZN => n102);
   U132 : NAND2_X1 port map( A1 => n41, A2 => n176, ZN => n174);
   U133 : NOR2_X1 port map( A1 => n42, A2 => B(19), ZN => n103);
   U134 : AOI211_X1 port map( C1 => n177, C2 => n178, A => n106, B => n46, ZN 
                           => n173);
   U135 : NAND2_X1 port map( A1 => B(17), A2 => n47, ZN => n108);
   U136 : NAND2_X1 port map( A1 => n176, A2 => n105, ZN => n106);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n45, ZN => n105);
   U138 : OR2_X1 port map( A1 => n45, A2 => B(18), ZN => n176);
   U139 : OAI211_X1 port map( C1 => n179, C2 => n180, A => n114, B => n111, ZN 
                           => n178);
   U140 : NOR2_X1 port map( A1 => n181, A2 => n112, ZN => n111);
   U141 : AND2_X1 port map( A1 => B(16), A2 => n48, ZN => n112);
   U142 : NAND2_X1 port map( A1 => B(15), A2 => n16, ZN => n114);
   U143 : NAND2_X1 port map( A1 => n49, A2 => n182, ZN => n180);
   U144 : NOR2_X1 port map( A1 => n16, A2 => B(15), ZN => n115);
   U145 : AOI211_X1 port map( C1 => n183, C2 => n184, A => n118, B => n52, ZN 
                           => n179);
   U146 : NAND2_X1 port map( A1 => B(13), A2 => n14, ZN => n120);
   U147 : NAND2_X1 port map( A1 => n182, A2 => n117, ZN => n118);
   U148 : NAND2_X1 port map( A1 => B(14), A2 => n15, ZN => n117);
   U149 : OR2_X1 port map( A1 => n15, A2 => B(14), ZN => n182);
   U150 : OAI211_X1 port map( C1 => n185, C2 => n186, A => n126, B => n123, ZN 
                           => n184);
   U151 : NOR2_X1 port map( A1 => n187, A2 => n124, ZN => n123);
   U152 : AND2_X1 port map( A1 => B(12), A2 => n13, ZN => n124);
   U153 : NAND2_X1 port map( A1 => B(11), A2 => n12, ZN => n126);
   U154 : NAND2_X1 port map( A1 => n53, A2 => n188, ZN => n186);
   U155 : NOR2_X1 port map( A1 => n12, A2 => B(11), ZN => n127);
   U156 : AOI211_X1 port map( C1 => n189, C2 => n190, A => n130, B => n56, ZN 
                           => n185);
   U157 : NAND2_X1 port map( A1 => B(9), A2 => n10, ZN => n132);
   U158 : NAND2_X1 port map( A1 => n188, A2 => n129, ZN => n130);
   U159 : NAND2_X1 port map( A1 => B(10), A2 => n11, ZN => n129);
   U160 : OR2_X1 port map( A1 => n11, A2 => B(10), ZN => n188);
   U161 : OAI211_X1 port map( C1 => n191, C2 => n192, A => n138, B => n135, ZN 
                           => n190);
   U162 : NOR2_X1 port map( A1 => n193, A2 => n136, ZN => n135);
   U163 : AND2_X1 port map( A1 => B(8), A2 => n9, ZN => n136);
   U164 : NAND2_X1 port map( A1 => B(7), A2 => n8, ZN => n138);
   U165 : NAND2_X1 port map( A1 => n57, A2 => n194, ZN => n192);
   U166 : NOR2_X1 port map( A1 => n8, A2 => B(7), ZN => n139);
   U167 : AOI211_X1 port map( C1 => n195, C2 => n196, A => n142, B => n60, ZN 
                           => n191);
   U168 : NAND2_X1 port map( A1 => B(5), A2 => n6, ZN => n144);
   U169 : NAND2_X1 port map( A1 => n194, A2 => n141, ZN => n142);
   U170 : NAND2_X1 port map( A1 => B(6), A2 => n7, ZN => n141);
   U171 : OR2_X1 port map( A1 => n7, A2 => B(6), ZN => n194);
   U172 : NAND3_X1 port map( A1 => n197, A2 => n150, A3 => n147, ZN => n196);
   U173 : NOR2_X1 port map( A1 => n198, A2 => n148, ZN => n147);
   U174 : AND2_X1 port map( A1 => B(4), A2 => n5, ZN => n148);
   U175 : NAND2_X1 port map( A1 => B(3), A2 => n4, ZN => n150);
   U176 : NAND3_X1 port map( A1 => n61, A2 => n199, A3 => n200, ZN => n197);
   U177 : OAI211_X1 port map( C1 => A(1), C2 => n201, A => n63, B => n153, ZN 
                           => n200);
   U178 : AND2_X1 port map( A1 => n199, A2 => n154, ZN => n153);
   U179 : NAND2_X1 port map( A1 => B(2), A2 => n3, ZN => n154);
   U180 : AOI21_X1 port map( B1 => A(1), B2 => n201, A => n1, ZN => n202);
   U181 : NOR2_X1 port map( A1 => n2, A2 => B(0), ZN => n201);
   U182 : OR2_X1 port map( A1 => n3, A2 => B(2), ZN => n199);
   U183 : NOR2_X1 port map( A1 => n4, A2 => B(3), ZN => n151);
   U184 : NOR2_X1 port map( A1 => n198, A2 => n145, ZN => n195);
   U185 : NOR2_X1 port map( A1 => n6, A2 => B(5), ZN => n145);
   U186 : NOR2_X1 port map( A1 => n5, A2 => B(4), ZN => n198);
   U187 : NOR2_X1 port map( A1 => n193, A2 => n133, ZN => n189);
   U188 : NOR2_X1 port map( A1 => n10, A2 => B(9), ZN => n133);
   U189 : NOR2_X1 port map( A1 => n9, A2 => B(8), ZN => n193);
   U190 : NOR2_X1 port map( A1 => n187, A2 => n121, ZN => n183);
   U191 : NOR2_X1 port map( A1 => n14, A2 => B(13), ZN => n121);
   U192 : NOR2_X1 port map( A1 => n13, A2 => B(12), ZN => n187);
   U193 : NOR2_X1 port map( A1 => n181, A2 => n109, ZN => n177);
   U194 : NOR2_X1 port map( A1 => n47, A2 => B(17), ZN => n109);
   U195 : NOR2_X1 port map( A1 => n48, A2 => B(16), ZN => n181);
   U196 : NOR2_X1 port map( A1 => n175, A2 => n97, ZN => n171);
   U197 : NOR2_X1 port map( A1 => n39, A2 => B(21), ZN => n97);
   U198 : NOR2_X1 port map( A1 => n40, A2 => B(20), ZN => n175);
   U199 : NOR2_X1 port map( A1 => n169, A2 => n85, ZN => n165);
   U200 : NOR2_X1 port map( A1 => n31, A2 => B(25), ZN => n85);
   U201 : NOR2_X1 port map( A1 => n32, A2 => B(24), ZN => n169);
   U202 : NOR2_X1 port map( A1 => n163, A2 => n73, ZN => n159);
   U203 : NOR2_X1 port map( A1 => n23, A2 => B(29), ZN => n73);
   U204 : NOR2_X1 port map( A1 => n24, A2 => B(28), ZN => n163);
   U205 : NOR2_X1 port map( A1 => n64, A2 => A(31), ZN => n67);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4;

architecture SYN_rpl of COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal LT_port, LE_port, n1, n2, n3, n4, n5, n6, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203 : std_logic;

begin
   LT <= LT_port;
   LE <= LE_port;
   
   U1 : INV_X1 port map( A => n139, ZN => n37);
   U2 : INV_X1 port map( A => n138, ZN => n36);
   U3 : INV_X1 port map( A => n123, ZN => n29);
   U4 : INV_X1 port map( A => n133, ZN => n33);
   U5 : INV_X1 port map( A => n134, ZN => n35);
   U6 : INV_X1 port map( A => n124, ZN => n31);
   U7 : INV_X1 port map( A => n119, ZN => n28);
   U8 : INV_X1 port map( A => n113, ZN => n25);
   U9 : INV_X1 port map( A => n114, ZN => n27);
   U10 : INV_X1 port map( A => n143, ZN => n39);
   U11 : INV_X1 port map( A => n195, ZN => n34);
   U12 : INV_X1 port map( A => n189, ZN => n30);
   U13 : INV_X1 port map( A => n183, ZN => n26);
   U14 : INV_X1 port map( A => n201, ZN => n38);
   U15 : INV_X1 port map( A => n103, ZN => n21);
   U16 : INV_X1 port map( A => n83, ZN => n13);
   U17 : INV_X1 port map( A => n129, ZN => n32);
   U18 : INV_X1 port map( A => n109, ZN => n24);
   U19 : INV_X1 port map( A => n5, ZN => n6);
   U20 : INV_X1 port map( A => B(0), ZN => n1);
   U21 : INV_X1 port map( A => B(2), ZN => n2);
   U22 : INV_X1 port map( A => B(4), ZN => n4);
   U23 : INV_X1 port map( A => B(3), ZN => n3);
   U24 : INV_X1 port map( A => n93, ZN => n17);
   U25 : INV_X1 port map( A => n94, ZN => n19);
   U26 : INV_X1 port map( A => n99, ZN => n20);
   U27 : INV_X1 port map( A => n79, ZN => n12);
   U28 : INV_X1 port map( A => n104, ZN => n23);
   U29 : INV_X1 port map( A => n84, ZN => n15);
   U30 : INV_X1 port map( A => n177, ZN => n22);
   U31 : INV_X1 port map( A => n171, ZN => n18);
   U32 : INV_X1 port map( A => n165, ZN => n14);
   U33 : INV_X1 port map( A => n89, ZN => n16);
   U34 : BUF_X1 port map( A => A(1), Z => n5);
   U35 : INV_X1 port map( A => n69, ZN => n9);
   U36 : INV_X1 port map( A => B(30), ZN => n41);
   U37 : INV_X1 port map( A => n74, ZN => n11);
   U38 : INV_X1 port map( A => LE_port, ZN => GT);
   U39 : INV_X1 port map( A => A(30), ZN => n10);
   U40 : INV_X1 port map( A => LT_port, ZN => GE);
   U41 : INV_X1 port map( A => B(5), ZN => n66);
   U42 : INV_X1 port map( A => B(9), ZN => n62);
   U43 : INV_X1 port map( A => B(13), ZN => n58);
   U44 : INV_X1 port map( A => B(8), ZN => n63);
   U45 : INV_X1 port map( A => B(12), ZN => n59);
   U46 : INV_X1 port map( A => B(7), ZN => n64);
   U47 : INV_X1 port map( A => B(11), ZN => n60);
   U48 : INV_X1 port map( A => B(15), ZN => n56);
   U49 : INV_X1 port map( A => B(16), ZN => n55);
   U50 : INV_X1 port map( A => B(20), ZN => n51);
   U51 : INV_X1 port map( A => B(24), ZN => n47);
   U52 : INV_X1 port map( A => B(28), ZN => n43);
   U53 : INV_X1 port map( A => B(6), ZN => n65);
   U54 : INV_X1 port map( A => B(10), ZN => n61);
   U55 : INV_X1 port map( A => B(14), ZN => n57);
   U56 : INV_X1 port map( A => B(18), ZN => n53);
   U57 : INV_X1 port map( A => B(22), ZN => n49);
   U58 : INV_X1 port map( A => B(26), ZN => n45);
   U59 : INV_X1 port map( A => B(31), ZN => n40);
   U60 : INV_X1 port map( A => B(17), ZN => n54);
   U61 : INV_X1 port map( A => B(21), ZN => n50);
   U62 : INV_X1 port map( A => B(25), ZN => n46);
   U63 : INV_X1 port map( A => B(29), ZN => n42);
   U64 : INV_X1 port map( A => B(19), ZN => n52);
   U65 : INV_X1 port map( A => B(23), ZN => n48);
   U66 : INV_X1 port map( A => B(27), ZN => n44);
   U67 : AOI21_X1 port map( B1 => n67, B2 => n9, A => n68, ZN => LE_port);
   U68 : AOI22_X1 port map( A1 => A(30), A2 => n41, B1 => n70, B2 => n71, ZN =>
                           n69);
   U69 : AOI21_X1 port map( B1 => n72, B2 => n73, A => n74, ZN => n70);
   U70 : OAI211_X1 port map( C1 => n75, C2 => n76, A => n77, B => n78, ZN => 
                           n73);
   U71 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n76);
   U72 : AOI211_X1 port map( C1 => n81, C2 => n82, A => n83, B => n84, ZN => 
                           n75);
   U73 : OAI211_X1 port map( C1 => n85, C2 => n86, A => n87, B => n88, ZN => 
                           n82);
   U74 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => n86);
   U75 : AOI211_X1 port map( C1 => n91, C2 => n92, A => n93, B => n94, ZN => 
                           n85);
   U76 : OAI211_X1 port map( C1 => n95, C2 => n96, A => n97, B => n98, ZN => 
                           n92);
   U77 : NAND2_X1 port map( A1 => n99, A2 => n100, ZN => n96);
   U78 : AOI211_X1 port map( C1 => n101, C2 => n102, A => n103, B => n104, ZN 
                           => n95);
   U79 : OAI211_X1 port map( C1 => n105, C2 => n106, A => n107, B => n108, ZN 
                           => n102);
   U80 : NAND2_X1 port map( A1 => n109, A2 => n110, ZN => n106);
   U81 : AOI211_X1 port map( C1 => n111, C2 => n112, A => n113, B => n114, ZN 
                           => n105);
   U82 : OAI211_X1 port map( C1 => n115, C2 => n116, A => n117, B => n118, ZN 
                           => n112);
   U83 : NAND2_X1 port map( A1 => n119, A2 => n120, ZN => n116);
   U84 : AOI211_X1 port map( C1 => n121, C2 => n122, A => n123, B => n124, ZN 
                           => n115);
   U85 : OAI211_X1 port map( C1 => n125, C2 => n126, A => n127, B => n128, ZN 
                           => n122);
   U86 : NAND2_X1 port map( A1 => n129, A2 => n130, ZN => n126);
   U87 : AOI211_X1 port map( C1 => n131, C2 => n132, A => n133, B => n134, ZN 
                           => n125);
   U88 : NAND3_X1 port map( A1 => n135, A2 => n136, A3 => n137, ZN => n132);
   U89 : NAND3_X1 port map( A1 => n138, A2 => n139, A3 => n140, ZN => n135);
   U90 : OAI211_X1 port map( C1 => n5, C2 => n39, A => n141, B => n142, ZN => 
                           n140);
   U91 : OAI21_X1 port map( B1 => n6, B2 => n143, A => B(1), ZN => n141);
   U92 : NAND2_X1 port map( A1 => A(0), A2 => n1, ZN => n143);
   U93 : NOR2_X1 port map( A1 => n144, A2 => n145, ZN => n131);
   U94 : NOR2_X1 port map( A1 => n146, A2 => n147, ZN => n121);
   U95 : NOR2_X1 port map( A1 => n148, A2 => n149, ZN => n111);
   U96 : NOR2_X1 port map( A1 => n150, A2 => n151, ZN => n101);
   U97 : NOR2_X1 port map( A1 => n152, A2 => n153, ZN => n91);
   U98 : NOR2_X1 port map( A1 => n154, A2 => n155, ZN => n81);
   U99 : NOR2_X1 port map( A1 => n156, A2 => n157, ZN => n72);
   U100 : OAI21_X1 port map( B1 => n68, B2 => n158, A => n67, ZN => LT_port);
   U101 : NAND2_X1 port map( A1 => A(31), A2 => n40, ZN => n67);
   U102 : AOI22_X1 port map( A1 => B(30), A2 => n10, B1 => n159, B2 => n71, ZN 
                           => n158);
   U103 : XOR2_X1 port map( A => n10, B => B(30), Z => n71);
   U104 : AOI21_X1 port map( B1 => n160, B2 => n11, A => n157, ZN => n159);
   U105 : AND2_X1 port map( A1 => A(29), A2 => n42, ZN => n157);
   U106 : NOR2_X1 port map( A1 => n42, A2 => A(29), ZN => n74);
   U107 : AOI21_X1 port map( B1 => n161, B2 => n78, A => n162, ZN => n160);
   U108 : NOR2_X1 port map( A1 => n162, A2 => n156, ZN => n78);
   U109 : AND2_X1 port map( A1 => A(28), A2 => n43, ZN => n156);
   U110 : NOR2_X1 port map( A1 => n43, A2 => A(28), ZN => n162);
   U111 : AOI21_X1 port map( B1 => n163, B2 => n77, A => n12, ZN => n161);
   U112 : NAND2_X1 port map( A1 => A(27), A2 => n44, ZN => n79);
   U113 : OR2_X1 port map( A1 => n44, A2 => A(27), ZN => n77);
   U114 : AOI21_X1 port map( B1 => n164, B2 => n13, A => n165, ZN => n163);
   U115 : NAND2_X1 port map( A1 => n14, A2 => n80, ZN => n83);
   U116 : NAND2_X1 port map( A1 => A(26), A2 => n45, ZN => n80);
   U117 : NOR2_X1 port map( A1 => n45, A2 => A(26), ZN => n165);
   U118 : AOI21_X1 port map( B1 => n166, B2 => n15, A => n155, ZN => n164);
   U119 : AND2_X1 port map( A1 => A(25), A2 => n46, ZN => n155);
   U120 : NOR2_X1 port map( A1 => n46, A2 => A(25), ZN => n84);
   U121 : AOI21_X1 port map( B1 => n167, B2 => n88, A => n168, ZN => n166);
   U122 : NOR2_X1 port map( A1 => n168, A2 => n154, ZN => n88);
   U123 : AND2_X1 port map( A1 => A(24), A2 => n47, ZN => n154);
   U124 : NOR2_X1 port map( A1 => n47, A2 => A(24), ZN => n168);
   U125 : AOI21_X1 port map( B1 => n169, B2 => n87, A => n16, ZN => n167);
   U126 : NAND2_X1 port map( A1 => A(23), A2 => n48, ZN => n89);
   U127 : OR2_X1 port map( A1 => n48, A2 => A(23), ZN => n87);
   U128 : AOI21_X1 port map( B1 => n170, B2 => n17, A => n171, ZN => n169);
   U129 : NAND2_X1 port map( A1 => n18, A2 => n90, ZN => n93);
   U130 : NAND2_X1 port map( A1 => A(22), A2 => n49, ZN => n90);
   U131 : NOR2_X1 port map( A1 => n49, A2 => A(22), ZN => n171);
   U132 : AOI21_X1 port map( B1 => n172, B2 => n19, A => n153, ZN => n170);
   U133 : AND2_X1 port map( A1 => A(21), A2 => n50, ZN => n153);
   U134 : NOR2_X1 port map( A1 => n50, A2 => A(21), ZN => n94);
   U135 : AOI21_X1 port map( B1 => n173, B2 => n98, A => n174, ZN => n172);
   U136 : NOR2_X1 port map( A1 => n174, A2 => n152, ZN => n98);
   U137 : AND2_X1 port map( A1 => A(20), A2 => n51, ZN => n152);
   U138 : NOR2_X1 port map( A1 => n51, A2 => A(20), ZN => n174);
   U139 : AOI21_X1 port map( B1 => n175, B2 => n97, A => n20, ZN => n173);
   U140 : NAND2_X1 port map( A1 => A(19), A2 => n52, ZN => n99);
   U141 : OR2_X1 port map( A1 => n52, A2 => A(19), ZN => n97);
   U142 : AOI21_X1 port map( B1 => n176, B2 => n21, A => n177, ZN => n175);
   U143 : NAND2_X1 port map( A1 => n22, A2 => n100, ZN => n103);
   U144 : NAND2_X1 port map( A1 => A(18), A2 => n53, ZN => n100);
   U145 : NOR2_X1 port map( A1 => n53, A2 => A(18), ZN => n177);
   U146 : AOI21_X1 port map( B1 => n178, B2 => n23, A => n151, ZN => n176);
   U147 : AND2_X1 port map( A1 => A(17), A2 => n54, ZN => n151);
   U148 : NOR2_X1 port map( A1 => n54, A2 => A(17), ZN => n104);
   U149 : AOI21_X1 port map( B1 => n179, B2 => n108, A => n180, ZN => n178);
   U150 : NOR2_X1 port map( A1 => n180, A2 => n150, ZN => n108);
   U151 : AND2_X1 port map( A1 => A(16), A2 => n55, ZN => n150);
   U152 : NOR2_X1 port map( A1 => n55, A2 => A(16), ZN => n180);
   U153 : AOI21_X1 port map( B1 => n181, B2 => n107, A => n24, ZN => n179);
   U154 : NAND2_X1 port map( A1 => A(15), A2 => n56, ZN => n109);
   U155 : OR2_X1 port map( A1 => n56, A2 => A(15), ZN => n107);
   U156 : AOI21_X1 port map( B1 => n182, B2 => n25, A => n183, ZN => n181);
   U157 : NAND2_X1 port map( A1 => n26, A2 => n110, ZN => n113);
   U158 : NAND2_X1 port map( A1 => A(14), A2 => n57, ZN => n110);
   U159 : NOR2_X1 port map( A1 => n57, A2 => A(14), ZN => n183);
   U160 : AOI21_X1 port map( B1 => n184, B2 => n27, A => n149, ZN => n182);
   U161 : AND2_X1 port map( A1 => A(13), A2 => n58, ZN => n149);
   U162 : NOR2_X1 port map( A1 => n58, A2 => A(13), ZN => n114);
   U163 : AOI21_X1 port map( B1 => n185, B2 => n118, A => n186, ZN => n184);
   U164 : NOR2_X1 port map( A1 => n186, A2 => n148, ZN => n118);
   U165 : AND2_X1 port map( A1 => A(12), A2 => n59, ZN => n148);
   U166 : NOR2_X1 port map( A1 => n59, A2 => A(12), ZN => n186);
   U167 : AOI21_X1 port map( B1 => n187, B2 => n117, A => n28, ZN => n185);
   U168 : NAND2_X1 port map( A1 => A(11), A2 => n60, ZN => n119);
   U169 : OR2_X1 port map( A1 => n60, A2 => A(11), ZN => n117);
   U170 : AOI21_X1 port map( B1 => n188, B2 => n29, A => n189, ZN => n187);
   U171 : NAND2_X1 port map( A1 => n30, A2 => n120, ZN => n123);
   U172 : NAND2_X1 port map( A1 => A(10), A2 => n61, ZN => n120);
   U173 : NOR2_X1 port map( A1 => n61, A2 => A(10), ZN => n189);
   U174 : AOI21_X1 port map( B1 => n190, B2 => n31, A => n147, ZN => n188);
   U175 : AND2_X1 port map( A1 => A(9), A2 => n62, ZN => n147);
   U176 : NOR2_X1 port map( A1 => n62, A2 => A(9), ZN => n124);
   U177 : AOI21_X1 port map( B1 => n191, B2 => n128, A => n192, ZN => n190);
   U178 : NOR2_X1 port map( A1 => n192, A2 => n146, ZN => n128);
   U179 : AND2_X1 port map( A1 => A(8), A2 => n63, ZN => n146);
   U180 : NOR2_X1 port map( A1 => n63, A2 => A(8), ZN => n192);
   U181 : AOI21_X1 port map( B1 => n193, B2 => n127, A => n32, ZN => n191);
   U182 : NAND2_X1 port map( A1 => A(7), A2 => n64, ZN => n129);
   U183 : OR2_X1 port map( A1 => n64, A2 => A(7), ZN => n127);
   U184 : AOI21_X1 port map( B1 => n194, B2 => n33, A => n195, ZN => n193);
   U185 : NAND2_X1 port map( A1 => n34, A2 => n130, ZN => n133);
   U186 : NAND2_X1 port map( A1 => A(6), A2 => n65, ZN => n130);
   U187 : NOR2_X1 port map( A1 => n65, A2 => A(6), ZN => n195);
   U188 : AOI21_X1 port map( B1 => n196, B2 => n35, A => n145, ZN => n194);
   U189 : AND2_X1 port map( A1 => A(5), A2 => n66, ZN => n145);
   U190 : NOR2_X1 port map( A1 => n66, A2 => A(5), ZN => n134);
   U191 : AOI21_X1 port map( B1 => n197, B2 => n137, A => n198, ZN => n196);
   U192 : NOR2_X1 port map( A1 => n198, A2 => n144, ZN => n137);
   U193 : AND2_X1 port map( A1 => A(4), A2 => n4, ZN => n144);
   U194 : NOR2_X1 port map( A1 => n4, A2 => A(4), ZN => n198);
   U195 : AOI21_X1 port map( B1 => n199, B2 => n136, A => n36, ZN => n197);
   U196 : NAND2_X1 port map( A1 => A(3), A2 => n3, ZN => n138);
   U197 : OR2_X1 port map( A1 => n3, A2 => A(3), ZN => n136);
   U198 : AOI21_X1 port map( B1 => n38, B2 => n142, A => n200, ZN => n199);
   U199 : NOR2_X1 port map( A1 => n200, A2 => n37, ZN => n142);
   U200 : NAND2_X1 port map( A1 => A(2), A2 => n2, ZN => n139);
   U201 : NOR2_X1 port map( A1 => n2, A2 => A(2), ZN => n200);
   U202 : OAI22_X1 port map( A1 => n202, A2 => B(1), B1 => n6, B2 => n203, ZN 
                           => n201);
   U203 : AND2_X1 port map( A1 => n203, A2 => n6, ZN => n202);
   U204 : NOR2_X1 port map( A1 => n1, A2 => A(0), ZN => n203);
   U205 : NOR2_X1 port map( A1 => n40, A2 => A(31), ZN => n68);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity 
   DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0 
   is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0
   ;

architecture SYN_rpl of 
   DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0 
   is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_3_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_8_port, SUM_7_port, SUM_6_port, SUM_5_port,
      SUM_4_port, SUM_31_port, SUM_9_port, n30, n31, n32, n33, n34, n35, n36, 
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U2 : XOR2_X1 port map( A => A(30), B => n30, Z => SUM_30_port);
   U3 : XOR2_X1 port map( A => A(29), B => n31, Z => SUM_29_port);
   U4 : XOR2_X1 port map( A => A(28), B => n32, Z => SUM_28_port);
   U5 : XOR2_X1 port map( A => A(27), B => n33, Z => SUM_27_port);
   U6 : XOR2_X1 port map( A => A(26), B => n34, Z => SUM_26_port);
   U7 : XOR2_X1 port map( A => A(25), B => n35, Z => SUM_25_port);
   U8 : XOR2_X1 port map( A => A(24), B => n36, Z => SUM_24_port);
   U9 : XOR2_X1 port map( A => A(23), B => n37, Z => SUM_23_port);
   U10 : XOR2_X1 port map( A => A(22), B => n38, Z => SUM_22_port);
   U11 : XOR2_X1 port map( A => A(21), B => n39, Z => SUM_21_port);
   U12 : XOR2_X1 port map( A => A(20), B => n40, Z => SUM_20_port);
   U13 : XOR2_X1 port map( A => A(19), B => n41, Z => SUM_19_port);
   U14 : XOR2_X1 port map( A => A(18), B => n42, Z => SUM_18_port);
   U15 : XOR2_X1 port map( A => A(17), B => n43, Z => SUM_17_port);
   U16 : XOR2_X1 port map( A => A(16), B => n44, Z => SUM_16_port);
   U17 : XOR2_X1 port map( A => A(15), B => n45, Z => SUM_15_port);
   U18 : XOR2_X1 port map( A => A(14), B => n46, Z => SUM_14_port);
   U19 : XOR2_X1 port map( A => A(13), B => n47, Z => SUM_13_port);
   U20 : XOR2_X1 port map( A => A(12), B => n48, Z => SUM_12_port);
   U21 : XOR2_X1 port map( A => A(11), B => n49, Z => SUM_11_port);
   U22 : XOR2_X1 port map( A => A(10), B => n50, Z => SUM_10_port);
   U23 : XOR2_X1 port map( A => A(8), B => n52, Z => SUM_8_port);
   U24 : XOR2_X1 port map( A => A(7), B => n53, Z => SUM_7_port);
   U25 : XOR2_X1 port map( A => A(6), B => n54, Z => SUM_6_port);
   U26 : XOR2_X1 port map( A => A(5), B => n55, Z => SUM_5_port);
   U27 : XOR2_X1 port map( A => A(4), B => n56, Z => SUM_4_port);
   U28 : XOR2_X1 port map( A => A(31), B => n57, Z => SUM_31_port);
   U29 : XOR2_X1 port map( A => A(9), B => n51, Z => SUM_9_port);
   U30 : AND2_X1 port map( A1 => A(29), A2 => n31, ZN => n30);
   U31 : AND2_X1 port map( A1 => A(28), A2 => n32, ZN => n31);
   U32 : AND2_X1 port map( A1 => A(27), A2 => n33, ZN => n32);
   U33 : AND2_X1 port map( A1 => A(26), A2 => n34, ZN => n33);
   U34 : AND2_X1 port map( A1 => A(25), A2 => n35, ZN => n34);
   U35 : AND2_X1 port map( A1 => A(24), A2 => n36, ZN => n35);
   U36 : AND2_X1 port map( A1 => A(23), A2 => n37, ZN => n36);
   U37 : AND2_X1 port map( A1 => A(22), A2 => n38, ZN => n37);
   U38 : AND2_X1 port map( A1 => A(21), A2 => n39, ZN => n38);
   U39 : AND2_X1 port map( A1 => A(20), A2 => n40, ZN => n39);
   U40 : AND2_X1 port map( A1 => A(19), A2 => n41, ZN => n40);
   U41 : AND2_X1 port map( A1 => A(18), A2 => n42, ZN => n41);
   U42 : AND2_X1 port map( A1 => A(17), A2 => n43, ZN => n42);
   U43 : AND2_X1 port map( A1 => A(16), A2 => n44, ZN => n43);
   U44 : AND2_X1 port map( A1 => A(15), A2 => n45, ZN => n44);
   U45 : AND2_X1 port map( A1 => A(14), A2 => n46, ZN => n45);
   U46 : AND2_X1 port map( A1 => A(13), A2 => n47, ZN => n46);
   U47 : AND2_X1 port map( A1 => A(12), A2 => n48, ZN => n47);
   U48 : AND2_X1 port map( A1 => A(11), A2 => n49, ZN => n48);
   U49 : AND2_X1 port map( A1 => A(10), A2 => n50, ZN => n49);
   U50 : AND2_X1 port map( A1 => A(9), A2 => n51, ZN => n50);
   U51 : AND2_X1 port map( A1 => A(8), A2 => n52, ZN => n51);
   U52 : AND2_X1 port map( A1 => A(7), A2 => n53, ZN => n52);
   U53 : AND2_X1 port map( A1 => A(6), A2 => n54, ZN => n53);
   U54 : AND2_X1 port map( A1 => A(5), A2 => n55, ZN => n54);
   U55 : AND2_X1 port map( A1 => A(4), A2 => n56, ZN => n55);
   U56 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n56);
   U57 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U58 : AND2_X1 port map( A1 => A(30), A2 => n30, ZN => n57);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_6;

architecture SYN_BEHAVIORAL of MUX21_N4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => S, B2 => B(3), ZN => n13
                           );
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => S, ZN => n11
                           );
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => S, ZN => n12
                           );
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => S, ZN => n10
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_5;

architecture SYN_BEHAVIORAL of MUX21_N4_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => S, B2 => B(3), ZN => n13
                           );
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => S, ZN => n10
                           );
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => S, ZN => n11
                           );
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => S, ZN => n12
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_4;

architecture SYN_BEHAVIORAL of MUX21_N4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => S, B2 => B(3), ZN => n13
                           );
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => S, ZN => n10
                           );
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => S, ZN => n11
                           );
   U8 : INV_X1 port map( A => n12, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => S, ZN => n12
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_3;

architecture SYN_BEHAVIORAL of MUX21_N4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => S, B2 => B(3), ZN => n13
                           );
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => S, ZN => n11
                           );
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => S, ZN => n12
                           );
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => S, ZN => n10
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_2;

architecture SYN_BEHAVIORAL of MUX21_N4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => S, B2 => B(3), ZN => n13
                           );
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => S, ZN => n11
                           );
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => S, ZN => n12
                           );
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => S, ZN => n10
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_1;

architecture SYN_BEHAVIORAL of MUX21_N4_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => S, B2 => B(3), ZN => n13
                           );
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => S, ZN => n11
                           );
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => S, ZN => n12
                           );
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => S, ZN => n10
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_0;

architecture SYN_BEHAVIORAL of MUX21_N4_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => S, B2 => B(3), ZN => n13
                           );
   U4 : INV_X1 port map( A => n11, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => S, ZN => n11
                           );
   U6 : INV_X1 port map( A => n12, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => S, ZN => n12
                           );
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => S, ZN => n10
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_BEHAVIORAL of RCA_N4_14 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27, n28, n29 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => n2, B => n5, Z => n28);
   U16 : XOR2_X1 port map( A => n18, B => n27, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n27);
   U18 : XOR2_X1 port map( A => n26, B => n25, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n25);
   U20 : XOR2_X1 port map( A => A(0), B => n24, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n24);
   U1 : INV_X1 port map( A => B(0), ZN => n1);
   U2 : INV_X1 port map( A => A(0), ZN => n4);
   U3 : INV_X1 port map( A => n5, ZN => n17);
   U4 : INV_X1 port map( A => n2, ZN => n3);
   U5 : OAI22_X1 port map( A1 => n29, A2 => n17, B1 => n23, B2 => n3, ZN => Co)
                           ;
   U6 : AND2_X1 port map( A1 => n17, A2 => n29, ZN => n23);
   U7 : BUF_X1 port map( A => A(3), Z => n5);
   U8 : BUF_X1 port map( A => B(3), Z => n2);
   U9 : AOI22_X1 port map( A1 => n18, A2 => A(2), B1 => n22, B2 => B(2), ZN => 
                           n29);
   U10 : OR2_X1 port map( A1 => A(2), A2 => n18, ZN => n22);
   U11 : INV_X1 port map( A => n21, ZN => n18);
   U12 : AOI22_X1 port map( A1 => n26, A2 => A(1), B1 => n20, B2 => B(1), ZN =>
                           n21);
   U13 : OR2_X1 port map( A1 => A(1), A2 => n26, ZN => n20);
   U14 : OAI21_X1 port map( B1 => n4, B2 => n1, A => n19, ZN => n26);
   U22 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n19);
   U23 : XNOR2_X1 port map( A => n29, B => n28, ZN => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_BEHAVIORAL of RCA_N4_13 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27, n28 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => n3, Z => n27);
   U16 : XOR2_X1 port map( A => n5, B => n26, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n26);
   U18 : XOR2_X1 port map( A => n25, B => n24, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n24);
   U20 : XOR2_X1 port map( A => A(0), B => n23, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n23);
   U1 : INV_X1 port map( A => n3, ZN => n4);
   U2 : BUF_X1 port map( A => A(3), Z => n3);
   U3 : INV_X1 port map( A => B(0), ZN => n1);
   U4 : INV_X1 port map( A => A(0), ZN => n2);
   U5 : OAI22_X1 port map( A1 => n28, A2 => n4, B1 => n22, B2 => n17, ZN => Co)
                           ;
   U6 : AND2_X1 port map( A1 => n4, A2 => n28, ZN => n22);
   U7 : XNOR2_X1 port map( A => n28, B => n27, ZN => S(3));
   U8 : AOI22_X1 port map( A1 => n5, A2 => A(2), B1 => n21, B2 => B(2), ZN => 
                           n28);
   U9 : OR2_X1 port map( A1 => A(2), A2 => n5, ZN => n21);
   U10 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n18, ZN => n25);
   U11 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n18);
   U12 : INV_X1 port map( A => B(3), ZN => n17);
   U13 : INV_X1 port map( A => n20, ZN => n5);
   U14 : AOI22_X1 port map( A1 => n25, A2 => A(1), B1 => n19, B2 => B(1), ZN =>
                           n20);
   U22 : OR2_X1 port map( A1 => A(1), A2 => n25, ZN => n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_BEHAVIORAL of RCA_N4_12 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27, n28 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => n3, Z => n27);
   U16 : XOR2_X1 port map( A => n5, B => n26, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n26);
   U18 : XOR2_X1 port map( A => n25, B => n24, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n24);
   U20 : XOR2_X1 port map( A => A(0), B => n23, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n23);
   U1 : INV_X1 port map( A => n3, ZN => n4);
   U2 : BUF_X1 port map( A => A(3), Z => n3);
   U3 : INV_X1 port map( A => B(0), ZN => n1);
   U4 : INV_X1 port map( A => A(0), ZN => n2);
   U5 : OAI22_X1 port map( A1 => n28, A2 => n4, B1 => n22, B2 => n17, ZN => Co)
                           ;
   U6 : AND2_X1 port map( A1 => n4, A2 => n28, ZN => n22);
   U7 : XNOR2_X1 port map( A => n28, B => n27, ZN => S(3));
   U8 : AOI22_X1 port map( A1 => n5, A2 => A(2), B1 => n21, B2 => B(2), ZN => 
                           n28);
   U9 : OR2_X1 port map( A1 => A(2), A2 => n5, ZN => n21);
   U10 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n18, ZN => n25);
   U11 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n18);
   U12 : INV_X1 port map( A => B(3), ZN => n17);
   U13 : INV_X1 port map( A => n20, ZN => n5);
   U14 : AOI22_X1 port map( A1 => n25, A2 => A(1), B1 => n19, B2 => B(1), ZN =>
                           n20);
   U22 : OR2_X1 port map( A1 => A(1), A2 => n25, ZN => n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_BEHAVIORAL of RCA_N4_11 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27, n28 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => n2, Z => n27);
   U16 : XOR2_X1 port map( A => n4, B => n26, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n26);
   U18 : XOR2_X1 port map( A => n25, B => n24, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n24);
   U20 : XOR2_X1 port map( A => A(0), B => n23, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n23);
   U1 : INV_X1 port map( A => n2, ZN => n3);
   U2 : BUF_X1 port map( A => A(3), Z => n2);
   U3 : INV_X1 port map( A => A(0), ZN => n1);
   U4 : OAI22_X1 port map( A1 => n28, A2 => n3, B1 => n22, B2 => n5, ZN => Co);
   U5 : XNOR2_X1 port map( A => n28, B => n27, ZN => S(3));
   U6 : AND2_X1 port map( A1 => n3, A2 => n28, ZN => n22);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A(2), B1 => n21, B2 => B(2), ZN => 
                           n28);
   U8 : OR2_X1 port map( A1 => A(2), A2 => n4, ZN => n21);
   U9 : OAI21_X1 port map( B1 => n1, B2 => n17, A => n18, ZN => n25);
   U10 : INV_X1 port map( A => B(0), ZN => n17);
   U11 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n18);
   U12 : INV_X1 port map( A => B(3), ZN => n5);
   U13 : INV_X1 port map( A => n20, ZN => n4);
   U14 : AOI22_X1 port map( A1 => n25, A2 => A(1), B1 => n19, B2 => B(1), ZN =>
                           n20);
   U22 : OR2_X1 port map( A1 => A(1), A2 => n25, ZN => n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_BEHAVIORAL of RCA_N4_10 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27, n28 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => n2, Z => n27);
   U16 : XOR2_X1 port map( A => n4, B => n26, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n26);
   U18 : XOR2_X1 port map( A => n25, B => n24, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n24);
   U20 : XOR2_X1 port map( A => A(0), B => n23, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n23);
   U1 : INV_X1 port map( A => n2, ZN => n3);
   U2 : BUF_X1 port map( A => A(3), Z => n2);
   U3 : INV_X1 port map( A => A(0), ZN => n1);
   U4 : OAI22_X1 port map( A1 => n28, A2 => n3, B1 => n22, B2 => n5, ZN => Co);
   U5 : XNOR2_X1 port map( A => n28, B => n27, ZN => S(3));
   U6 : AND2_X1 port map( A1 => n3, A2 => n28, ZN => n22);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A(2), B1 => n21, B2 => B(2), ZN => 
                           n28);
   U8 : OR2_X1 port map( A1 => A(2), A2 => n4, ZN => n21);
   U9 : OAI21_X1 port map( B1 => n1, B2 => n17, A => n18, ZN => n25);
   U10 : INV_X1 port map( A => B(0), ZN => n17);
   U11 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n18);
   U12 : INV_X1 port map( A => B(3), ZN => n5);
   U13 : INV_X1 port map( A => n20, ZN => n4);
   U14 : AOI22_X1 port map( A1 => n25, A2 => A(1), B1 => n19, B2 => B(1), ZN =>
                           n20);
   U22 : OR2_X1 port map( A1 => A(1), A2 => n25, ZN => n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_BEHAVIORAL of RCA_N4_9 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27, n28 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => n2, Z => n27);
   U16 : XOR2_X1 port map( A => n4, B => n26, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n26);
   U18 : XOR2_X1 port map( A => n25, B => n24, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n24);
   U20 : XOR2_X1 port map( A => A(0), B => n23, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n23);
   U1 : INV_X1 port map( A => n2, ZN => n3);
   U2 : BUF_X1 port map( A => A(3), Z => n2);
   U3 : INV_X1 port map( A => A(0), ZN => n1);
   U4 : OAI22_X1 port map( A1 => n28, A2 => n3, B1 => n22, B2 => n5, ZN => Co);
   U5 : XNOR2_X1 port map( A => n28, B => n27, ZN => S(3));
   U6 : AND2_X1 port map( A1 => n3, A2 => n28, ZN => n22);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A(2), B1 => n21, B2 => B(2), ZN => 
                           n28);
   U8 : OR2_X1 port map( A1 => A(2), A2 => n4, ZN => n21);
   U9 : OAI21_X1 port map( B1 => n1, B2 => n17, A => n18, ZN => n25);
   U10 : INV_X1 port map( A => B(0), ZN => n17);
   U11 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n18);
   U12 : INV_X1 port map( A => B(3), ZN => n5);
   U13 : INV_X1 port map( A => n20, ZN => n4);
   U14 : AOI22_X1 port map( A1 => n25, A2 => A(1), B1 => n19, B2 => B(1), ZN =>
                           n20);
   U22 : OR2_X1 port map( A1 => A(1), A2 => n25, ZN => n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_BEHAVIORAL of RCA_N4_8 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27, n28 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => n2, Z => n27);
   U16 : XOR2_X1 port map( A => n4, B => n26, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n26);
   U18 : XOR2_X1 port map( A => n25, B => n24, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n24);
   U20 : XOR2_X1 port map( A => A(0), B => n23, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n23);
   U1 : INV_X1 port map( A => n2, ZN => n3);
   U2 : BUF_X1 port map( A => A(3), Z => n2);
   U3 : INV_X1 port map( A => A(0), ZN => n1);
   U4 : OAI22_X1 port map( A1 => n28, A2 => n3, B1 => n22, B2 => n5, ZN => Co);
   U5 : XNOR2_X1 port map( A => n28, B => n27, ZN => S(3));
   U6 : AND2_X1 port map( A1 => n3, A2 => n28, ZN => n22);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A(2), B1 => n21, B2 => B(2), ZN => 
                           n28);
   U8 : OR2_X1 port map( A1 => A(2), A2 => n4, ZN => n21);
   U9 : OAI21_X1 port map( B1 => n1, B2 => n17, A => n18, ZN => n25);
   U10 : INV_X1 port map( A => B(0), ZN => n17);
   U11 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n18);
   U12 : INV_X1 port map( A => B(3), ZN => n5);
   U13 : INV_X1 port map( A => n20, ZN => n4);
   U14 : AOI22_X1 port map( A1 => n25, A2 => A(1), B1 => n19, B2 => B(1), ZN =>
                           n20);
   U22 : OR2_X1 port map( A1 => A(1), A2 => n25, ZN => n19);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_BEHAVIORAL of RCA_N4_7 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => A(3), Z => n26);
   U16 : XOR2_X1 port map( A => n1, B => n25, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n25);
   U18 : XOR2_X1 port map( A => n24, B => n23, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n23);
   U20 : XOR2_X1 port map( A => A(0), B => n22, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n22);
   U1 : OAI22_X1 port map( A1 => n27, A2 => n2, B1 => n21, B2 => n4, ZN => Co);
   U2 : AND2_X1 port map( A1 => n2, A2 => n27, ZN => n21);
   U3 : XNOR2_X1 port map( A => n27, B => n26, ZN => S(3));
   U4 : AOI22_X1 port map( A1 => n1, A2 => A(2), B1 => n20, B2 => B(2), ZN => 
                           n27);
   U5 : OR2_X1 port map( A1 => A(2), A2 => n1, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n5, A => n17, ZN => n24);
   U7 : INV_X1 port map( A => B(0), ZN => n5);
   U8 : INV_X1 port map( A => A(0), ZN => n3);
   U9 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U10 : INV_X1 port map( A => A(3), ZN => n2);
   U11 : INV_X1 port map( A => B(3), ZN => n4);
   U12 : INV_X1 port map( A => n19, ZN => n1);
   U13 : AOI22_X1 port map( A1 => n24, A2 => A(1), B1 => n18, B2 => B(1), ZN =>
                           n19);
   U14 : OR2_X1 port map( A1 => A(1), A2 => n24, ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_BEHAVIORAL of RCA_N4_6 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => A(3), Z => n26);
   U16 : XOR2_X1 port map( A => n1, B => n25, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n25);
   U18 : XOR2_X1 port map( A => n24, B => n23, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n23);
   U20 : XOR2_X1 port map( A => A(0), B => n22, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n22);
   U1 : OAI22_X1 port map( A1 => n27, A2 => n2, B1 => n21, B2 => n4, ZN => Co);
   U2 : AND2_X1 port map( A1 => n2, A2 => n27, ZN => n21);
   U3 : XNOR2_X1 port map( A => n27, B => n26, ZN => S(3));
   U4 : AOI22_X1 port map( A1 => n1, A2 => A(2), B1 => n20, B2 => B(2), ZN => 
                           n27);
   U5 : OR2_X1 port map( A1 => A(2), A2 => n1, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n5, A => n17, ZN => n24);
   U7 : INV_X1 port map( A => B(0), ZN => n5);
   U8 : INV_X1 port map( A => A(0), ZN => n3);
   U9 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U10 : INV_X1 port map( A => A(3), ZN => n2);
   U11 : INV_X1 port map( A => B(3), ZN => n4);
   U12 : INV_X1 port map( A => n19, ZN => n1);
   U13 : AOI22_X1 port map( A1 => n24, A2 => A(1), B1 => n18, B2 => B(1), ZN =>
                           n19);
   U14 : OR2_X1 port map( A1 => A(1), A2 => n24, ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_BEHAVIORAL of RCA_N4_5 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => A(3), Z => n26);
   U16 : XOR2_X1 port map( A => n1, B => n25, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n25);
   U18 : XOR2_X1 port map( A => n24, B => n23, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n23);
   U20 : XOR2_X1 port map( A => A(0), B => n22, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n22);
   U1 : OAI22_X1 port map( A1 => n27, A2 => n2, B1 => n21, B2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => n27, B => n26, ZN => S(3));
   U3 : AND2_X1 port map( A1 => n2, A2 => n27, ZN => n21);
   U4 : AOI22_X1 port map( A1 => n1, A2 => A(2), B1 => n20, B2 => B(2), ZN => 
                           n27);
   U5 : OR2_X1 port map( A1 => A(2), A2 => n1, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n5, A => n17, ZN => n24);
   U7 : INV_X1 port map( A => B(0), ZN => n5);
   U8 : INV_X1 port map( A => A(0), ZN => n3);
   U9 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U10 : INV_X1 port map( A => A(3), ZN => n2);
   U11 : INV_X1 port map( A => B(3), ZN => n4);
   U12 : INV_X1 port map( A => n19, ZN => n1);
   U13 : AOI22_X1 port map( A1 => n24, A2 => A(1), B1 => n18, B2 => B(1), ZN =>
                           n19);
   U14 : OR2_X1 port map( A1 => A(1), A2 => n24, ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_BEHAVIORAL of RCA_N4_4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => A(3), Z => n26);
   U16 : XOR2_X1 port map( A => n1, B => n25, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n25);
   U18 : XOR2_X1 port map( A => n24, B => n23, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n23);
   U20 : XOR2_X1 port map( A => A(0), B => n22, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n22);
   U1 : OAI22_X1 port map( A1 => n27, A2 => n2, B1 => n21, B2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => n27, B => n26, ZN => S(3));
   U3 : AND2_X1 port map( A1 => n2, A2 => n27, ZN => n21);
   U4 : AOI22_X1 port map( A1 => n1, A2 => A(2), B1 => n20, B2 => B(2), ZN => 
                           n27);
   U5 : OR2_X1 port map( A1 => A(2), A2 => n1, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n5, A => n17, ZN => n24);
   U7 : INV_X1 port map( A => B(0), ZN => n5);
   U8 : INV_X1 port map( A => A(0), ZN => n3);
   U9 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U10 : INV_X1 port map( A => A(3), ZN => n2);
   U11 : INV_X1 port map( A => B(3), ZN => n4);
   U12 : INV_X1 port map( A => n19, ZN => n1);
   U13 : AOI22_X1 port map( A1 => n24, A2 => A(1), B1 => n18, B2 => B(1), ZN =>
                           n19);
   U14 : OR2_X1 port map( A1 => A(1), A2 => n24, ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_BEHAVIORAL of RCA_N4_3 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => A(3), Z => n26);
   U16 : XOR2_X1 port map( A => n1, B => n25, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n25);
   U18 : XOR2_X1 port map( A => n24, B => n23, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n23);
   U20 : XOR2_X1 port map( A => A(0), B => n22, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n22);
   U1 : OAI22_X1 port map( A1 => n27, A2 => n2, B1 => n21, B2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => n27, B => n26, ZN => S(3));
   U3 : AND2_X1 port map( A1 => n2, A2 => n27, ZN => n21);
   U4 : AOI22_X1 port map( A1 => n1, A2 => A(2), B1 => n20, B2 => B(2), ZN => 
                           n27);
   U5 : OR2_X1 port map( A1 => A(2), A2 => n1, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n5, A => n17, ZN => n24);
   U7 : INV_X1 port map( A => B(0), ZN => n5);
   U8 : INV_X1 port map( A => A(0), ZN => n3);
   U9 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U10 : INV_X1 port map( A => A(3), ZN => n2);
   U11 : INV_X1 port map( A => B(3), ZN => n4);
   U12 : INV_X1 port map( A => n19, ZN => n1);
   U13 : AOI22_X1 port map( A1 => n24, A2 => A(1), B1 => n18, B2 => B(1), ZN =>
                           n19);
   U14 : OR2_X1 port map( A1 => A(1), A2 => n24, ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_BEHAVIORAL of RCA_N4_2 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => A(3), Z => n26);
   U16 : XOR2_X1 port map( A => n1, B => n25, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n25);
   U18 : XOR2_X1 port map( A => n24, B => n23, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n23);
   U20 : XOR2_X1 port map( A => A(0), B => n22, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n22);
   U1 : OAI22_X1 port map( A1 => n27, A2 => n2, B1 => n21, B2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => n27, B => n26, ZN => S(3));
   U3 : AND2_X1 port map( A1 => n2, A2 => n27, ZN => n21);
   U4 : AOI22_X1 port map( A1 => n1, A2 => A(2), B1 => n20, B2 => B(2), ZN => 
                           n27);
   U5 : OR2_X1 port map( A1 => A(2), A2 => n1, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n5, A => n17, ZN => n24);
   U7 : INV_X1 port map( A => B(0), ZN => n5);
   U8 : INV_X1 port map( A => A(0), ZN => n3);
   U9 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U10 : INV_X1 port map( A => A(3), ZN => n2);
   U11 : INV_X1 port map( A => B(3), ZN => n4);
   U12 : INV_X1 port map( A => n19, ZN => n1);
   U13 : AOI22_X1 port map( A1 => n24, A2 => A(1), B1 => n18, B2 => B(1), ZN =>
                           n19);
   U14 : OR2_X1 port map( A1 => A(1), A2 => n24, ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_BEHAVIORAL of RCA_N4_1 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => A(3), Z => n26);
   U16 : XOR2_X1 port map( A => n1, B => n25, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n25);
   U18 : XOR2_X1 port map( A => n24, B => n23, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n23);
   U20 : XOR2_X1 port map( A => A(0), B => n22, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n22);
   U1 : OAI22_X1 port map( A1 => n27, A2 => n2, B1 => n21, B2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => n27, B => n26, ZN => S(3));
   U3 : AND2_X1 port map( A1 => n2, A2 => n27, ZN => n21);
   U4 : AOI22_X1 port map( A1 => n1, A2 => A(2), B1 => n20, B2 => B(2), ZN => 
                           n27);
   U5 : OR2_X1 port map( A1 => A(2), A2 => n1, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n5, A => n17, ZN => n24);
   U7 : INV_X1 port map( A => B(0), ZN => n5);
   U8 : INV_X1 port map( A => A(0), ZN => n3);
   U9 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U10 : INV_X1 port map( A => A(3), ZN => n2);
   U11 : INV_X1 port map( A => B(3), ZN => n4);
   U12 : INV_X1 port map( A => n19, ZN => n1);
   U13 : AOI22_X1 port map( A1 => n24, A2 => A(1), B1 => n18, B2 => B(1), ZN =>
                           n19);
   U14 : OR2_X1 port map( A1 => A(1), A2 => n24, ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_BEHAVIORAL of RCA_N4_0 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => B(3), B => A(3), Z => n26);
   U16 : XOR2_X1 port map( A => n1, B => n25, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n25);
   U18 : XOR2_X1 port map( A => n24, B => n23, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n23);
   U20 : XOR2_X1 port map( A => A(0), B => n22, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n22);
   U1 : OAI22_X1 port map( A1 => n27, A2 => n2, B1 => n21, B2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => n27, B => n26, ZN => S(3));
   U3 : AND2_X1 port map( A1 => n2, A2 => n27, ZN => n21);
   U4 : AOI22_X1 port map( A1 => n1, A2 => A(2), B1 => n20, B2 => B(2), ZN => 
                           n27);
   U5 : OR2_X1 port map( A1 => A(2), A2 => n1, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n5, A => n17, ZN => n24);
   U7 : INV_X1 port map( A => B(0), ZN => n5);
   U8 : INV_X1 port map( A => A(0), ZN => n3);
   U9 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U10 : INV_X1 port map( A => A(3), ZN => n2);
   U11 : INV_X1 port map( A => B(3), ZN => n4);
   U12 : INV_X1 port map( A => n19, ZN => n1);
   U13 : AOI22_X1 port map( A1 => n24, A2 => A(1), B1 => n18, B2 => B(1), ZN =>
                           n19);
   U14 : OR2_X1 port map( A1 => A(1), A2 => n24, ZN => n18);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_6 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_6;

architecture SYN_BEHAVIORAL of ENCODER_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8, n9 : std_logic;

begin
   
   U10 : XOR2_X1 port map( A => B(0), B => B(1), Z => n8);
   U3 : NOR3_X1 port map( A1 => n2, A2 => n9, A3 => n8, ZN => Y(2));
   U4 : OAI21_X1 port map( B1 => n6, B2 => n2, A => n7, ZN => Y(1));
   U5 : OAI21_X1 port map( B1 => n1, B2 => n6, A => n7, ZN => Y(0));
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n9, A2 => n2, ZN => n7);
   U8 : INV_X1 port map( A => n1, ZN => n2);
   U9 : AND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n9);
   U11 : BUF_X1 port map( A => B(2), Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_5 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_5;

architecture SYN_BEHAVIORAL of ENCODER_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U10 : XOR2_X1 port map( A => B(0), B => B(1), Z => n7);
   U3 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => Y(2));
   U4 : INV_X1 port map( A => n7, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => Y(1));
   U6 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U7 : AND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n8);
   U8 : OAI21_X1 port map( B1 => B(2), B2 => n2, A => n6, ZN => Y(0));
   U9 : INV_X1 port map( A => B(2), ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_4 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_4;

architecture SYN_BEHAVIORAL of ENCODER_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U10 : XOR2_X1 port map( A => B(0), B => B(1), Z => n7);
   U3 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => Y(2));
   U4 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => Y(1));
   U5 : INV_X1 port map( A => n7, ZN => n2);
   U6 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U7 : OAI21_X1 port map( B1 => B(2), B2 => n2, A => n6, ZN => Y(0));
   U8 : INV_X1 port map( A => B(2), ZN => n1);
   U9 : AND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_3 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_3;

architecture SYN_BEHAVIORAL of ENCODER_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U10 : XOR2_X1 port map( A => B(0), B => B(1), Z => n7);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => n2, A => n6, ZN => Y(0));
   U4 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => Y(2));
   U5 : INV_X1 port map( A => n7, ZN => n2);
   U6 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U7 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => Y(1));
   U8 : INV_X1 port map( A => B(2), ZN => n1);
   U9 : AND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_2 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_2;

architecture SYN_BEHAVIORAL of ENCODER_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U10 : XOR2_X1 port map( A => B(0), B => B(1), Z => n7);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => n2, A => n6, ZN => Y(0));
   U4 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => Y(2));
   U5 : INV_X1 port map( A => n7, ZN => n2);
   U6 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U7 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => Y(1));
   U8 : INV_X1 port map( A => B(2), ZN => n1);
   U9 : AND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_1 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_1;

architecture SYN_BEHAVIORAL of ENCODER_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U10 : XOR2_X1 port map( A => B(0), B => B(1), Z => n7);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => n2, A => n6, ZN => Y(0));
   U4 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => Y(2));
   U5 : INV_X1 port map( A => n7, ZN => n2);
   U6 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U7 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => Y(1));
   U8 : INV_X1 port map( A => B(2), ZN => n1);
   U9 : AND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_0 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_0;

architecture SYN_BEHAVIORAL of ENCODER_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n6, n7, n8 : std_logic;

begin
   
   U10 : XOR2_X1 port map( A => B(0), B => B(1), Z => n7);
   U3 : OAI21_X1 port map( B1 => B(2), B2 => n2, A => n6, ZN => Y(0));
   U4 : NOR3_X1 port map( A1 => n1, A2 => n8, A3 => n7, ZN => Y(2));
   U5 : INV_X1 port map( A => n7, ZN => n2);
   U6 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => n6);
   U7 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n6, ZN => Y(1));
   U8 : INV_X1 port map( A => B(2), ZN => n1);
   U9 : AND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_5;

architecture SYN_STRUCTURAL of CSB_N4_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n1, n2, 
      n_1203, n_1204 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_11 port map( A(3) => n2, A(2) => A(2), A(1) => A(1), A(0) => 
                           n1, B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0) 
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1203);
   RCA1 : RCA_N4_10 port map( A(3) => n2, A(2) => A(2), A(1) => A(1), A(0) => 
                           n1, B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0) 
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1204);
   MUX : MUX21_N4_5 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : BUF_X1 port map( A => A(0), Z => n1);
   U4 : BUF_X1 port map( A => A(3), Z => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_4;

architecture SYN_STRUCTURAL of CSB_N4_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n1, n2, 
      n_1205, n_1206 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_9 port map( A(3) => n2, A(2) => A(2), A(1) => A(1), A(0) => n1
                           , B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0) => 
                           B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, S(2)
                           => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1205);
   RCA1 : RCA_N4_8 port map( A(3) => n2, A(2) => A(2), A(1) => A(1), A(0) => n1
                           , B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0) => 
                           B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, S(2)
                           => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1206);
   MUX : MUX21_N4_4 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : BUF_X1 port map( A => A(0), Z => n1);
   U4 : BUF_X1 port map( A => A(3), Z => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_3;

architecture SYN_STRUCTURAL of CSB_N4_3 is

   component MUX21_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1207, 
      n_1208 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1207);
   RCA1 : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1208);
   MUX : MUX21_N4_3 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_2;

architecture SYN_STRUCTURAL of CSB_N4_2 is

   component MUX21_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1209, 
      n_1210 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1209);
   RCA1 : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1210);
   MUX : MUX21_N4_2 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_1;

architecture SYN_STRUCTURAL of CSB_N4_1 is

   component MUX21_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1211, 
      n_1212 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1211);
   RCA1 : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1212);
   MUX : MUX21_N4_1 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_0;

architecture SYN_STRUCTURAL of CSB_N4_0 is

   component MUX21_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1213, 
      n_1214 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1213);
   RCA1 : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1214);
   MUX : MUX21_N4_0 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_32 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_32;

architecture SYN_BEHAVIORAL of PG_BLOCK_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_31 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_31;

architecture SYN_BEHAVIORAL of PG_BLOCK_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_30 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_30;

architecture SYN_BEHAVIORAL of PG_BLOCK_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_29 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_29;

architecture SYN_BEHAVIORAL of PG_BLOCK_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_28 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_28;

architecture SYN_BEHAVIORAL of PG_BLOCK_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_27 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_27;

architecture SYN_BEHAVIORAL of PG_BLOCK_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_26 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_26;

architecture SYN_BEHAVIORAL of PG_BLOCK_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_25 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_25;

architecture SYN_BEHAVIORAL of PG_BLOCK_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_24 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_24;

architecture SYN_BEHAVIORAL of PG_BLOCK_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_23 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_23;

architecture SYN_BEHAVIORAL of PG_BLOCK_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_22 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_22;

architecture SYN_BEHAVIORAL of PG_BLOCK_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_21 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_21;

architecture SYN_BEHAVIORAL of PG_BLOCK_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_20 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_20;

architecture SYN_BEHAVIORAL of PG_BLOCK_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_19 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_19;

architecture SYN_BEHAVIORAL of PG_BLOCK_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_18 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_18;

architecture SYN_BEHAVIORAL of PG_BLOCK_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_17 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_17;

architecture SYN_BEHAVIORAL of PG_BLOCK_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_16 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_16;

architecture SYN_BEHAVIORAL of PG_BLOCK_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_15 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_15;

architecture SYN_BEHAVIORAL of PG_BLOCK_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_14 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_14;

architecture SYN_BEHAVIORAL of PG_BLOCK_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_13 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_13;

architecture SYN_BEHAVIORAL of PG_BLOCK_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_12 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_12;

architecture SYN_BEHAVIORAL of PG_BLOCK_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_11 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_11;

architecture SYN_BEHAVIORAL of PG_BLOCK_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_10 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_10;

architecture SYN_BEHAVIORAL of PG_BLOCK_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_9 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_9;

architecture SYN_BEHAVIORAL of PG_BLOCK_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_8 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_8;

architecture SYN_BEHAVIORAL of PG_BLOCK_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_7 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_7;

architecture SYN_BEHAVIORAL of PG_BLOCK_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_6 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_6;

architecture SYN_BEHAVIORAL of PG_BLOCK_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_5 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_5;

architecture SYN_BEHAVIORAL of PG_BLOCK_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_4 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_4;

architecture SYN_BEHAVIORAL of PG_BLOCK_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_3 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_3;

architecture SYN_BEHAVIORAL of PG_BLOCK_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_2 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_2;

architecture SYN_BEHAVIORAL of PG_BLOCK_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_1 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_1;

architecture SYN_BEHAVIORAL of PG_BLOCK_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_0 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_0;

architecture SYN_BEHAVIORAL of PG_BLOCK_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_7 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_7;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_6 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_6;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_5 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_5;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_4 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_4;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_3 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_3;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_2 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_2;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_1 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_1;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_0 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_0;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_N32_1;

architecture SYN_BEHAVIORAL of RCA_N32_1 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237 : std_logic;

begin
   
   U129 : XOR2_X1 port map( A => n237, B => n236, Z => S(9));
   U130 : XOR2_X1 port map( A => B(9), B => A(9), Z => n236);
   U131 : XOR2_X1 port map( A => B(8), B => A(8), Z => n234);
   U132 : XOR2_X1 port map( A => n233, B => n232, Z => S(7));
   U133 : XOR2_X1 port map( A => B(7), B => A(7), Z => n232);
   U134 : XOR2_X1 port map( A => B(6), B => A(6), Z => n230);
   U135 : XOR2_X1 port map( A => n229, B => n228, Z => S(5));
   U136 : XOR2_X1 port map( A => B(5), B => A(5), Z => n228);
   U137 : XOR2_X1 port map( A => B(4), B => A(4), Z => n226);
   U138 : XOR2_X1 port map( A => B(3), B => A(3), Z => n224);
   U139 : XOR2_X1 port map( A => n1, B => n223, Z => S(31));
   U140 : XOR2_X1 port map( A => B(31), B => A(31), Z => n223);
   U141 : XOR2_X1 port map( A => n222, B => n221, Z => S(30));
   U142 : XOR2_X1 port map( A => B(30), B => A(30), Z => n221);
   U143 : XOR2_X1 port map( A => B(2), B => A(2), Z => n219);
   U144 : XOR2_X1 port map( A => B(28), B => A(28), Z => n216);
   U145 : XOR2_X1 port map( A => n215, B => n214, Z => S(27));
   U146 : XOR2_X1 port map( A => B(27), B => A(27), Z => n214);
   U147 : XOR2_X1 port map( A => B(26), B => A(26), Z => n212);
   U148 : XOR2_X1 port map( A => n211, B => n210, Z => S(25));
   U149 : XOR2_X1 port map( A => B(25), B => A(25), Z => n210);
   U150 : XOR2_X1 port map( A => B(24), B => A(24), Z => n208);
   U151 : XOR2_X1 port map( A => n207, B => n206, Z => S(23));
   U152 : XOR2_X1 port map( A => B(23), B => A(23), Z => n206);
   U153 : XOR2_X1 port map( A => B(22), B => A(22), Z => n204);
   U154 : XOR2_X1 port map( A => n203, B => n202, Z => S(21));
   U155 : XOR2_X1 port map( A => B(21), B => A(21), Z => n202);
   U156 : XOR2_X1 port map( A => B(20), B => A(20), Z => n200);
   U157 : XOR2_X1 port map( A => B(1), B => A(1), Z => n198);
   U158 : XOR2_X1 port map( A => n197, B => n196, Z => S(19));
   U159 : XOR2_X1 port map( A => B(19), B => A(19), Z => n196);
   U160 : XOR2_X1 port map( A => B(18), B => A(18), Z => n194);
   U161 : XOR2_X1 port map( A => n193, B => n192, Z => S(17));
   U162 : XOR2_X1 port map( A => B(17), B => A(17), Z => n192);
   U163 : XOR2_X1 port map( A => B(16), B => A(16), Z => n190);
   U164 : XOR2_X1 port map( A => n189, B => n188, Z => S(15));
   U165 : XOR2_X1 port map( A => B(15), B => A(15), Z => n188);
   U166 : XOR2_X1 port map( A => B(14), B => A(14), Z => n186);
   U167 : XOR2_X1 port map( A => n185, B => n184, Z => S(13));
   U168 : XOR2_X1 port map( A => B(13), B => A(13), Z => n184);
   U169 : XOR2_X1 port map( A => B(12), B => A(12), Z => n182);
   U170 : XOR2_X1 port map( A => n181, B => n180, Z => S(11));
   U171 : XOR2_X1 port map( A => B(11), B => A(11), Z => n180);
   U172 : XOR2_X1 port map( A => n22, B => n179, Z => S(10));
   U173 : XOR2_X1 port map( A => B(10), B => A(10), Z => n179);
   U174 : XOR2_X1 port map( A => A(0), B => n178, Z => S(0));
   U175 : XOR2_X1 port map( A => Ci, B => B(0), Z => n178);
   U1 : XNOR2_X1 port map( A => n3, B => n218, ZN => S(29));
   U2 : XNOR2_X1 port map( A => B(29), B => n31, ZN => n218);
   U3 : INV_X1 port map( A => n173, ZN => n3);
   U4 : OAI21_X1 port map( B1 => n177, B2 => n30, A => n176, ZN => Co);
   U5 : INV_X1 port map( A => n154, ZN => n22);
   U6 : INV_X1 port map( A => n177, ZN => n1);
   U7 : AOI21_X1 port map( B1 => n229, B2 => A(5), A => n27, ZN => n231);
   U8 : INV_X1 port map( A => n148, ZN => n27);
   U9 : OAI21_X1 port map( B1 => A(5), B2 => n229, A => B(5), ZN => n148);
   U10 : AOI21_X1 port map( B1 => n233, B2 => A(7), A => n25, ZN => n235);
   U11 : INV_X1 port map( A => n150, ZN => n25);
   U12 : OAI21_X1 port map( B1 => A(7), B2 => n233, A => B(7), ZN => n150);
   U13 : AOI21_X1 port map( B1 => n181, B2 => A(11), A => n21, ZN => n183);
   U14 : INV_X1 port map( A => n155, ZN => n21);
   U15 : OAI21_X1 port map( B1 => A(11), B2 => n181, A => B(11), ZN => n155);
   U16 : AOI21_X1 port map( B1 => n185, B2 => A(13), A => n19, ZN => n187);
   U17 : INV_X1 port map( A => n157, ZN => n19);
   U18 : OAI21_X1 port map( B1 => A(13), B2 => n185, A => B(13), ZN => n157);
   U19 : AOI21_X1 port map( B1 => n189, B2 => A(15), A => n17, ZN => n191);
   U20 : INV_X1 port map( A => n159, ZN => n17);
   U21 : OAI21_X1 port map( B1 => A(15), B2 => n189, A => B(15), ZN => n159);
   U22 : AOI21_X1 port map( B1 => n193, B2 => A(17), A => n15, ZN => n195);
   U23 : INV_X1 port map( A => n161, ZN => n15);
   U24 : OAI21_X1 port map( B1 => A(17), B2 => n193, A => B(17), ZN => n161);
   U25 : AOI21_X1 port map( B1 => n197, B2 => A(19), A => n13, ZN => n201);
   U26 : INV_X1 port map( A => n163, ZN => n13);
   U27 : OAI21_X1 port map( B1 => A(19), B2 => n197, A => B(19), ZN => n163);
   U28 : AOI21_X1 port map( B1 => n203, B2 => A(21), A => n11, ZN => n205);
   U29 : INV_X1 port map( A => n165, ZN => n11);
   U30 : OAI21_X1 port map( B1 => A(21), B2 => n203, A => B(21), ZN => n165);
   U31 : AOI21_X1 port map( B1 => n207, B2 => A(23), A => n9, ZN => n209);
   U32 : INV_X1 port map( A => n167, ZN => n9);
   U33 : OAI21_X1 port map( B1 => A(23), B2 => n207, A => B(23), ZN => n167);
   U34 : AOI21_X1 port map( B1 => n211, B2 => A(25), A => n7, ZN => n213);
   U35 : INV_X1 port map( A => n169, ZN => n7);
   U36 : OAI21_X1 port map( B1 => A(25), B2 => n211, A => B(25), ZN => n169);
   U37 : AOI21_X1 port map( B1 => n215, B2 => A(27), A => n5, ZN => n217);
   U38 : INV_X1 port map( A => n171, ZN => n5);
   U39 : OAI21_X1 port map( B1 => A(27), B2 => n215, A => B(27), ZN => n171);
   U40 : OAI21_X1 port map( B1 => n235, B2 => n42, A => n151, ZN => n237);
   U41 : INV_X1 port map( A => A(8), ZN => n42);
   U42 : OAI21_X1 port map( B1 => A(8), B2 => n24, A => B(8), ZN => n151);
   U43 : INV_X1 port map( A => n235, ZN => n24);
   U44 : OAI21_X1 port map( B1 => n183, B2 => n40, A => n156, ZN => n185);
   U45 : INV_X1 port map( A => A(12), ZN => n40);
   U46 : OAI21_X1 port map( B1 => A(12), B2 => n20, A => B(12), ZN => n156);
   U47 : INV_X1 port map( A => n183, ZN => n20);
   U48 : OAI21_X1 port map( B1 => n187, B2 => n39, A => n158, ZN => n189);
   U49 : INV_X1 port map( A => A(14), ZN => n39);
   U50 : OAI21_X1 port map( B1 => A(14), B2 => n18, A => B(14), ZN => n158);
   U51 : INV_X1 port map( A => n187, ZN => n18);
   U52 : OAI21_X1 port map( B1 => n191, B2 => n38, A => n160, ZN => n193);
   U53 : INV_X1 port map( A => A(16), ZN => n38);
   U54 : OAI21_X1 port map( B1 => A(16), B2 => n16, A => B(16), ZN => n160);
   U55 : INV_X1 port map( A => n191, ZN => n16);
   U56 : OAI21_X1 port map( B1 => n195, B2 => n37, A => n162, ZN => n197);
   U57 : INV_X1 port map( A => A(18), ZN => n37);
   U58 : OAI21_X1 port map( B1 => A(18), B2 => n14, A => B(18), ZN => n162);
   U59 : INV_X1 port map( A => n195, ZN => n14);
   U60 : OAI21_X1 port map( B1 => n201, B2 => n36, A => n164, ZN => n203);
   U61 : INV_X1 port map( A => A(20), ZN => n36);
   U62 : OAI21_X1 port map( B1 => A(20), B2 => n12, A => B(20), ZN => n164);
   U63 : INV_X1 port map( A => n201, ZN => n12);
   U64 : OAI21_X1 port map( B1 => n205, B2 => n35, A => n166, ZN => n207);
   U65 : INV_X1 port map( A => A(22), ZN => n35);
   U66 : OAI21_X1 port map( B1 => A(22), B2 => n10, A => B(22), ZN => n166);
   U67 : INV_X1 port map( A => n205, ZN => n10);
   U68 : OAI21_X1 port map( B1 => n209, B2 => n34, A => n168, ZN => n211);
   U69 : INV_X1 port map( A => A(24), ZN => n34);
   U70 : OAI21_X1 port map( B1 => A(24), B2 => n8, A => B(24), ZN => n168);
   U71 : INV_X1 port map( A => n209, ZN => n8);
   U72 : OAI21_X1 port map( B1 => n213, B2 => n33, A => n170, ZN => n215);
   U73 : INV_X1 port map( A => A(26), ZN => n33);
   U74 : OAI21_X1 port map( B1 => A(26), B2 => n6, A => B(26), ZN => n170);
   U75 : INV_X1 port map( A => n213, ZN => n6);
   U76 : OAI21_X1 port map( B1 => n231, B2 => n43, A => n149, ZN => n233);
   U77 : INV_X1 port map( A => A(6), ZN => n43);
   U78 : OAI21_X1 port map( B1 => A(6), B2 => n26, A => B(6), ZN => n149);
   U79 : INV_X1 port map( A => n231, ZN => n26);
   U80 : OAI21_X1 port map( B1 => n154, B2 => n41, A => n153, ZN => n181);
   U81 : INV_X1 port map( A => A(10), ZN => n41);
   U82 : OAI21_X1 port map( B1 => A(10), B2 => n22, A => B(10), ZN => n153);
   U83 : OAI21_X1 port map( B1 => n3, B2 => n31, A => n174, ZN => n222);
   U84 : OAI21_X1 port map( B1 => A(29), B2 => n173, A => B(29), ZN => n174);
   U85 : AOI21_X1 port map( B1 => n237, B2 => A(9), A => n23, ZN => n154);
   U86 : INV_X1 port map( A => n152, ZN => n23);
   U87 : OAI21_X1 port map( B1 => A(9), B2 => n237, A => B(9), ZN => n152);
   U88 : AOI21_X1 port map( B1 => n222, B2 => A(30), A => n2, ZN => n177);
   U89 : INV_X1 port map( A => n175, ZN => n2);
   U90 : OAI21_X1 port map( B1 => A(30), B2 => n222, A => B(30), ZN => n175);
   U91 : AOI22_X1 port map( A1 => n29, A2 => A(3), B1 => n146, B2 => B(3), ZN 
                           => n227);
   U92 : OR2_X1 port map( A1 => A(3), A2 => n29, ZN => n146);
   U93 : INV_X1 port map( A => n225, ZN => n29);
   U94 : OAI21_X1 port map( B1 => n217, B2 => n32, A => n172, ZN => n173);
   U95 : INV_X1 port map( A => A(28), ZN => n32);
   U96 : OAI21_X1 port map( B1 => A(28), B2 => n4, A => B(28), ZN => n172);
   U97 : INV_X1 port map( A => n217, ZN => n4);
   U98 : XNOR2_X1 port map( A => n235, B => n234, ZN => S(8));
   U99 : XNOR2_X1 port map( A => n183, B => n182, ZN => S(12));
   U100 : XNOR2_X1 port map( A => n187, B => n186, ZN => S(14));
   U101 : XNOR2_X1 port map( A => n191, B => n190, ZN => S(16));
   U102 : XNOR2_X1 port map( A => n195, B => n194, ZN => S(18));
   U103 : XNOR2_X1 port map( A => n201, B => n200, ZN => S(20));
   U104 : XNOR2_X1 port map( A => n205, B => n204, ZN => S(22));
   U105 : XNOR2_X1 port map( A => n209, B => n208, ZN => S(24));
   U106 : XNOR2_X1 port map( A => n213, B => n212, ZN => S(26));
   U107 : XNOR2_X1 port map( A => n217, B => n216, ZN => S(28));
   U108 : XNOR2_X1 port map( A => n231, B => n230, ZN => S(6));
   U109 : AOI22_X1 port map( A1 => n46, A2 => A(1), B1 => n144, B2 => B(1), ZN 
                           => n220);
   U110 : OR2_X1 port map( A1 => A(1), A2 => n46, ZN => n144);
   U111 : INV_X1 port map( A => n199, ZN => n46);
   U112 : AOI22_X1 port map( A1 => n45, A2 => A(2), B1 => n145, B2 => B(2), ZN 
                           => n225);
   U113 : OR2_X1 port map( A1 => A(2), A2 => n45, ZN => n145);
   U114 : INV_X1 port map( A => n220, ZN => n45);
   U115 : OAI21_X1 port map( B1 => A(31), B2 => n1, A => B(31), ZN => n176);
   U116 : OAI21_X1 port map( B1 => n227, B2 => n44, A => n147, ZN => n229);
   U117 : INV_X1 port map( A => A(4), ZN => n44);
   U118 : OAI21_X1 port map( B1 => A(4), B2 => n28, A => B(4), ZN => n147);
   U119 : INV_X1 port map( A => n227, ZN => n28);
   U120 : XNOR2_X1 port map( A => n199, B => n198, ZN => S(1));
   U121 : XNOR2_X1 port map( A => n220, B => n219, ZN => S(2));
   U122 : XNOR2_X1 port map( A => n225, B => n224, ZN => S(3));
   U123 : XNOR2_X1 port map( A => n227, B => n226, ZN => S(4));
   U124 : INV_X1 port map( A => A(29), ZN => n31);
   U125 : INV_X1 port map( A => A(31), ZN => n30);
   U126 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n47, ZN => n199);
   U127 : INV_X1 port map( A => n143, ZN => n47);
   U128 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n143);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_N32_0;

architecture SYN_BEHAVIORAL of RCA_N32_0 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237 : std_logic;

begin
   
   U129 : XOR2_X1 port map( A => n237, B => n236, Z => S(9));
   U130 : XOR2_X1 port map( A => B(9), B => A(9), Z => n236);
   U131 : XOR2_X1 port map( A => B(8), B => A(8), Z => n234);
   U132 : XOR2_X1 port map( A => n233, B => n232, Z => S(7));
   U133 : XOR2_X1 port map( A => B(7), B => A(7), Z => n232);
   U134 : XOR2_X1 port map( A => B(6), B => A(6), Z => n230);
   U135 : XOR2_X1 port map( A => n229, B => n228, Z => S(5));
   U136 : XOR2_X1 port map( A => B(5), B => A(5), Z => n228);
   U137 : XOR2_X1 port map( A => B(4), B => A(4), Z => n226);
   U138 : XOR2_X1 port map( A => B(3), B => A(3), Z => n224);
   U139 : XOR2_X1 port map( A => n1, B => n223, Z => S(31));
   U140 : XOR2_X1 port map( A => B(31), B => A(31), Z => n223);
   U141 : XOR2_X1 port map( A => n222, B => n221, Z => S(30));
   U142 : XOR2_X1 port map( A => B(30), B => A(30), Z => n221);
   U143 : XOR2_X1 port map( A => B(2), B => A(2), Z => n219);
   U144 : XOR2_X1 port map( A => B(28), B => A(28), Z => n216);
   U145 : XOR2_X1 port map( A => n215, B => n214, Z => S(27));
   U146 : XOR2_X1 port map( A => B(27), B => A(27), Z => n214);
   U147 : XOR2_X1 port map( A => B(26), B => A(26), Z => n212);
   U148 : XOR2_X1 port map( A => n211, B => n210, Z => S(25));
   U149 : XOR2_X1 port map( A => B(25), B => A(25), Z => n210);
   U150 : XOR2_X1 port map( A => B(24), B => A(24), Z => n208);
   U151 : XOR2_X1 port map( A => n207, B => n206, Z => S(23));
   U152 : XOR2_X1 port map( A => B(23), B => A(23), Z => n206);
   U153 : XOR2_X1 port map( A => B(22), B => A(22), Z => n204);
   U154 : XOR2_X1 port map( A => n203, B => n202, Z => S(21));
   U155 : XOR2_X1 port map( A => B(21), B => A(21), Z => n202);
   U156 : XOR2_X1 port map( A => B(20), B => A(20), Z => n200);
   U157 : XOR2_X1 port map( A => B(1), B => A(1), Z => n198);
   U158 : XOR2_X1 port map( A => n197, B => n196, Z => S(19));
   U159 : XOR2_X1 port map( A => B(19), B => A(19), Z => n196);
   U160 : XOR2_X1 port map( A => B(18), B => A(18), Z => n194);
   U161 : XOR2_X1 port map( A => n193, B => n192, Z => S(17));
   U162 : XOR2_X1 port map( A => B(17), B => A(17), Z => n192);
   U163 : XOR2_X1 port map( A => B(16), B => A(16), Z => n190);
   U164 : XOR2_X1 port map( A => n189, B => n188, Z => S(15));
   U165 : XOR2_X1 port map( A => B(15), B => A(15), Z => n188);
   U166 : XOR2_X1 port map( A => B(14), B => A(14), Z => n186);
   U167 : XOR2_X1 port map( A => n185, B => n184, Z => S(13));
   U168 : XOR2_X1 port map( A => B(13), B => A(13), Z => n184);
   U169 : XOR2_X1 port map( A => B(12), B => A(12), Z => n182);
   U170 : XOR2_X1 port map( A => n181, B => n180, Z => S(11));
   U171 : XOR2_X1 port map( A => B(11), B => A(11), Z => n180);
   U172 : XOR2_X1 port map( A => n22, B => n179, Z => S(10));
   U173 : XOR2_X1 port map( A => B(10), B => A(10), Z => n179);
   U174 : XOR2_X1 port map( A => A(0), B => n178, Z => S(0));
   U175 : XOR2_X1 port map( A => Ci, B => B(0), Z => n178);
   U1 : XNOR2_X1 port map( A => n3, B => n218, ZN => S(29));
   U2 : XNOR2_X1 port map( A => B(29), B => n31, ZN => n218);
   U3 : INV_X1 port map( A => n173, ZN => n3);
   U4 : OAI21_X1 port map( B1 => n177, B2 => n30, A => n176, ZN => Co);
   U5 : INV_X1 port map( A => n154, ZN => n22);
   U6 : INV_X1 port map( A => n177, ZN => n1);
   U7 : AOI21_X1 port map( B1 => n233, B2 => A(7), A => n25, ZN => n235);
   U8 : INV_X1 port map( A => n150, ZN => n25);
   U9 : OAI21_X1 port map( B1 => A(7), B2 => n233, A => B(7), ZN => n150);
   U10 : AOI21_X1 port map( B1 => n181, B2 => A(11), A => n21, ZN => n183);
   U11 : INV_X1 port map( A => n155, ZN => n21);
   U12 : OAI21_X1 port map( B1 => A(11), B2 => n181, A => B(11), ZN => n155);
   U13 : AOI21_X1 port map( B1 => n185, B2 => A(13), A => n19, ZN => n187);
   U14 : INV_X1 port map( A => n157, ZN => n19);
   U15 : OAI21_X1 port map( B1 => A(13), B2 => n185, A => B(13), ZN => n157);
   U16 : AOI21_X1 port map( B1 => n189, B2 => A(15), A => n17, ZN => n191);
   U17 : INV_X1 port map( A => n159, ZN => n17);
   U18 : OAI21_X1 port map( B1 => A(15), B2 => n189, A => B(15), ZN => n159);
   U19 : AOI21_X1 port map( B1 => n193, B2 => A(17), A => n15, ZN => n195);
   U20 : INV_X1 port map( A => n161, ZN => n15);
   U21 : OAI21_X1 port map( B1 => A(17), B2 => n193, A => B(17), ZN => n161);
   U22 : AOI21_X1 port map( B1 => n197, B2 => A(19), A => n13, ZN => n201);
   U23 : INV_X1 port map( A => n163, ZN => n13);
   U24 : OAI21_X1 port map( B1 => A(19), B2 => n197, A => B(19), ZN => n163);
   U25 : AOI21_X1 port map( B1 => n203, B2 => A(21), A => n11, ZN => n205);
   U26 : INV_X1 port map( A => n165, ZN => n11);
   U27 : OAI21_X1 port map( B1 => A(21), B2 => n203, A => B(21), ZN => n165);
   U28 : AOI21_X1 port map( B1 => n207, B2 => A(23), A => n9, ZN => n209);
   U29 : INV_X1 port map( A => n167, ZN => n9);
   U30 : OAI21_X1 port map( B1 => A(23), B2 => n207, A => B(23), ZN => n167);
   U31 : AOI21_X1 port map( B1 => n211, B2 => A(25), A => n7, ZN => n213);
   U32 : INV_X1 port map( A => n169, ZN => n7);
   U33 : OAI21_X1 port map( B1 => A(25), B2 => n211, A => B(25), ZN => n169);
   U34 : AOI21_X1 port map( B1 => n215, B2 => A(27), A => n5, ZN => n217);
   U35 : INV_X1 port map( A => n171, ZN => n5);
   U36 : OAI21_X1 port map( B1 => A(27), B2 => n215, A => B(27), ZN => n171);
   U37 : AOI21_X1 port map( B1 => n229, B2 => A(5), A => n27, ZN => n231);
   U38 : INV_X1 port map( A => n148, ZN => n27);
   U39 : OAI21_X1 port map( B1 => A(5), B2 => n229, A => B(5), ZN => n148);
   U40 : OAI21_X1 port map( B1 => n183, B2 => n40, A => n156, ZN => n185);
   U41 : INV_X1 port map( A => A(12), ZN => n40);
   U42 : OAI21_X1 port map( B1 => A(12), B2 => n20, A => B(12), ZN => n156);
   U43 : INV_X1 port map( A => n183, ZN => n20);
   U44 : OAI21_X1 port map( B1 => n187, B2 => n39, A => n158, ZN => n189);
   U45 : INV_X1 port map( A => A(14), ZN => n39);
   U46 : OAI21_X1 port map( B1 => A(14), B2 => n18, A => B(14), ZN => n158);
   U47 : INV_X1 port map( A => n187, ZN => n18);
   U48 : OAI21_X1 port map( B1 => n191, B2 => n38, A => n160, ZN => n193);
   U49 : INV_X1 port map( A => A(16), ZN => n38);
   U50 : OAI21_X1 port map( B1 => A(16), B2 => n16, A => B(16), ZN => n160);
   U51 : INV_X1 port map( A => n191, ZN => n16);
   U52 : OAI21_X1 port map( B1 => n195, B2 => n37, A => n162, ZN => n197);
   U53 : INV_X1 port map( A => A(18), ZN => n37);
   U54 : OAI21_X1 port map( B1 => A(18), B2 => n14, A => B(18), ZN => n162);
   U55 : INV_X1 port map( A => n195, ZN => n14);
   U56 : OAI21_X1 port map( B1 => n201, B2 => n36, A => n164, ZN => n203);
   U57 : INV_X1 port map( A => A(20), ZN => n36);
   U58 : OAI21_X1 port map( B1 => A(20), B2 => n12, A => B(20), ZN => n164);
   U59 : INV_X1 port map( A => n201, ZN => n12);
   U60 : OAI21_X1 port map( B1 => n205, B2 => n35, A => n166, ZN => n207);
   U61 : INV_X1 port map( A => A(22), ZN => n35);
   U62 : OAI21_X1 port map( B1 => A(22), B2 => n10, A => B(22), ZN => n166);
   U63 : INV_X1 port map( A => n205, ZN => n10);
   U64 : OAI21_X1 port map( B1 => n209, B2 => n34, A => n168, ZN => n211);
   U65 : INV_X1 port map( A => A(24), ZN => n34);
   U66 : OAI21_X1 port map( B1 => A(24), B2 => n8, A => B(24), ZN => n168);
   U67 : INV_X1 port map( A => n209, ZN => n8);
   U68 : OAI21_X1 port map( B1 => n213, B2 => n33, A => n170, ZN => n215);
   U69 : INV_X1 port map( A => A(26), ZN => n33);
   U70 : OAI21_X1 port map( B1 => A(26), B2 => n6, A => B(26), ZN => n170);
   U71 : INV_X1 port map( A => n213, ZN => n6);
   U72 : OAI21_X1 port map( B1 => n227, B2 => n47, A => n147, ZN => n229);
   U73 : INV_X1 port map( A => A(4), ZN => n47);
   U74 : OAI21_X1 port map( B1 => A(4), B2 => n28, A => B(4), ZN => n147);
   U75 : INV_X1 port map( A => n227, ZN => n28);
   U76 : OAI21_X1 port map( B1 => n235, B2 => n42, A => n151, ZN => n237);
   U77 : INV_X1 port map( A => A(8), ZN => n42);
   U78 : OAI21_X1 port map( B1 => A(8), B2 => n24, A => B(8), ZN => n151);
   U79 : INV_X1 port map( A => n235, ZN => n24);
   U80 : OAI21_X1 port map( B1 => n154, B2 => n41, A => n153, ZN => n181);
   U81 : INV_X1 port map( A => A(10), ZN => n41);
   U82 : OAI21_X1 port map( B1 => A(10), B2 => n22, A => B(10), ZN => n153);
   U83 : OAI21_X1 port map( B1 => n3, B2 => n31, A => n174, ZN => n222);
   U84 : OAI21_X1 port map( B1 => A(29), B2 => n173, A => B(29), ZN => n174);
   U85 : AOI21_X1 port map( B1 => n237, B2 => A(9), A => n23, ZN => n154);
   U86 : INV_X1 port map( A => n152, ZN => n23);
   U87 : OAI21_X1 port map( B1 => A(9), B2 => n237, A => B(9), ZN => n152);
   U88 : AOI21_X1 port map( B1 => n222, B2 => A(30), A => n2, ZN => n177);
   U89 : INV_X1 port map( A => n175, ZN => n2);
   U90 : OAI21_X1 port map( B1 => A(30), B2 => n222, A => B(30), ZN => n175);
   U91 : AOI22_X1 port map( A1 => n29, A2 => A(3), B1 => n146, B2 => B(3), ZN 
                           => n227);
   U92 : OR2_X1 port map( A1 => A(3), A2 => n29, ZN => n146);
   U93 : INV_X1 port map( A => n225, ZN => n29);
   U94 : OAI21_X1 port map( B1 => n217, B2 => n32, A => n172, ZN => n173);
   U95 : INV_X1 port map( A => A(28), ZN => n32);
   U96 : OAI21_X1 port map( B1 => A(28), B2 => n4, A => B(28), ZN => n172);
   U97 : INV_X1 port map( A => n217, ZN => n4);
   U98 : AOI22_X1 port map( A1 => n45, A2 => A(1), B1 => n144, B2 => B(1), ZN 
                           => n220);
   U99 : OR2_X1 port map( A1 => A(1), A2 => n45, ZN => n144);
   U100 : INV_X1 port map( A => n199, ZN => n45);
   U101 : AOI22_X1 port map( A1 => n44, A2 => A(2), B1 => n145, B2 => B(2), ZN 
                           => n225);
   U102 : OR2_X1 port map( A1 => A(2), A2 => n44, ZN => n145);
   U103 : INV_X1 port map( A => n220, ZN => n44);
   U104 : OAI21_X1 port map( B1 => A(31), B2 => n1, A => B(31), ZN => n176);
   U105 : XNOR2_X1 port map( A => n183, B => n182, ZN => S(12));
   U106 : XNOR2_X1 port map( A => n187, B => n186, ZN => S(14));
   U107 : XNOR2_X1 port map( A => n191, B => n190, ZN => S(16));
   U108 : XNOR2_X1 port map( A => n195, B => n194, ZN => S(18));
   U109 : XNOR2_X1 port map( A => n201, B => n200, ZN => S(20));
   U110 : XNOR2_X1 port map( A => n205, B => n204, ZN => S(22));
   U111 : XNOR2_X1 port map( A => n209, B => n208, ZN => S(24));
   U112 : XNOR2_X1 port map( A => n213, B => n212, ZN => S(26));
   U113 : XNOR2_X1 port map( A => n217, B => n216, ZN => S(28));
   U114 : XNOR2_X1 port map( A => n235, B => n234, ZN => S(8));
   U115 : OAI21_X1 port map( B1 => n231, B2 => n43, A => n149, ZN => n233);
   U116 : INV_X1 port map( A => A(6), ZN => n43);
   U117 : OAI21_X1 port map( B1 => A(6), B2 => n26, A => B(6), ZN => n149);
   U118 : INV_X1 port map( A => n231, ZN => n26);
   U119 : INV_X1 port map( A => A(29), ZN => n31);
   U120 : XNOR2_X1 port map( A => n199, B => n198, ZN => S(1));
   U121 : XNOR2_X1 port map( A => n220, B => n219, ZN => S(2));
   U122 : XNOR2_X1 port map( A => n225, B => n224, ZN => S(3));
   U123 : XNOR2_X1 port map( A => n227, B => n226, ZN => S(4));
   U124 : XNOR2_X1 port map( A => n231, B => n230, ZN => S(6));
   U125 : INV_X1 port map( A => A(31), ZN => n30);
   U126 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n46, ZN => n199);
   U127 : INV_X1 port map( A => n143, ZN => n46);
   U128 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n143);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX81_N32_2 is

   port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX81_N32_2;

architecture SYN_BEHAVIORAL of MUX81_N32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n298, Z => n152);
   U2 : BUF_X1 port map( A => n297, Z => n148);
   U3 : BUF_X1 port map( A => n296, Z => n144);
   U4 : BUF_X1 port map( A => n295, Z => n140);
   U5 : BUF_X1 port map( A => n300, Z => n157);
   U6 : BUF_X1 port map( A => n299, Z => n153);
   U7 : BUF_X1 port map( A => n302, Z => n165);
   U8 : BUF_X1 port map( A => n301, Z => n161);
   U9 : AOI22_X1 port map( A1 => D(18), A2 => n149, B1 => C(18), B2 => n145, ZN
                           => n209);
   U10 : AOI22_X1 port map( A1 => D(19), A2 => n149, B1 => C(19), B2 => n145, 
                           ZN => n213);
   U11 : AOI22_X1 port map( A1 => D(20), A2 => n150, B1 => C(20), B2 => n146, 
                           ZN => n221);
   U12 : AOI22_X1 port map( A1 => D(21), A2 => n150, B1 => C(21), B2 => n146, 
                           ZN => n225);
   U13 : AOI22_X1 port map( A1 => D(22), A2 => n150, B1 => C(22), B2 => n146, 
                           ZN => n229);
   U14 : AOI22_X1 port map( A1 => D(23), A2 => n150, B1 => C(23), B2 => n146, 
                           ZN => n233);
   U15 : AOI22_X1 port map( A1 => D(24), A2 => n150, B1 => C(24), B2 => n146, 
                           ZN => n237);
   U16 : AOI22_X1 port map( A1 => D(25), A2 => n150, B1 => C(25), B2 => n146, 
                           ZN => n241);
   U17 : AOI22_X1 port map( A1 => D(26), A2 => n150, B1 => C(26), B2 => n146, 
                           ZN => n245);
   U18 : AOI22_X1 port map( A1 => D(27), A2 => n150, B1 => C(27), B2 => n146, 
                           ZN => n249);
   U19 : AOI22_X1 port map( A1 => D(28), A2 => n150, B1 => C(28), B2 => n146, 
                           ZN => n253);
   U20 : AOI22_X1 port map( A1 => D(29), A2 => n150, B1 => C(29), B2 => n146, 
                           ZN => n257);
   U21 : AOI22_X1 port map( A1 => D(30), A2 => n150, B1 => C(30), B2 => n146, 
                           ZN => n265);
   U22 : AOI22_X1 port map( A1 => D(31), A2 => n151, B1 => C(31), B2 => n147, 
                           ZN => n269);
   U23 : INV_X1 port map( A => S(1), ZN => n169);
   U24 : BUF_X1 port map( A => n152, Z => n149);
   U25 : BUF_X1 port map( A => n144, Z => n141);
   U26 : BUF_X1 port map( A => n152, Z => n150);
   U27 : BUF_X1 port map( A => n144, Z => n142);
   U28 : BUF_X1 port map( A => n157, Z => n158);
   U29 : BUF_X1 port map( A => n165, Z => n166);
   U30 : BUF_X1 port map( A => n157, Z => n159);
   U31 : BUF_X1 port map( A => n165, Z => n167);
   U32 : BUF_X1 port map( A => n148, Z => n145);
   U33 : BUF_X1 port map( A => n140, Z => n1);
   U34 : BUF_X1 port map( A => n148, Z => n146);
   U35 : BUF_X1 port map( A => n140, Z => n2);
   U36 : BUF_X1 port map( A => n153, Z => n154);
   U37 : BUF_X1 port map( A => n161, Z => n162);
   U38 : BUF_X1 port map( A => n153, Z => n155);
   U39 : BUF_X1 port map( A => n161, Z => n163);
   U40 : BUF_X1 port map( A => n152, Z => n151);
   U41 : BUF_X1 port map( A => n144, Z => n143);
   U42 : BUF_X1 port map( A => n148, Z => n147);
   U43 : BUF_X1 port map( A => n140, Z => n139);
   U44 : BUF_X1 port map( A => n157, Z => n160);
   U45 : BUF_X1 port map( A => n165, Z => n168);
   U46 : BUF_X1 port map( A => n153, Z => n156);
   U47 : BUF_X1 port map( A => n161, Z => n164);
   U48 : AOI22_X1 port map( A1 => D(3), A2 => n151, B1 => C(3), B2 => n147, ZN 
                           => n273);
   U49 : AOI22_X1 port map( A1 => D(4), A2 => n151, B1 => C(4), B2 => n147, ZN 
                           => n277);
   U50 : AOI22_X1 port map( A1 => D(5), A2 => n151, B1 => C(5), B2 => n147, ZN 
                           => n281);
   U51 : AOI22_X1 port map( A1 => D(6), A2 => n151, B1 => C(6), B2 => n147, ZN 
                           => n285);
   U52 : AOI22_X1 port map( A1 => D(7), A2 => n151, B1 => C(7), B2 => n147, ZN 
                           => n289);
   U53 : AOI22_X1 port map( A1 => D(8), A2 => n151, B1 => C(8), B2 => n147, ZN 
                           => n293);
   U54 : AOI22_X1 port map( A1 => D(9), A2 => n151, B1 => C(9), B2 => n147, ZN 
                           => n305);
   U55 : AOI22_X1 port map( A1 => D(10), A2 => n149, B1 => C(10), B2 => n145, 
                           ZN => n177);
   U56 : AOI22_X1 port map( A1 => D(11), A2 => n149, B1 => C(11), B2 => n145, 
                           ZN => n181);
   U57 : AOI22_X1 port map( A1 => D(12), A2 => n149, B1 => C(12), B2 => n145, 
                           ZN => n185);
   U58 : AOI22_X1 port map( A1 => D(13), A2 => n149, B1 => C(13), B2 => n145, 
                           ZN => n189);
   U59 : AOI22_X1 port map( A1 => D(14), A2 => n149, B1 => C(14), B2 => n145, 
                           ZN => n193);
   U60 : AOI22_X1 port map( A1 => D(15), A2 => n149, B1 => C(15), B2 => n145, 
                           ZN => n197);
   U61 : AOI22_X1 port map( A1 => D(16), A2 => n149, B1 => C(16), B2 => n145, 
                           ZN => n201);
   U62 : AOI22_X1 port map( A1 => D(17), A2 => n149, B1 => C(17), B2 => n145, 
                           ZN => n205);
   U63 : INV_X1 port map( A => S(0), ZN => n170);
   U64 : NOR3_X1 port map( A1 => n170, A2 => S(2), A3 => n169, ZN => n298);
   U65 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n169, ZN => n297);
   U66 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n170, ZN => n296);
   U67 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => S(0), ZN => n295);
   U68 : AND3_X1 port map( A1 => S(0), A2 => n169, A3 => S(2), ZN => n300);
   U69 : AND3_X1 port map( A1 => n170, A2 => n169, A3 => S(2), ZN => n299);
   U70 : AND3_X1 port map( A1 => S(1), A2 => S(0), A3 => S(2), ZN => n302);
   U71 : AND3_X1 port map( A1 => S(1), A2 => n170, A3 => S(2), ZN => n301);
   U72 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(19));
   U73 : AOI22_X1 port map( A1 => H(19), A2 => n166, B1 => G(19), B2 => n162, 
                           ZN => n211);
   U74 : AOI22_X1 port map( A1 => B(19), A2 => n141, B1 => A(19), B2 => n1, ZN 
                           => n214);
   U75 : AOI22_X1 port map( A1 => F(19), A2 => n158, B1 => E(19), B2 => n154, 
                           ZN => n212);
   U76 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN 
                           => Y(21));
   U77 : AOI22_X1 port map( A1 => H(21), A2 => n167, B1 => G(21), B2 => n163, 
                           ZN => n223);
   U78 : AOI22_X1 port map( A1 => B(21), A2 => n142, B1 => A(21), B2 => n2, ZN 
                           => n226);
   U79 : AOI22_X1 port map( A1 => F(21), A2 => n159, B1 => E(21), B2 => n155, 
                           ZN => n224);
   U80 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN 
                           => Y(23));
   U81 : AOI22_X1 port map( A1 => H(23), A2 => n167, B1 => G(23), B2 => n163, 
                           ZN => n231);
   U82 : AOI22_X1 port map( A1 => B(23), A2 => n142, B1 => A(23), B2 => n2, ZN 
                           => n234);
   U83 : AOI22_X1 port map( A1 => F(23), A2 => n159, B1 => E(23), B2 => n155, 
                           ZN => n232);
   U84 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN 
                           => Y(25));
   U85 : AOI22_X1 port map( A1 => H(25), A2 => n167, B1 => G(25), B2 => n163, 
                           ZN => n239);
   U86 : AOI22_X1 port map( A1 => B(25), A2 => n142, B1 => A(25), B2 => n2, ZN 
                           => n242);
   U87 : AOI22_X1 port map( A1 => F(25), A2 => n159, B1 => E(25), B2 => n155, 
                           ZN => n240);
   U88 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN 
                           => Y(27));
   U89 : AOI22_X1 port map( A1 => H(27), A2 => n167, B1 => G(27), B2 => n163, 
                           ZN => n247);
   U90 : AOI22_X1 port map( A1 => B(27), A2 => n142, B1 => A(27), B2 => n2, ZN 
                           => n250);
   U91 : AOI22_X1 port map( A1 => F(27), A2 => n159, B1 => E(27), B2 => n155, 
                           ZN => n248);
   U92 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN 
                           => Y(30));
   U93 : AOI22_X1 port map( A1 => H(30), A2 => n167, B1 => G(30), B2 => n163, 
                           ZN => n263);
   U94 : AOI22_X1 port map( A1 => B(30), A2 => n142, B1 => A(30), B2 => n2, ZN 
                           => n266);
   U95 : AOI22_X1 port map( A1 => F(30), A2 => n159, B1 => E(30), B2 => n155, 
                           ZN => n264);
   U96 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(18));
   U97 : AOI22_X1 port map( A1 => H(18), A2 => n166, B1 => G(18), B2 => n162, 
                           ZN => n207);
   U98 : AOI22_X1 port map( A1 => B(18), A2 => n141, B1 => A(18), B2 => n1, ZN 
                           => n210);
   U99 : AOI22_X1 port map( A1 => F(18), A2 => n158, B1 => E(18), B2 => n154, 
                           ZN => n208);
   U100 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(20));
   U101 : AOI22_X1 port map( A1 => H(20), A2 => n167, B1 => G(20), B2 => n163, 
                           ZN => n219);
   U102 : AOI22_X1 port map( A1 => B(20), A2 => n142, B1 => A(20), B2 => n2, ZN
                           => n222);
   U103 : AOI22_X1 port map( A1 => F(20), A2 => n159, B1 => E(20), B2 => n155, 
                           ZN => n220);
   U104 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(22));
   U105 : AOI22_X1 port map( A1 => H(22), A2 => n167, B1 => G(22), B2 => n163, 
                           ZN => n227);
   U106 : AOI22_X1 port map( A1 => B(22), A2 => n142, B1 => A(22), B2 => n2, ZN
                           => n230);
   U107 : AOI22_X1 port map( A1 => F(22), A2 => n159, B1 => E(22), B2 => n155, 
                           ZN => n228);
   U108 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(24));
   U109 : AOI22_X1 port map( A1 => H(24), A2 => n167, B1 => G(24), B2 => n163, 
                           ZN => n235);
   U110 : AOI22_X1 port map( A1 => B(24), A2 => n142, B1 => A(24), B2 => n2, ZN
                           => n238);
   U111 : AOI22_X1 port map( A1 => F(24), A2 => n159, B1 => E(24), B2 => n155, 
                           ZN => n236);
   U112 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(26));
   U113 : AOI22_X1 port map( A1 => H(26), A2 => n167, B1 => G(26), B2 => n163, 
                           ZN => n243);
   U114 : AOI22_X1 port map( A1 => B(26), A2 => n142, B1 => A(26), B2 => n2, ZN
                           => n246);
   U115 : AOI22_X1 port map( A1 => F(26), A2 => n159, B1 => E(26), B2 => n155, 
                           ZN => n244);
   U116 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(28));
   U117 : AOI22_X1 port map( A1 => H(28), A2 => n167, B1 => G(28), B2 => n163, 
                           ZN => n251);
   U118 : AOI22_X1 port map( A1 => B(28), A2 => n142, B1 => A(28), B2 => n2, ZN
                           => n254);
   U119 : AOI22_X1 port map( A1 => F(28), A2 => n159, B1 => E(28), B2 => n155, 
                           ZN => n252);
   U120 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(31));
   U121 : AOI22_X1 port map( A1 => H(31), A2 => n168, B1 => G(31), B2 => n164, 
                           ZN => n267);
   U122 : AOI22_X1 port map( A1 => B(31), A2 => n143, B1 => A(31), B2 => n139, 
                           ZN => n270);
   U123 : AOI22_X1 port map( A1 => F(31), A2 => n160, B1 => E(31), B2 => n156, 
                           ZN => n268);
   U124 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(5));
   U125 : AOI22_X1 port map( A1 => H(5), A2 => n168, B1 => G(5), B2 => n164, ZN
                           => n279);
   U126 : AOI22_X1 port map( A1 => B(5), A2 => n143, B1 => A(5), B2 => n139, ZN
                           => n282);
   U127 : AOI22_X1 port map( A1 => F(5), A2 => n160, B1 => E(5), B2 => n156, ZN
                           => n280);
   U128 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(7));
   U129 : AOI22_X1 port map( A1 => H(7), A2 => n168, B1 => G(7), B2 => n164, ZN
                           => n287);
   U130 : AOI22_X1 port map( A1 => B(7), A2 => n143, B1 => A(7), B2 => n139, ZN
                           => n290);
   U131 : AOI22_X1 port map( A1 => F(7), A2 => n160, B1 => E(7), B2 => n156, ZN
                           => n288);
   U132 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(9));
   U133 : AOI22_X1 port map( A1 => H(9), A2 => n168, B1 => G(9), B2 => n164, ZN
                           => n303);
   U134 : AOI22_X1 port map( A1 => B(9), A2 => n143, B1 => A(9), B2 => n139, ZN
                           => n306);
   U135 : AOI22_X1 port map( A1 => F(9), A2 => n160, B1 => E(9), B2 => n156, ZN
                           => n304);
   U136 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN
                           => Y(11));
   U137 : AOI22_X1 port map( A1 => H(11), A2 => n166, B1 => G(11), B2 => n162, 
                           ZN => n179);
   U138 : AOI22_X1 port map( A1 => B(11), A2 => n141, B1 => A(11), B2 => n1, ZN
                           => n182);
   U139 : AOI22_X1 port map( A1 => F(11), A2 => n158, B1 => E(11), B2 => n154, 
                           ZN => n180);
   U140 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN
                           => Y(13));
   U141 : AOI22_X1 port map( A1 => H(13), A2 => n166, B1 => G(13), B2 => n162, 
                           ZN => n187);
   U142 : AOI22_X1 port map( A1 => B(13), A2 => n141, B1 => A(13), B2 => n1, ZN
                           => n190);
   U143 : AOI22_X1 port map( A1 => F(13), A2 => n158, B1 => E(13), B2 => n154, 
                           ZN => n188);
   U144 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN
                           => Y(15));
   U145 : AOI22_X1 port map( A1 => H(15), A2 => n166, B1 => G(15), B2 => n162, 
                           ZN => n195);
   U146 : AOI22_X1 port map( A1 => B(15), A2 => n141, B1 => A(15), B2 => n1, ZN
                           => n198);
   U147 : AOI22_X1 port map( A1 => F(15), A2 => n158, B1 => E(15), B2 => n154, 
                           ZN => n196);
   U148 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN
                           => Y(17));
   U149 : AOI22_X1 port map( A1 => H(17), A2 => n166, B1 => G(17), B2 => n162, 
                           ZN => n203);
   U150 : AOI22_X1 port map( A1 => B(17), A2 => n141, B1 => A(17), B2 => n1, ZN
                           => n206);
   U151 : AOI22_X1 port map( A1 => F(17), A2 => n158, B1 => E(17), B2 => n154, 
                           ZN => n204);
   U152 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(4));
   U153 : AOI22_X1 port map( A1 => H(4), A2 => n168, B1 => G(4), B2 => n164, ZN
                           => n275);
   U154 : AOI22_X1 port map( A1 => B(4), A2 => n143, B1 => A(4), B2 => n139, ZN
                           => n278);
   U155 : AOI22_X1 port map( A1 => F(4), A2 => n160, B1 => E(4), B2 => n156, ZN
                           => n276);
   U156 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(6));
   U157 : AOI22_X1 port map( A1 => H(6), A2 => n168, B1 => G(6), B2 => n164, ZN
                           => n283);
   U158 : AOI22_X1 port map( A1 => B(6), A2 => n143, B1 => A(6), B2 => n139, ZN
                           => n286);
   U159 : AOI22_X1 port map( A1 => F(6), A2 => n160, B1 => E(6), B2 => n156, ZN
                           => n284);
   U160 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(8));
   U161 : AOI22_X1 port map( A1 => H(8), A2 => n168, B1 => G(8), B2 => n164, ZN
                           => n291);
   U162 : AOI22_X1 port map( A1 => B(8), A2 => n143, B1 => A(8), B2 => n139, ZN
                           => n294);
   U163 : AOI22_X1 port map( A1 => F(8), A2 => n160, B1 => E(8), B2 => n156, ZN
                           => n292);
   U164 : NAND4_X1 port map( A1 => n178, A2 => n177, A3 => n176, A4 => n175, ZN
                           => Y(10));
   U165 : AOI22_X1 port map( A1 => H(10), A2 => n166, B1 => G(10), B2 => n162, 
                           ZN => n175);
   U166 : AOI22_X1 port map( A1 => B(10), A2 => n141, B1 => A(10), B2 => n1, ZN
                           => n178);
   U167 : AOI22_X1 port map( A1 => F(10), A2 => n158, B1 => E(10), B2 => n154, 
                           ZN => n176);
   U168 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN
                           => Y(12));
   U169 : AOI22_X1 port map( A1 => H(12), A2 => n166, B1 => G(12), B2 => n162, 
                           ZN => n183);
   U170 : AOI22_X1 port map( A1 => B(12), A2 => n141, B1 => A(12), B2 => n1, ZN
                           => n186);
   U171 : AOI22_X1 port map( A1 => F(12), A2 => n158, B1 => E(12), B2 => n154, 
                           ZN => n184);
   U172 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN
                           => Y(14));
   U173 : AOI22_X1 port map( A1 => H(14), A2 => n166, B1 => G(14), B2 => n162, 
                           ZN => n191);
   U174 : AOI22_X1 port map( A1 => B(14), A2 => n141, B1 => A(14), B2 => n1, ZN
                           => n194);
   U175 : AOI22_X1 port map( A1 => F(14), A2 => n158, B1 => E(14), B2 => n154, 
                           ZN => n192);
   U176 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN
                           => Y(16));
   U177 : AOI22_X1 port map( A1 => H(16), A2 => n166, B1 => G(16), B2 => n162, 
                           ZN => n199);
   U178 : AOI22_X1 port map( A1 => B(16), A2 => n141, B1 => A(16), B2 => n1, ZN
                           => n202);
   U179 : AOI22_X1 port map( A1 => F(16), A2 => n158, B1 => E(16), B2 => n154, 
                           ZN => n200);
   U180 : NAND4_X1 port map( A1 => n174, A2 => n173, A3 => n172, A4 => n171, ZN
                           => Y(0));
   U181 : AOI22_X1 port map( A1 => B(0), A2 => n141, B1 => A(0), B2 => n1, ZN 
                           => n174);
   U182 : AOI22_X1 port map( A1 => D(0), A2 => n149, B1 => C(0), B2 => n145, ZN
                           => n173);
   U183 : AOI22_X1 port map( A1 => F(0), A2 => n158, B1 => E(0), B2 => n154, ZN
                           => n172);
   U184 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(29));
   U185 : AOI22_X1 port map( A1 => H(29), A2 => n167, B1 => G(29), B2 => n163, 
                           ZN => n255);
   U186 : AOI22_X1 port map( A1 => B(29), A2 => n142, B1 => A(29), B2 => n2, ZN
                           => n258);
   U187 : AOI22_X1 port map( A1 => F(29), A2 => n159, B1 => E(29), B2 => n155, 
                           ZN => n256);
   U188 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(3));
   U189 : AOI22_X1 port map( A1 => H(3), A2 => n168, B1 => G(3), B2 => n164, ZN
                           => n271);
   U190 : AOI22_X1 port map( A1 => B(3), A2 => n143, B1 => A(3), B2 => n139, ZN
                           => n274);
   U191 : AOI22_X1 port map( A1 => F(3), A2 => n160, B1 => E(3), B2 => n156, ZN
                           => n272);
   U192 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(2));
   U193 : AOI22_X1 port map( A1 => F(2), A2 => n159, B1 => E(2), B2 => n155, ZN
                           => n260);
   U194 : AOI22_X1 port map( A1 => H(2), A2 => n167, B1 => G(2), B2 => n163, ZN
                           => n259);
   U195 : AOI22_X1 port map( A1 => B(2), A2 => n142, B1 => A(2), B2 => n2, ZN 
                           => n262);
   U196 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN
                           => Y(1));
   U197 : AOI22_X1 port map( A1 => B(1), A2 => n141, B1 => A(1), B2 => n1, ZN 
                           => n218);
   U198 : AOI22_X1 port map( A1 => D(1), A2 => n149, B1 => C(1), B2 => n145, ZN
                           => n217);
   U199 : AOI22_X1 port map( A1 => F(1), A2 => n158, B1 => E(1), B2 => n154, ZN
                           => n216);
   U200 : AOI22_X1 port map( A1 => D(2), A2 => n150, B1 => C(2), B2 => n146, ZN
                           => n261);
   U201 : AOI22_X1 port map( A1 => H(0), A2 => n166, B1 => G(0), B2 => n162, ZN
                           => n171);
   U202 : AOI22_X1 port map( A1 => H(1), A2 => n166, B1 => G(1), B2 => n162, ZN
                           => n215);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX81_N32_1 is

   port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX81_N32_1;

architecture SYN_BEHAVIORAL of MUX81_N32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n296, Z => n144);
   U2 : BUF_X1 port map( A => n298, Z => n152);
   U3 : BUF_X1 port map( A => n299, Z => n153);
   U4 : BUF_X1 port map( A => n301, Z => n161);
   U5 : BUF_X1 port map( A => n297, Z => n148);
   U6 : BUF_X1 port map( A => n295, Z => n140);
   U7 : BUF_X1 port map( A => n300, Z => n157);
   U8 : BUF_X1 port map( A => n302, Z => n165);
   U9 : AOI22_X1 port map( A1 => D(5), A2 => n151, B1 => C(5), B2 => n147, ZN 
                           => n281);
   U10 : AOI22_X1 port map( A1 => D(6), A2 => n151, B1 => C(6), B2 => n147, ZN 
                           => n285);
   U11 : AOI22_X1 port map( A1 => D(7), A2 => n151, B1 => C(7), B2 => n147, ZN 
                           => n289);
   U12 : AOI22_X1 port map( A1 => D(8), A2 => n151, B1 => C(8), B2 => n147, ZN 
                           => n293);
   U13 : AOI22_X1 port map( A1 => D(9), A2 => n151, B1 => C(9), B2 => n147, ZN 
                           => n305);
   U14 : AOI22_X1 port map( A1 => D(10), A2 => n149, B1 => C(10), B2 => n145, 
                           ZN => n177);
   U15 : AOI22_X1 port map( A1 => D(11), A2 => n149, B1 => C(11), B2 => n145, 
                           ZN => n181);
   U16 : AOI22_X1 port map( A1 => D(12), A2 => n149, B1 => C(12), B2 => n145, 
                           ZN => n185);
   U17 : AOI22_X1 port map( A1 => D(13), A2 => n149, B1 => C(13), B2 => n145, 
                           ZN => n189);
   U18 : AOI22_X1 port map( A1 => D(14), A2 => n149, B1 => C(14), B2 => n145, 
                           ZN => n193);
   U19 : AOI22_X1 port map( A1 => D(15), A2 => n149, B1 => C(15), B2 => n145, 
                           ZN => n197);
   U20 : AOI22_X1 port map( A1 => D(16), A2 => n149, B1 => C(16), B2 => n145, 
                           ZN => n201);
   U21 : AOI22_X1 port map( A1 => D(17), A2 => n149, B1 => C(17), B2 => n145, 
                           ZN => n205);
   U22 : AOI22_X1 port map( A1 => D(18), A2 => n149, B1 => C(18), B2 => n145, 
                           ZN => n209);
   U23 : AOI22_X1 port map( A1 => D(19), A2 => n149, B1 => C(19), B2 => n145, 
                           ZN => n213);
   U24 : AOI22_X1 port map( A1 => D(20), A2 => n150, B1 => C(20), B2 => n146, 
                           ZN => n221);
   U25 : AOI22_X1 port map( A1 => D(21), A2 => n150, B1 => C(21), B2 => n146, 
                           ZN => n225);
   U26 : AOI22_X1 port map( A1 => D(22), A2 => n150, B1 => C(22), B2 => n146, 
                           ZN => n229);
   U27 : AOI22_X1 port map( A1 => D(23), A2 => n150, B1 => C(23), B2 => n146, 
                           ZN => n233);
   U28 : AOI22_X1 port map( A1 => D(24), A2 => n150, B1 => C(24), B2 => n146, 
                           ZN => n237);
   U29 : AOI22_X1 port map( A1 => D(25), A2 => n150, B1 => C(25), B2 => n146, 
                           ZN => n241);
   U30 : AOI22_X1 port map( A1 => D(26), A2 => n150, B1 => C(26), B2 => n146, 
                           ZN => n245);
   U31 : AOI22_X1 port map( A1 => D(27), A2 => n150, B1 => C(27), B2 => n146, 
                           ZN => n249);
   U32 : AOI22_X1 port map( A1 => D(28), A2 => n150, B1 => C(28), B2 => n146, 
                           ZN => n253);
   U33 : AOI22_X1 port map( A1 => D(29), A2 => n150, B1 => C(29), B2 => n146, 
                           ZN => n257);
   U34 : AOI22_X1 port map( A1 => D(30), A2 => n150, B1 => C(30), B2 => n146, 
                           ZN => n265);
   U35 : AOI22_X1 port map( A1 => D(31), A2 => n151, B1 => C(31), B2 => n147, 
                           ZN => n269);
   U36 : BUF_X1 port map( A => n152, Z => n149);
   U37 : BUF_X1 port map( A => n144, Z => n141);
   U38 : BUF_X1 port map( A => n152, Z => n150);
   U39 : BUF_X1 port map( A => n144, Z => n142);
   U40 : BUF_X1 port map( A => n153, Z => n154);
   U41 : BUF_X1 port map( A => n161, Z => n162);
   U42 : BUF_X1 port map( A => n153, Z => n155);
   U43 : BUF_X1 port map( A => n161, Z => n163);
   U44 : BUF_X1 port map( A => n152, Z => n151);
   U45 : BUF_X1 port map( A => n144, Z => n143);
   U46 : BUF_X1 port map( A => n153, Z => n156);
   U47 : BUF_X1 port map( A => n161, Z => n164);
   U48 : INV_X1 port map( A => S(1), ZN => n169);
   U49 : NOR3_X1 port map( A1 => n170, A2 => S(2), A3 => n169, ZN => n298);
   U50 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n170, ZN => n296);
   U51 : AND3_X1 port map( A1 => n170, A2 => n169, A3 => S(2), ZN => n299);
   U52 : AND3_X1 port map( A1 => S(1), A2 => n170, A3 => S(2), ZN => n301);
   U53 : BUF_X1 port map( A => n157, Z => n158);
   U54 : BUF_X1 port map( A => n165, Z => n166);
   U55 : BUF_X1 port map( A => n157, Z => n159);
   U56 : BUF_X1 port map( A => n165, Z => n167);
   U57 : BUF_X1 port map( A => n148, Z => n145);
   U58 : BUF_X1 port map( A => n140, Z => n1);
   U59 : BUF_X1 port map( A => n148, Z => n146);
   U60 : BUF_X1 port map( A => n140, Z => n2);
   U61 : BUF_X1 port map( A => n148, Z => n147);
   U62 : BUF_X1 port map( A => n140, Z => n139);
   U63 : BUF_X1 port map( A => n157, Z => n160);
   U64 : BUF_X1 port map( A => n165, Z => n168);
   U65 : INV_X1 port map( A => S(0), ZN => n170);
   U66 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n169, ZN => n297);
   U67 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => S(0), ZN => n295);
   U68 : AND3_X1 port map( A1 => S(0), A2 => n169, A3 => S(2), ZN => n300);
   U69 : AND3_X1 port map( A1 => S(1), A2 => S(0), A3 => S(2), ZN => n302);
   U70 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN 
                           => Y(5));
   U71 : AOI22_X1 port map( A1 => H(5), A2 => n168, B1 => G(5), B2 => n164, ZN 
                           => n279);
   U72 : AOI22_X1 port map( A1 => B(5), A2 => n143, B1 => A(5), B2 => n139, ZN 
                           => n282);
   U73 : AOI22_X1 port map( A1 => F(5), A2 => n160, B1 => E(5), B2 => n156, ZN 
                           => n280);
   U74 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN 
                           => Y(7));
   U75 : AOI22_X1 port map( A1 => H(7), A2 => n168, B1 => G(7), B2 => n164, ZN 
                           => n287);
   U76 : AOI22_X1 port map( A1 => B(7), A2 => n143, B1 => A(7), B2 => n139, ZN 
                           => n290);
   U77 : AOI22_X1 port map( A1 => F(7), A2 => n160, B1 => E(7), B2 => n156, ZN 
                           => n288);
   U78 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN 
                           => Y(9));
   U79 : AOI22_X1 port map( A1 => H(9), A2 => n168, B1 => G(9), B2 => n164, ZN 
                           => n303);
   U80 : AOI22_X1 port map( A1 => B(9), A2 => n143, B1 => A(9), B2 => n139, ZN 
                           => n306);
   U81 : AOI22_X1 port map( A1 => F(9), A2 => n160, B1 => E(9), B2 => n156, ZN 
                           => n304);
   U82 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(11));
   U83 : AOI22_X1 port map( A1 => H(11), A2 => n166, B1 => G(11), B2 => n162, 
                           ZN => n179);
   U84 : AOI22_X1 port map( A1 => B(11), A2 => n141, B1 => A(11), B2 => n1, ZN 
                           => n182);
   U85 : AOI22_X1 port map( A1 => F(11), A2 => n158, B1 => E(11), B2 => n154, 
                           ZN => n180);
   U86 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(13));
   U87 : AOI22_X1 port map( A1 => H(13), A2 => n166, B1 => G(13), B2 => n162, 
                           ZN => n187);
   U88 : AOI22_X1 port map( A1 => B(13), A2 => n141, B1 => A(13), B2 => n1, ZN 
                           => n190);
   U89 : AOI22_X1 port map( A1 => F(13), A2 => n158, B1 => E(13), B2 => n154, 
                           ZN => n188);
   U90 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(15));
   U91 : AOI22_X1 port map( A1 => H(15), A2 => n166, B1 => G(15), B2 => n162, 
                           ZN => n195);
   U92 : AOI22_X1 port map( A1 => B(15), A2 => n141, B1 => A(15), B2 => n1, ZN 
                           => n198);
   U93 : AOI22_X1 port map( A1 => F(15), A2 => n158, B1 => E(15), B2 => n154, 
                           ZN => n196);
   U94 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(17));
   U95 : AOI22_X1 port map( A1 => H(17), A2 => n166, B1 => G(17), B2 => n162, 
                           ZN => n203);
   U96 : AOI22_X1 port map( A1 => B(17), A2 => n141, B1 => A(17), B2 => n1, ZN 
                           => n206);
   U97 : AOI22_X1 port map( A1 => F(17), A2 => n158, B1 => E(17), B2 => n154, 
                           ZN => n204);
   U98 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(19));
   U99 : AOI22_X1 port map( A1 => H(19), A2 => n166, B1 => G(19), B2 => n162, 
                           ZN => n211);
   U100 : AOI22_X1 port map( A1 => B(19), A2 => n141, B1 => A(19), B2 => n1, ZN
                           => n214);
   U101 : AOI22_X1 port map( A1 => F(19), A2 => n158, B1 => E(19), B2 => n154, 
                           ZN => n212);
   U102 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(21));
   U103 : AOI22_X1 port map( A1 => H(21), A2 => n167, B1 => G(21), B2 => n163, 
                           ZN => n223);
   U104 : AOI22_X1 port map( A1 => B(21), A2 => n142, B1 => A(21), B2 => n2, ZN
                           => n226);
   U105 : AOI22_X1 port map( A1 => F(21), A2 => n159, B1 => E(21), B2 => n155, 
                           ZN => n224);
   U106 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(23));
   U107 : AOI22_X1 port map( A1 => H(23), A2 => n167, B1 => G(23), B2 => n163, 
                           ZN => n231);
   U108 : AOI22_X1 port map( A1 => B(23), A2 => n142, B1 => A(23), B2 => n2, ZN
                           => n234);
   U109 : AOI22_X1 port map( A1 => F(23), A2 => n159, B1 => E(23), B2 => n155, 
                           ZN => n232);
   U110 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(25));
   U111 : AOI22_X1 port map( A1 => H(25), A2 => n167, B1 => G(25), B2 => n163, 
                           ZN => n239);
   U112 : AOI22_X1 port map( A1 => B(25), A2 => n142, B1 => A(25), B2 => n2, ZN
                           => n242);
   U113 : AOI22_X1 port map( A1 => F(25), A2 => n159, B1 => E(25), B2 => n155, 
                           ZN => n240);
   U114 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(27));
   U115 : AOI22_X1 port map( A1 => H(27), A2 => n167, B1 => G(27), B2 => n163, 
                           ZN => n247);
   U116 : AOI22_X1 port map( A1 => B(27), A2 => n142, B1 => A(27), B2 => n2, ZN
                           => n250);
   U117 : AOI22_X1 port map( A1 => F(27), A2 => n159, B1 => E(27), B2 => n155, 
                           ZN => n248);
   U118 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(30));
   U119 : AOI22_X1 port map( A1 => H(30), A2 => n167, B1 => G(30), B2 => n163, 
                           ZN => n263);
   U120 : AOI22_X1 port map( A1 => B(30), A2 => n142, B1 => A(30), B2 => n2, ZN
                           => n266);
   U121 : AOI22_X1 port map( A1 => F(30), A2 => n159, B1 => E(30), B2 => n155, 
                           ZN => n264);
   U122 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(6));
   U123 : AOI22_X1 port map( A1 => H(6), A2 => n168, B1 => G(6), B2 => n164, ZN
                           => n283);
   U124 : AOI22_X1 port map( A1 => B(6), A2 => n143, B1 => A(6), B2 => n139, ZN
                           => n286);
   U125 : AOI22_X1 port map( A1 => F(6), A2 => n160, B1 => E(6), B2 => n156, ZN
                           => n284);
   U126 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(8));
   U127 : AOI22_X1 port map( A1 => H(8), A2 => n168, B1 => G(8), B2 => n164, ZN
                           => n291);
   U128 : AOI22_X1 port map( A1 => B(8), A2 => n143, B1 => A(8), B2 => n139, ZN
                           => n294);
   U129 : AOI22_X1 port map( A1 => F(8), A2 => n160, B1 => E(8), B2 => n156, ZN
                           => n292);
   U130 : NAND4_X1 port map( A1 => n178, A2 => n177, A3 => n176, A4 => n175, ZN
                           => Y(10));
   U131 : AOI22_X1 port map( A1 => H(10), A2 => n166, B1 => G(10), B2 => n162, 
                           ZN => n175);
   U132 : AOI22_X1 port map( A1 => B(10), A2 => n141, B1 => A(10), B2 => n1, ZN
                           => n178);
   U133 : AOI22_X1 port map( A1 => F(10), A2 => n158, B1 => E(10), B2 => n154, 
                           ZN => n176);
   U134 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN
                           => Y(12));
   U135 : AOI22_X1 port map( A1 => H(12), A2 => n166, B1 => G(12), B2 => n162, 
                           ZN => n183);
   U136 : AOI22_X1 port map( A1 => B(12), A2 => n141, B1 => A(12), B2 => n1, ZN
                           => n186);
   U137 : AOI22_X1 port map( A1 => F(12), A2 => n158, B1 => E(12), B2 => n154, 
                           ZN => n184);
   U138 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN
                           => Y(14));
   U139 : AOI22_X1 port map( A1 => H(14), A2 => n166, B1 => G(14), B2 => n162, 
                           ZN => n191);
   U140 : AOI22_X1 port map( A1 => B(14), A2 => n141, B1 => A(14), B2 => n1, ZN
                           => n194);
   U141 : AOI22_X1 port map( A1 => F(14), A2 => n158, B1 => E(14), B2 => n154, 
                           ZN => n192);
   U142 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN
                           => Y(16));
   U143 : AOI22_X1 port map( A1 => H(16), A2 => n166, B1 => G(16), B2 => n162, 
                           ZN => n199);
   U144 : AOI22_X1 port map( A1 => B(16), A2 => n141, B1 => A(16), B2 => n1, ZN
                           => n202);
   U145 : AOI22_X1 port map( A1 => F(16), A2 => n158, B1 => E(16), B2 => n154, 
                           ZN => n200);
   U146 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN
                           => Y(18));
   U147 : AOI22_X1 port map( A1 => H(18), A2 => n166, B1 => G(18), B2 => n162, 
                           ZN => n207);
   U148 : AOI22_X1 port map( A1 => B(18), A2 => n141, B1 => A(18), B2 => n1, ZN
                           => n210);
   U149 : AOI22_X1 port map( A1 => F(18), A2 => n158, B1 => E(18), B2 => n154, 
                           ZN => n208);
   U150 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(20));
   U151 : AOI22_X1 port map( A1 => H(20), A2 => n167, B1 => G(20), B2 => n163, 
                           ZN => n219);
   U152 : AOI22_X1 port map( A1 => B(20), A2 => n142, B1 => A(20), B2 => n2, ZN
                           => n222);
   U153 : AOI22_X1 port map( A1 => F(20), A2 => n159, B1 => E(20), B2 => n155, 
                           ZN => n220);
   U154 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(22));
   U155 : AOI22_X1 port map( A1 => H(22), A2 => n167, B1 => G(22), B2 => n163, 
                           ZN => n227);
   U156 : AOI22_X1 port map( A1 => B(22), A2 => n142, B1 => A(22), B2 => n2, ZN
                           => n230);
   U157 : AOI22_X1 port map( A1 => F(22), A2 => n159, B1 => E(22), B2 => n155, 
                           ZN => n228);
   U158 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(24));
   U159 : AOI22_X1 port map( A1 => H(24), A2 => n167, B1 => G(24), B2 => n163, 
                           ZN => n235);
   U160 : AOI22_X1 port map( A1 => B(24), A2 => n142, B1 => A(24), B2 => n2, ZN
                           => n238);
   U161 : AOI22_X1 port map( A1 => F(24), A2 => n159, B1 => E(24), B2 => n155, 
                           ZN => n236);
   U162 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(26));
   U163 : AOI22_X1 port map( A1 => H(26), A2 => n167, B1 => G(26), B2 => n163, 
                           ZN => n243);
   U164 : AOI22_X1 port map( A1 => B(26), A2 => n142, B1 => A(26), B2 => n2, ZN
                           => n246);
   U165 : AOI22_X1 port map( A1 => F(26), A2 => n159, B1 => E(26), B2 => n155, 
                           ZN => n244);
   U166 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(28));
   U167 : AOI22_X1 port map( A1 => H(28), A2 => n167, B1 => G(28), B2 => n163, 
                           ZN => n251);
   U168 : AOI22_X1 port map( A1 => B(28), A2 => n142, B1 => A(28), B2 => n2, ZN
                           => n254);
   U169 : AOI22_X1 port map( A1 => F(28), A2 => n159, B1 => E(28), B2 => n155, 
                           ZN => n252);
   U170 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(31));
   U171 : AOI22_X1 port map( A1 => H(31), A2 => n168, B1 => G(31), B2 => n164, 
                           ZN => n267);
   U172 : AOI22_X1 port map( A1 => B(31), A2 => n143, B1 => A(31), B2 => n139, 
                           ZN => n270);
   U173 : AOI22_X1 port map( A1 => F(31), A2 => n160, B1 => E(31), B2 => n156, 
                           ZN => n268);
   U174 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(4));
   U175 : AOI22_X1 port map( A1 => F(4), A2 => n160, B1 => E(4), B2 => n156, ZN
                           => n276);
   U176 : AOI22_X1 port map( A1 => H(4), A2 => n168, B1 => G(4), B2 => n164, ZN
                           => n275);
   U177 : AOI22_X1 port map( A1 => B(4), A2 => n143, B1 => A(4), B2 => n139, ZN
                           => n278);
   U178 : NAND4_X1 port map( A1 => n174, A2 => n173, A3 => n172, A4 => n171, ZN
                           => Y(0));
   U179 : AOI22_X1 port map( A1 => B(0), A2 => n141, B1 => A(0), B2 => n1, ZN 
                           => n174);
   U180 : AOI22_X1 port map( A1 => D(0), A2 => n149, B1 => C(0), B2 => n145, ZN
                           => n173);
   U181 : AOI22_X1 port map( A1 => F(0), A2 => n158, B1 => E(0), B2 => n154, ZN
                           => n172);
   U182 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN
                           => Y(1));
   U183 : AOI22_X1 port map( A1 => B(1), A2 => n141, B1 => A(1), B2 => n1, ZN 
                           => n218);
   U184 : AOI22_X1 port map( A1 => D(1), A2 => n149, B1 => C(1), B2 => n145, ZN
                           => n217);
   U185 : AOI22_X1 port map( A1 => F(1), A2 => n158, B1 => E(1), B2 => n154, ZN
                           => n216);
   U186 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(2));
   U187 : AOI22_X1 port map( A1 => B(2), A2 => n142, B1 => A(2), B2 => n2, ZN 
                           => n262);
   U188 : AOI22_X1 port map( A1 => D(2), A2 => n150, B1 => C(2), B2 => n146, ZN
                           => n261);
   U189 : AOI22_X1 port map( A1 => F(2), A2 => n159, B1 => E(2), B2 => n155, ZN
                           => n260);
   U190 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(3));
   U191 : AOI22_X1 port map( A1 => B(3), A2 => n143, B1 => A(3), B2 => n139, ZN
                           => n274);
   U192 : AOI22_X1 port map( A1 => D(3), A2 => n151, B1 => C(3), B2 => n147, ZN
                           => n273);
   U193 : AOI22_X1 port map( A1 => F(3), A2 => n160, B1 => E(3), B2 => n156, ZN
                           => n272);
   U194 : AOI22_X1 port map( A1 => D(4), A2 => n151, B1 => C(4), B2 => n147, ZN
                           => n277);
   U195 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(29));
   U196 : AOI22_X1 port map( A1 => H(29), A2 => n167, B1 => G(29), B2 => n163, 
                           ZN => n255);
   U197 : AOI22_X1 port map( A1 => B(29), A2 => n142, B1 => A(29), B2 => n2, ZN
                           => n258);
   U198 : AOI22_X1 port map( A1 => F(29), A2 => n159, B1 => E(29), B2 => n155, 
                           ZN => n256);
   U199 : AOI22_X1 port map( A1 => H(0), A2 => n166, B1 => G(0), B2 => n162, ZN
                           => n171);
   U200 : AOI22_X1 port map( A1 => H(1), A2 => n166, B1 => G(1), B2 => n162, ZN
                           => n215);
   U201 : AOI22_X1 port map( A1 => H(2), A2 => n167, B1 => G(2), B2 => n163, ZN
                           => n259);
   U202 : AOI22_X1 port map( A1 => H(3), A2 => n168, B1 => G(3), B2 => n164, ZN
                           => n271);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX81_N32_0 is

   port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX81_N32_0;

architecture SYN_BEHAVIORAL of MUX81_N32_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n296, Z => n144);
   U2 : BUF_X1 port map( A => n298, Z => n152);
   U3 : BUF_X1 port map( A => n299, Z => n153);
   U4 : BUF_X1 port map( A => n301, Z => n161);
   U5 : BUF_X1 port map( A => n297, Z => n148);
   U6 : BUF_X1 port map( A => n295, Z => n140);
   U7 : BUF_X1 port map( A => n300, Z => n157);
   U8 : BUF_X1 port map( A => n302, Z => n165);
   U9 : AOI22_X1 port map( A1 => D(7), A2 => n151, B1 => C(7), B2 => n147, ZN 
                           => n289);
   U10 : AOI22_X1 port map( A1 => D(8), A2 => n151, B1 => C(8), B2 => n147, ZN 
                           => n293);
   U11 : AOI22_X1 port map( A1 => D(9), A2 => n151, B1 => C(9), B2 => n147, ZN 
                           => n305);
   U12 : AOI22_X1 port map( A1 => D(10), A2 => n149, B1 => C(10), B2 => n145, 
                           ZN => n177);
   U13 : AOI22_X1 port map( A1 => D(11), A2 => n149, B1 => C(11), B2 => n145, 
                           ZN => n181);
   U14 : AOI22_X1 port map( A1 => D(12), A2 => n149, B1 => C(12), B2 => n145, 
                           ZN => n185);
   U15 : AOI22_X1 port map( A1 => D(13), A2 => n149, B1 => C(13), B2 => n145, 
                           ZN => n189);
   U16 : AOI22_X1 port map( A1 => D(14), A2 => n149, B1 => C(14), B2 => n145, 
                           ZN => n193);
   U17 : AOI22_X1 port map( A1 => D(15), A2 => n149, B1 => C(15), B2 => n145, 
                           ZN => n197);
   U18 : AOI22_X1 port map( A1 => D(16), A2 => n149, B1 => C(16), B2 => n145, 
                           ZN => n201);
   U19 : AOI22_X1 port map( A1 => D(17), A2 => n149, B1 => C(17), B2 => n145, 
                           ZN => n205);
   U20 : AOI22_X1 port map( A1 => D(18), A2 => n149, B1 => C(18), B2 => n145, 
                           ZN => n209);
   U21 : AOI22_X1 port map( A1 => D(19), A2 => n149, B1 => C(19), B2 => n145, 
                           ZN => n213);
   U22 : AOI22_X1 port map( A1 => D(20), A2 => n150, B1 => C(20), B2 => n146, 
                           ZN => n221);
   U23 : AOI22_X1 port map( A1 => D(21), A2 => n150, B1 => C(21), B2 => n146, 
                           ZN => n225);
   U24 : AOI22_X1 port map( A1 => D(22), A2 => n150, B1 => C(22), B2 => n146, 
                           ZN => n229);
   U25 : AOI22_X1 port map( A1 => D(23), A2 => n150, B1 => C(23), B2 => n146, 
                           ZN => n233);
   U26 : AOI22_X1 port map( A1 => D(24), A2 => n150, B1 => C(24), B2 => n146, 
                           ZN => n237);
   U27 : AOI22_X1 port map( A1 => D(25), A2 => n150, B1 => C(25), B2 => n146, 
                           ZN => n241);
   U28 : AOI22_X1 port map( A1 => D(26), A2 => n150, B1 => C(26), B2 => n146, 
                           ZN => n245);
   U29 : AOI22_X1 port map( A1 => D(27), A2 => n150, B1 => C(27), B2 => n146, 
                           ZN => n249);
   U30 : AOI22_X1 port map( A1 => D(28), A2 => n150, B1 => C(28), B2 => n146, 
                           ZN => n253);
   U31 : AOI22_X1 port map( A1 => D(29), A2 => n150, B1 => C(29), B2 => n146, 
                           ZN => n257);
   U32 : AOI22_X1 port map( A1 => D(30), A2 => n150, B1 => C(30), B2 => n146, 
                           ZN => n265);
   U33 : AOI22_X1 port map( A1 => D(31), A2 => n151, B1 => C(31), B2 => n147, 
                           ZN => n269);
   U34 : BUF_X1 port map( A => n152, Z => n149);
   U35 : BUF_X1 port map( A => n144, Z => n141);
   U36 : BUF_X1 port map( A => n152, Z => n150);
   U37 : BUF_X1 port map( A => n144, Z => n142);
   U38 : BUF_X1 port map( A => n153, Z => n154);
   U39 : BUF_X1 port map( A => n161, Z => n162);
   U40 : BUF_X1 port map( A => n153, Z => n155);
   U41 : BUF_X1 port map( A => n161, Z => n163);
   U42 : BUF_X1 port map( A => n152, Z => n151);
   U43 : BUF_X1 port map( A => n144, Z => n143);
   U44 : BUF_X1 port map( A => n153, Z => n156);
   U45 : BUF_X1 port map( A => n161, Z => n164);
   U46 : INV_X1 port map( A => S(1), ZN => n169);
   U47 : NOR3_X1 port map( A1 => n170, A2 => S(2), A3 => n169, ZN => n298);
   U48 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n170, ZN => n296);
   U49 : AND3_X1 port map( A1 => n170, A2 => n169, A3 => S(2), ZN => n299);
   U50 : AND3_X1 port map( A1 => S(1), A2 => n170, A3 => S(2), ZN => n301);
   U51 : BUF_X1 port map( A => n157, Z => n158);
   U52 : BUF_X1 port map( A => n165, Z => n166);
   U53 : BUF_X1 port map( A => n157, Z => n159);
   U54 : BUF_X1 port map( A => n165, Z => n167);
   U55 : BUF_X1 port map( A => n148, Z => n145);
   U56 : BUF_X1 port map( A => n140, Z => n1);
   U57 : BUF_X1 port map( A => n148, Z => n146);
   U58 : BUF_X1 port map( A => n140, Z => n2);
   U59 : BUF_X1 port map( A => n148, Z => n147);
   U60 : BUF_X1 port map( A => n140, Z => n139);
   U61 : BUF_X1 port map( A => n157, Z => n160);
   U62 : BUF_X1 port map( A => n165, Z => n168);
   U63 : INV_X1 port map( A => S(0), ZN => n170);
   U64 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n169, ZN => n297);
   U65 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => S(0), ZN => n295);
   U66 : AND3_X1 port map( A1 => S(0), A2 => n169, A3 => S(2), ZN => n300);
   U67 : AND3_X1 port map( A1 => S(1), A2 => S(0), A3 => S(2), ZN => n302);
   U68 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN 
                           => Y(7));
   U69 : AOI22_X1 port map( A1 => H(7), A2 => n168, B1 => G(7), B2 => n164, ZN 
                           => n287);
   U70 : AOI22_X1 port map( A1 => B(7), A2 => n143, B1 => A(7), B2 => n139, ZN 
                           => n290);
   U71 : AOI22_X1 port map( A1 => F(7), A2 => n160, B1 => E(7), B2 => n156, ZN 
                           => n288);
   U72 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN 
                           => Y(9));
   U73 : AOI22_X1 port map( A1 => H(9), A2 => n168, B1 => G(9), B2 => n164, ZN 
                           => n303);
   U74 : AOI22_X1 port map( A1 => B(9), A2 => n143, B1 => A(9), B2 => n139, ZN 
                           => n306);
   U75 : AOI22_X1 port map( A1 => F(9), A2 => n160, B1 => E(9), B2 => n156, ZN 
                           => n304);
   U76 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(11));
   U77 : AOI22_X1 port map( A1 => H(11), A2 => n166, B1 => G(11), B2 => n162, 
                           ZN => n179);
   U78 : AOI22_X1 port map( A1 => B(11), A2 => n141, B1 => A(11), B2 => n1, ZN 
                           => n182);
   U79 : AOI22_X1 port map( A1 => F(11), A2 => n158, B1 => E(11), B2 => n154, 
                           ZN => n180);
   U80 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(13));
   U81 : AOI22_X1 port map( A1 => H(13), A2 => n166, B1 => G(13), B2 => n162, 
                           ZN => n187);
   U82 : AOI22_X1 port map( A1 => B(13), A2 => n141, B1 => A(13), B2 => n1, ZN 
                           => n190);
   U83 : AOI22_X1 port map( A1 => F(13), A2 => n158, B1 => E(13), B2 => n154, 
                           ZN => n188);
   U84 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(15));
   U85 : AOI22_X1 port map( A1 => H(15), A2 => n166, B1 => G(15), B2 => n162, 
                           ZN => n195);
   U86 : AOI22_X1 port map( A1 => B(15), A2 => n141, B1 => A(15), B2 => n1, ZN 
                           => n198);
   U87 : AOI22_X1 port map( A1 => F(15), A2 => n158, B1 => E(15), B2 => n154, 
                           ZN => n196);
   U88 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(17));
   U89 : AOI22_X1 port map( A1 => H(17), A2 => n166, B1 => G(17), B2 => n162, 
                           ZN => n203);
   U90 : AOI22_X1 port map( A1 => B(17), A2 => n141, B1 => A(17), B2 => n1, ZN 
                           => n206);
   U91 : AOI22_X1 port map( A1 => F(17), A2 => n158, B1 => E(17), B2 => n154, 
                           ZN => n204);
   U92 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(19));
   U93 : AOI22_X1 port map( A1 => H(19), A2 => n166, B1 => G(19), B2 => n162, 
                           ZN => n211);
   U94 : AOI22_X1 port map( A1 => B(19), A2 => n141, B1 => A(19), B2 => n1, ZN 
                           => n214);
   U95 : AOI22_X1 port map( A1 => F(19), A2 => n158, B1 => E(19), B2 => n154, 
                           ZN => n212);
   U96 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN 
                           => Y(21));
   U97 : AOI22_X1 port map( A1 => H(21), A2 => n167, B1 => G(21), B2 => n163, 
                           ZN => n223);
   U98 : AOI22_X1 port map( A1 => B(21), A2 => n142, B1 => A(21), B2 => n2, ZN 
                           => n226);
   U99 : AOI22_X1 port map( A1 => F(21), A2 => n159, B1 => E(21), B2 => n155, 
                           ZN => n224);
   U100 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(23));
   U101 : AOI22_X1 port map( A1 => H(23), A2 => n167, B1 => G(23), B2 => n163, 
                           ZN => n231);
   U102 : AOI22_X1 port map( A1 => B(23), A2 => n142, B1 => A(23), B2 => n2, ZN
                           => n234);
   U103 : AOI22_X1 port map( A1 => F(23), A2 => n159, B1 => E(23), B2 => n155, 
                           ZN => n232);
   U104 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(25));
   U105 : AOI22_X1 port map( A1 => H(25), A2 => n167, B1 => G(25), B2 => n163, 
                           ZN => n239);
   U106 : AOI22_X1 port map( A1 => B(25), A2 => n142, B1 => A(25), B2 => n2, ZN
                           => n242);
   U107 : AOI22_X1 port map( A1 => F(25), A2 => n159, B1 => E(25), B2 => n155, 
                           ZN => n240);
   U108 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(27));
   U109 : AOI22_X1 port map( A1 => H(27), A2 => n167, B1 => G(27), B2 => n163, 
                           ZN => n247);
   U110 : AOI22_X1 port map( A1 => B(27), A2 => n142, B1 => A(27), B2 => n2, ZN
                           => n250);
   U111 : AOI22_X1 port map( A1 => F(27), A2 => n159, B1 => E(27), B2 => n155, 
                           ZN => n248);
   U112 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(30));
   U113 : AOI22_X1 port map( A1 => H(30), A2 => n167, B1 => G(30), B2 => n163, 
                           ZN => n263);
   U114 : AOI22_X1 port map( A1 => B(30), A2 => n142, B1 => A(30), B2 => n2, ZN
                           => n266);
   U115 : AOI22_X1 port map( A1 => F(30), A2 => n159, B1 => E(30), B2 => n155, 
                           ZN => n264);
   U116 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(8));
   U117 : AOI22_X1 port map( A1 => H(8), A2 => n168, B1 => G(8), B2 => n164, ZN
                           => n291);
   U118 : AOI22_X1 port map( A1 => B(8), A2 => n143, B1 => A(8), B2 => n139, ZN
                           => n294);
   U119 : AOI22_X1 port map( A1 => F(8), A2 => n160, B1 => E(8), B2 => n156, ZN
                           => n292);
   U120 : NAND4_X1 port map( A1 => n178, A2 => n177, A3 => n176, A4 => n175, ZN
                           => Y(10));
   U121 : AOI22_X1 port map( A1 => H(10), A2 => n166, B1 => G(10), B2 => n162, 
                           ZN => n175);
   U122 : AOI22_X1 port map( A1 => B(10), A2 => n141, B1 => A(10), B2 => n1, ZN
                           => n178);
   U123 : AOI22_X1 port map( A1 => F(10), A2 => n158, B1 => E(10), B2 => n154, 
                           ZN => n176);
   U124 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN
                           => Y(12));
   U125 : AOI22_X1 port map( A1 => H(12), A2 => n166, B1 => G(12), B2 => n162, 
                           ZN => n183);
   U126 : AOI22_X1 port map( A1 => B(12), A2 => n141, B1 => A(12), B2 => n1, ZN
                           => n186);
   U127 : AOI22_X1 port map( A1 => F(12), A2 => n158, B1 => E(12), B2 => n154, 
                           ZN => n184);
   U128 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN
                           => Y(14));
   U129 : AOI22_X1 port map( A1 => H(14), A2 => n166, B1 => G(14), B2 => n162, 
                           ZN => n191);
   U130 : AOI22_X1 port map( A1 => B(14), A2 => n141, B1 => A(14), B2 => n1, ZN
                           => n194);
   U131 : AOI22_X1 port map( A1 => F(14), A2 => n158, B1 => E(14), B2 => n154, 
                           ZN => n192);
   U132 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN
                           => Y(16));
   U133 : AOI22_X1 port map( A1 => H(16), A2 => n166, B1 => G(16), B2 => n162, 
                           ZN => n199);
   U134 : AOI22_X1 port map( A1 => B(16), A2 => n141, B1 => A(16), B2 => n1, ZN
                           => n202);
   U135 : AOI22_X1 port map( A1 => F(16), A2 => n158, B1 => E(16), B2 => n154, 
                           ZN => n200);
   U136 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN
                           => Y(18));
   U137 : AOI22_X1 port map( A1 => H(18), A2 => n166, B1 => G(18), B2 => n162, 
                           ZN => n207);
   U138 : AOI22_X1 port map( A1 => B(18), A2 => n141, B1 => A(18), B2 => n1, ZN
                           => n210);
   U139 : AOI22_X1 port map( A1 => F(18), A2 => n158, B1 => E(18), B2 => n154, 
                           ZN => n208);
   U140 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(20));
   U141 : AOI22_X1 port map( A1 => H(20), A2 => n167, B1 => G(20), B2 => n163, 
                           ZN => n219);
   U142 : AOI22_X1 port map( A1 => B(20), A2 => n142, B1 => A(20), B2 => n2, ZN
                           => n222);
   U143 : AOI22_X1 port map( A1 => F(20), A2 => n159, B1 => E(20), B2 => n155, 
                           ZN => n220);
   U144 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(22));
   U145 : AOI22_X1 port map( A1 => H(22), A2 => n167, B1 => G(22), B2 => n163, 
                           ZN => n227);
   U146 : AOI22_X1 port map( A1 => B(22), A2 => n142, B1 => A(22), B2 => n2, ZN
                           => n230);
   U147 : AOI22_X1 port map( A1 => F(22), A2 => n159, B1 => E(22), B2 => n155, 
                           ZN => n228);
   U148 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(24));
   U149 : AOI22_X1 port map( A1 => H(24), A2 => n167, B1 => G(24), B2 => n163, 
                           ZN => n235);
   U150 : AOI22_X1 port map( A1 => B(24), A2 => n142, B1 => A(24), B2 => n2, ZN
                           => n238);
   U151 : AOI22_X1 port map( A1 => F(24), A2 => n159, B1 => E(24), B2 => n155, 
                           ZN => n236);
   U152 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(26));
   U153 : AOI22_X1 port map( A1 => H(26), A2 => n167, B1 => G(26), B2 => n163, 
                           ZN => n243);
   U154 : AOI22_X1 port map( A1 => B(26), A2 => n142, B1 => A(26), B2 => n2, ZN
                           => n246);
   U155 : AOI22_X1 port map( A1 => F(26), A2 => n159, B1 => E(26), B2 => n155, 
                           ZN => n244);
   U156 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(28));
   U157 : AOI22_X1 port map( A1 => H(28), A2 => n167, B1 => G(28), B2 => n163, 
                           ZN => n251);
   U158 : AOI22_X1 port map( A1 => B(28), A2 => n142, B1 => A(28), B2 => n2, ZN
                           => n254);
   U159 : AOI22_X1 port map( A1 => F(28), A2 => n159, B1 => E(28), B2 => n155, 
                           ZN => n252);
   U160 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(31));
   U161 : AOI22_X1 port map( A1 => H(31), A2 => n168, B1 => G(31), B2 => n164, 
                           ZN => n267);
   U162 : AOI22_X1 port map( A1 => B(31), A2 => n143, B1 => A(31), B2 => n139, 
                           ZN => n270);
   U163 : AOI22_X1 port map( A1 => F(31), A2 => n160, B1 => E(31), B2 => n156, 
                           ZN => n268);
   U164 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(6));
   U165 : AOI22_X1 port map( A1 => F(6), A2 => n160, B1 => E(6), B2 => n156, ZN
                           => n284);
   U166 : AOI22_X1 port map( A1 => H(6), A2 => n168, B1 => G(6), B2 => n164, ZN
                           => n283);
   U167 : AOI22_X1 port map( A1 => B(6), A2 => n143, B1 => A(6), B2 => n139, ZN
                           => n286);
   U168 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(5));
   U169 : AOI22_X1 port map( A1 => B(5), A2 => n143, B1 => A(5), B2 => n139, ZN
                           => n282);
   U170 : AOI22_X1 port map( A1 => D(5), A2 => n151, B1 => C(5), B2 => n147, ZN
                           => n281);
   U171 : AOI22_X1 port map( A1 => F(5), A2 => n160, B1 => E(5), B2 => n156, ZN
                           => n280);
   U172 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(4));
   U173 : AOI22_X1 port map( A1 => B(4), A2 => n143, B1 => A(4), B2 => n139, ZN
                           => n278);
   U174 : AOI22_X1 port map( A1 => D(4), A2 => n151, B1 => C(4), B2 => n147, ZN
                           => n277);
   U175 : AOI22_X1 port map( A1 => F(4), A2 => n160, B1 => E(4), B2 => n156, ZN
                           => n276);
   U176 : NAND4_X1 port map( A1 => n174, A2 => n173, A3 => n172, A4 => n171, ZN
                           => Y(0));
   U177 : AOI22_X1 port map( A1 => B(0), A2 => n141, B1 => A(0), B2 => n1, ZN 
                           => n174);
   U178 : AOI22_X1 port map( A1 => D(0), A2 => n149, B1 => C(0), B2 => n145, ZN
                           => n173);
   U179 : AOI22_X1 port map( A1 => F(0), A2 => n158, B1 => E(0), B2 => n154, ZN
                           => n172);
   U180 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN
                           => Y(1));
   U181 : AOI22_X1 port map( A1 => B(1), A2 => n141, B1 => A(1), B2 => n1, ZN 
                           => n218);
   U182 : AOI22_X1 port map( A1 => D(1), A2 => n149, B1 => C(1), B2 => n145, ZN
                           => n217);
   U183 : AOI22_X1 port map( A1 => F(1), A2 => n158, B1 => E(1), B2 => n154, ZN
                           => n216);
   U184 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(2));
   U185 : AOI22_X1 port map( A1 => B(2), A2 => n142, B1 => A(2), B2 => n2, ZN 
                           => n262);
   U186 : AOI22_X1 port map( A1 => D(2), A2 => n150, B1 => C(2), B2 => n146, ZN
                           => n261);
   U187 : AOI22_X1 port map( A1 => F(2), A2 => n159, B1 => E(2), B2 => n155, ZN
                           => n260);
   U188 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(3));
   U189 : AOI22_X1 port map( A1 => B(3), A2 => n143, B1 => A(3), B2 => n139, ZN
                           => n274);
   U190 : AOI22_X1 port map( A1 => D(3), A2 => n151, B1 => C(3), B2 => n147, ZN
                           => n273);
   U191 : AOI22_X1 port map( A1 => F(3), A2 => n160, B1 => E(3), B2 => n156, ZN
                           => n272);
   U192 : AOI22_X1 port map( A1 => D(6), A2 => n151, B1 => C(6), B2 => n147, ZN
                           => n285);
   U193 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(29));
   U194 : AOI22_X1 port map( A1 => H(29), A2 => n167, B1 => G(29), B2 => n163, 
                           ZN => n255);
   U195 : AOI22_X1 port map( A1 => B(29), A2 => n142, B1 => A(29), B2 => n2, ZN
                           => n258);
   U196 : AOI22_X1 port map( A1 => F(29), A2 => n159, B1 => E(29), B2 => n155, 
                           ZN => n256);
   U197 : AOI22_X1 port map( A1 => H(0), A2 => n166, B1 => G(0), B2 => n162, ZN
                           => n171);
   U198 : AOI22_X1 port map( A1 => H(1), A2 => n166, B1 => G(1), B2 => n162, ZN
                           => n215);
   U199 : AOI22_X1 port map( A1 => H(2), A2 => n167, B1 => G(2), B2 => n163, ZN
                           => n259);
   U200 : AOI22_X1 port map( A1 => H(3), A2 => n168, B1 => G(3), B2 => n164, ZN
                           => n271);
   U201 : AOI22_X1 port map( A1 => H(4), A2 => n168, B1 => G(4), B2 => n164, ZN
                           => n275);
   U202 : AOI22_X1 port map( A1 => H(5), A2 => n168, B1 => G(5), B2 => n164, ZN
                           => n279);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_60;

architecture SYN_BEHAVIORAL of AND2_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_59;

architecture SYN_BEHAVIORAL of AND2_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_58;

architecture SYN_BEHAVIORAL of AND2_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_57;

architecture SYN_BEHAVIORAL of AND2_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_56;

architecture SYN_BEHAVIORAL of AND2_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_55;

architecture SYN_BEHAVIORAL of AND2_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_54;

architecture SYN_BEHAVIORAL of AND2_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_53;

architecture SYN_BEHAVIORAL of AND2_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_52;

architecture SYN_BEHAVIORAL of AND2_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_51;

architecture SYN_BEHAVIORAL of AND2_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_50;

architecture SYN_BEHAVIORAL of AND2_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_49;

architecture SYN_BEHAVIORAL of AND2_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_48;

architecture SYN_BEHAVIORAL of AND2_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_47;

architecture SYN_BEHAVIORAL of AND2_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_46;

architecture SYN_BEHAVIORAL of AND2_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_45;

architecture SYN_BEHAVIORAL of AND2_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_44;

architecture SYN_BEHAVIORAL of AND2_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_43;

architecture SYN_BEHAVIORAL of AND2_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_42;

architecture SYN_BEHAVIORAL of AND2_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_41;

architecture SYN_BEHAVIORAL of AND2_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_40;

architecture SYN_BEHAVIORAL of AND2_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_39;

architecture SYN_BEHAVIORAL of AND2_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_38;

architecture SYN_BEHAVIORAL of AND2_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_37;

architecture SYN_BEHAVIORAL of AND2_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_36;

architecture SYN_BEHAVIORAL of AND2_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_35;

architecture SYN_BEHAVIORAL of AND2_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_34;

architecture SYN_BEHAVIORAL of AND2_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_33;

architecture SYN_BEHAVIORAL of AND2_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_32;

architecture SYN_BEHAVIORAL of AND2_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_31;

architecture SYN_BEHAVIORAL of AND2_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_30;

architecture SYN_BEHAVIORAL of AND2_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_29;

architecture SYN_BEHAVIORAL of AND2_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_28;

architecture SYN_BEHAVIORAL of AND2_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_27;

architecture SYN_BEHAVIORAL of AND2_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_26;

architecture SYN_BEHAVIORAL of AND2_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_25;

architecture SYN_BEHAVIORAL of AND2_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_24;

architecture SYN_BEHAVIORAL of AND2_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_23;

architecture SYN_BEHAVIORAL of AND2_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_22;

architecture SYN_BEHAVIORAL of AND2_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_21;

architecture SYN_BEHAVIORAL of AND2_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_20;

architecture SYN_BEHAVIORAL of AND2_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_19;

architecture SYN_BEHAVIORAL of AND2_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_18;

architecture SYN_BEHAVIORAL of AND2_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_17;

architecture SYN_BEHAVIORAL of AND2_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_16;

architecture SYN_BEHAVIORAL of AND2_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_15;

architecture SYN_BEHAVIORAL of AND2_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_14;

architecture SYN_BEHAVIORAL of AND2_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_13;

architecture SYN_BEHAVIORAL of AND2_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_12;

architecture SYN_BEHAVIORAL of AND2_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_11;

architecture SYN_BEHAVIORAL of AND2_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_10;

architecture SYN_BEHAVIORAL of AND2_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_9;

architecture SYN_BEHAVIORAL of AND2_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_8;

architecture SYN_BEHAVIORAL of AND2_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_7;

architecture SYN_BEHAVIORAL of AND2_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_6;

architecture SYN_BEHAVIORAL of AND2_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_5;

architecture SYN_BEHAVIORAL of AND2_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_4;

architecture SYN_BEHAVIORAL of AND2_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_3;

architecture SYN_BEHAVIORAL of AND2_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_2;

architecture SYN_BEHAVIORAL of AND2_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_1;

architecture SYN_BEHAVIORAL of AND2_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_0;

architecture SYN_BEHAVIORAL of AND2_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_62;

architecture SYN_BEHAVIORAL of XNOR2_62 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_61;

architecture SYN_BEHAVIORAL of XNOR2_61 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_60;

architecture SYN_BEHAVIORAL of XNOR2_60 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_59;

architecture SYN_BEHAVIORAL of XNOR2_59 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_58;

architecture SYN_BEHAVIORAL of XNOR2_58 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_57;

architecture SYN_BEHAVIORAL of XNOR2_57 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_56;

architecture SYN_BEHAVIORAL of XNOR2_56 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_55;

architecture SYN_BEHAVIORAL of XNOR2_55 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_54;

architecture SYN_BEHAVIORAL of XNOR2_54 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_53;

architecture SYN_BEHAVIORAL of XNOR2_53 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_52;

architecture SYN_BEHAVIORAL of XNOR2_52 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_51;

architecture SYN_BEHAVIORAL of XNOR2_51 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_50;

architecture SYN_BEHAVIORAL of XNOR2_50 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_49;

architecture SYN_BEHAVIORAL of XNOR2_49 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_48;

architecture SYN_BEHAVIORAL of XNOR2_48 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_47;

architecture SYN_BEHAVIORAL of XNOR2_47 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_46;

architecture SYN_BEHAVIORAL of XNOR2_46 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_45;

architecture SYN_BEHAVIORAL of XNOR2_45 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_44;

architecture SYN_BEHAVIORAL of XNOR2_44 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_43;

architecture SYN_BEHAVIORAL of XNOR2_43 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_42;

architecture SYN_BEHAVIORAL of XNOR2_42 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_41;

architecture SYN_BEHAVIORAL of XNOR2_41 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_40;

architecture SYN_BEHAVIORAL of XNOR2_40 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_39;

architecture SYN_BEHAVIORAL of XNOR2_39 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_38;

architecture SYN_BEHAVIORAL of XNOR2_38 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_37;

architecture SYN_BEHAVIORAL of XNOR2_37 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_36;

architecture SYN_BEHAVIORAL of XNOR2_36 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_35;

architecture SYN_BEHAVIORAL of XNOR2_35 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_34;

architecture SYN_BEHAVIORAL of XNOR2_34 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_33;

architecture SYN_BEHAVIORAL of XNOR2_33 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_32;

architecture SYN_BEHAVIORAL of XNOR2_32 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_31;

architecture SYN_BEHAVIORAL of XNOR2_31 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_30;

architecture SYN_BEHAVIORAL of XNOR2_30 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_29;

architecture SYN_BEHAVIORAL of XNOR2_29 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_28;

architecture SYN_BEHAVIORAL of XNOR2_28 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_27;

architecture SYN_BEHAVIORAL of XNOR2_27 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_26;

architecture SYN_BEHAVIORAL of XNOR2_26 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_25;

architecture SYN_BEHAVIORAL of XNOR2_25 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_24;

architecture SYN_BEHAVIORAL of XNOR2_24 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_23;

architecture SYN_BEHAVIORAL of XNOR2_23 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_22;

architecture SYN_BEHAVIORAL of XNOR2_22 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_21;

architecture SYN_BEHAVIORAL of XNOR2_21 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_20;

architecture SYN_BEHAVIORAL of XNOR2_20 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_19;

architecture SYN_BEHAVIORAL of XNOR2_19 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_18;

architecture SYN_BEHAVIORAL of XNOR2_18 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_17;

architecture SYN_BEHAVIORAL of XNOR2_17 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_16;

architecture SYN_BEHAVIORAL of XNOR2_16 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_15;

architecture SYN_BEHAVIORAL of XNOR2_15 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_14;

architecture SYN_BEHAVIORAL of XNOR2_14 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_13;

architecture SYN_BEHAVIORAL of XNOR2_13 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_12;

architecture SYN_BEHAVIORAL of XNOR2_12 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_11;

architecture SYN_BEHAVIORAL of XNOR2_11 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_10;

architecture SYN_BEHAVIORAL of XNOR2_10 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_9;

architecture SYN_BEHAVIORAL of XNOR2_9 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_8;

architecture SYN_BEHAVIORAL of XNOR2_8 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_7;

architecture SYN_BEHAVIORAL of XNOR2_7 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_6;

architecture SYN_BEHAVIORAL of XNOR2_6 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_5;

architecture SYN_BEHAVIORAL of XNOR2_5 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_4;

architecture SYN_BEHAVIORAL of XNOR2_4 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_3;

architecture SYN_BEHAVIORAL of XNOR2_3 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_2;

architecture SYN_BEHAVIORAL of XNOR2_2 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_1;

architecture SYN_BEHAVIORAL of XNOR2_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_0;

architecture SYN_BEHAVIORAL of XNOR2_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_30 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_30;

architecture SYN_BEHAVIORAL of FFD_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1215 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1215);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_29 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_29;

architecture SYN_BEHAVIORAL of FFD_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1216 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1216);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_28 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_28;

architecture SYN_BEHAVIORAL of FFD_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1217 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1217);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_27 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_27;

architecture SYN_BEHAVIORAL of FFD_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1218 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1218);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_26 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_26;

architecture SYN_BEHAVIORAL of FFD_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1219 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1219);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_25 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_25;

architecture SYN_BEHAVIORAL of FFD_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1220 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1220);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_24 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_24;

architecture SYN_BEHAVIORAL of FFD_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1221 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1221);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_23 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_23;

architecture SYN_BEHAVIORAL of FFD_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1222 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1222);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_22 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_22;

architecture SYN_BEHAVIORAL of FFD_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1223 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1223);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_21 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_21;

architecture SYN_BEHAVIORAL of FFD_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1224 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1224);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_20 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_20;

architecture SYN_BEHAVIORAL of FFD_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1225 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1225);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_19 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_19;

architecture SYN_BEHAVIORAL of FFD_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1226 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1226);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_18 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_18;

architecture SYN_BEHAVIORAL of FFD_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1227 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1227);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_17 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_17;

architecture SYN_BEHAVIORAL of FFD_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1228 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1228);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_16 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_16;

architecture SYN_BEHAVIORAL of FFD_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1229 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1229);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_15 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_15;

architecture SYN_BEHAVIORAL of FFD_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1230 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1230);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_14 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_14;

architecture SYN_BEHAVIORAL of FFD_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1231 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1231);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_13 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_13;

architecture SYN_BEHAVIORAL of FFD_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1232 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1232);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_12 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_12;

architecture SYN_BEHAVIORAL of FFD_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1233 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1233);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_11 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_11;

architecture SYN_BEHAVIORAL of FFD_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1234 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1234);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_10 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_10;

architecture SYN_BEHAVIORAL of FFD_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1235 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1235);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_9 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_9;

architecture SYN_BEHAVIORAL of FFD_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1236 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1236);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_8 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_8;

architecture SYN_BEHAVIORAL of FFD_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1237 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1237);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_7 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_7;

architecture SYN_BEHAVIORAL of FFD_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1238 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1238);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_6 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_6;

architecture SYN_BEHAVIORAL of FFD_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1239 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1239);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_5 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_5;

architecture SYN_BEHAVIORAL of FFD_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1240 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1240);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_4 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_4;

architecture SYN_BEHAVIORAL of FFD_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1241 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1241);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_3 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_3;

architecture SYN_BEHAVIORAL of FFD_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1242 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1242);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_2 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_2;

architecture SYN_BEHAVIORAL of FFD_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1243 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1243);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_1 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_1;

architecture SYN_BEHAVIORAL of FFD_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1244 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1244);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_0 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_0;

architecture SYN_BEHAVIORAL of FFD_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1245 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1245);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_223 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_223;

architecture SYN_BEHAVIORAL of LD_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_222 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_222;

architecture SYN_BEHAVIORAL of LD_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_221 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_221;

architecture SYN_BEHAVIORAL of LD_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_220 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_220;

architecture SYN_BEHAVIORAL of LD_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_219 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_219;

architecture SYN_BEHAVIORAL of LD_219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_218 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_218;

architecture SYN_BEHAVIORAL of LD_218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_217 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_217;

architecture SYN_BEHAVIORAL of LD_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_216 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_216;

architecture SYN_BEHAVIORAL of LD_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_215 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_215;

architecture SYN_BEHAVIORAL of LD_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_214 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_214;

architecture SYN_BEHAVIORAL of LD_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_213 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_213;

architecture SYN_BEHAVIORAL of LD_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_212 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_212;

architecture SYN_BEHAVIORAL of LD_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_211 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_211;

architecture SYN_BEHAVIORAL of LD_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_210 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_210;

architecture SYN_BEHAVIORAL of LD_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_209 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_209;

architecture SYN_BEHAVIORAL of LD_209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_208 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_208;

architecture SYN_BEHAVIORAL of LD_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_207 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_207;

architecture SYN_BEHAVIORAL of LD_207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_206 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_206;

architecture SYN_BEHAVIORAL of LD_206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_205 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_205;

architecture SYN_BEHAVIORAL of LD_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_204 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_204;

architecture SYN_BEHAVIORAL of LD_204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_203 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_203;

architecture SYN_BEHAVIORAL of LD_203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_202 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_202;

architecture SYN_BEHAVIORAL of LD_202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_201 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_201;

architecture SYN_BEHAVIORAL of LD_201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_200 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_200;

architecture SYN_BEHAVIORAL of LD_200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_199 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_199;

architecture SYN_BEHAVIORAL of LD_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_198 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_198;

architecture SYN_BEHAVIORAL of LD_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_197 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_197;

architecture SYN_BEHAVIORAL of LD_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_196 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_196;

architecture SYN_BEHAVIORAL of LD_196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_195 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_195;

architecture SYN_BEHAVIORAL of LD_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_194 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_194;

architecture SYN_BEHAVIORAL of LD_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_193 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_193;

architecture SYN_BEHAVIORAL of LD_193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_192 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_192;

architecture SYN_BEHAVIORAL of LD_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_191 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_191;

architecture SYN_BEHAVIORAL of LD_191 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_190 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_190;

architecture SYN_BEHAVIORAL of LD_190 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_189 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_189;

architecture SYN_BEHAVIORAL of LD_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_188 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_188;

architecture SYN_BEHAVIORAL of LD_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_187 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_187;

architecture SYN_BEHAVIORAL of LD_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_186 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_186;

architecture SYN_BEHAVIORAL of LD_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_185 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_185;

architecture SYN_BEHAVIORAL of LD_185 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_184 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_184;

architecture SYN_BEHAVIORAL of LD_184 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_183 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_183;

architecture SYN_BEHAVIORAL of LD_183 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_182 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_182;

architecture SYN_BEHAVIORAL of LD_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_181 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_181;

architecture SYN_BEHAVIORAL of LD_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_180 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_180;

architecture SYN_BEHAVIORAL of LD_180 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_179 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_179;

architecture SYN_BEHAVIORAL of LD_179 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_178 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_178;

architecture SYN_BEHAVIORAL of LD_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_177 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_177;

architecture SYN_BEHAVIORAL of LD_177 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_176 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_176;

architecture SYN_BEHAVIORAL of LD_176 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_175 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_175;

architecture SYN_BEHAVIORAL of LD_175 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_174 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_174;

architecture SYN_BEHAVIORAL of LD_174 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_173 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_173;

architecture SYN_BEHAVIORAL of LD_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_172 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_172;

architecture SYN_BEHAVIORAL of LD_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_171 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_171;

architecture SYN_BEHAVIORAL of LD_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_170 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_170;

architecture SYN_BEHAVIORAL of LD_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_169 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_169;

architecture SYN_BEHAVIORAL of LD_169 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_168 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_168;

architecture SYN_BEHAVIORAL of LD_168 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_167 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_167;

architecture SYN_BEHAVIORAL of LD_167 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_166 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_166;

architecture SYN_BEHAVIORAL of LD_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_165 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_165;

architecture SYN_BEHAVIORAL of LD_165 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_164 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_164;

architecture SYN_BEHAVIORAL of LD_164 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_163 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_163;

architecture SYN_BEHAVIORAL of LD_163 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_162 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_162;

architecture SYN_BEHAVIORAL of LD_162 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_161 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_161;

architecture SYN_BEHAVIORAL of LD_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_160 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_160;

architecture SYN_BEHAVIORAL of LD_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_159 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_159;

architecture SYN_BEHAVIORAL of LD_159 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_158 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_158;

architecture SYN_BEHAVIORAL of LD_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_157 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_157;

architecture SYN_BEHAVIORAL of LD_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_156 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_156;

architecture SYN_BEHAVIORAL of LD_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_155 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_155;

architecture SYN_BEHAVIORAL of LD_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_154 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_154;

architecture SYN_BEHAVIORAL of LD_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_153 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_153;

architecture SYN_BEHAVIORAL of LD_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_152 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_152;

architecture SYN_BEHAVIORAL of LD_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_151 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_151;

architecture SYN_BEHAVIORAL of LD_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_150 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_150;

architecture SYN_BEHAVIORAL of LD_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_149 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_149;

architecture SYN_BEHAVIORAL of LD_149 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_148 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_148;

architecture SYN_BEHAVIORAL of LD_148 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_147 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_147;

architecture SYN_BEHAVIORAL of LD_147 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_146 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_146;

architecture SYN_BEHAVIORAL of LD_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_145 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_145;

architecture SYN_BEHAVIORAL of LD_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_144 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_144;

architecture SYN_BEHAVIORAL of LD_144 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_143 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_143;

architecture SYN_BEHAVIORAL of LD_143 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_142 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_142;

architecture SYN_BEHAVIORAL of LD_142 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_141 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_141;

architecture SYN_BEHAVIORAL of LD_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_140 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_140;

architecture SYN_BEHAVIORAL of LD_140 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_139 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_139;

architecture SYN_BEHAVIORAL of LD_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_138 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_138;

architecture SYN_BEHAVIORAL of LD_138 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_137 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_137;

architecture SYN_BEHAVIORAL of LD_137 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_136 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_136;

architecture SYN_BEHAVIORAL of LD_136 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_135 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_135;

architecture SYN_BEHAVIORAL of LD_135 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_134 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_134;

architecture SYN_BEHAVIORAL of LD_134 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_133 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_133;

architecture SYN_BEHAVIORAL of LD_133 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_132 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_132;

architecture SYN_BEHAVIORAL of LD_132 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_131 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_131;

architecture SYN_BEHAVIORAL of LD_131 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_130 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_130;

architecture SYN_BEHAVIORAL of LD_130 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_129 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_129;

architecture SYN_BEHAVIORAL of LD_129 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_128 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_128;

architecture SYN_BEHAVIORAL of LD_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_127 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_127;

architecture SYN_BEHAVIORAL of LD_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_126 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_126;

architecture SYN_BEHAVIORAL of LD_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_125 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_125;

architecture SYN_BEHAVIORAL of LD_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_124 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_124;

architecture SYN_BEHAVIORAL of LD_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_123 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_123;

architecture SYN_BEHAVIORAL of LD_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_122 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_122;

architecture SYN_BEHAVIORAL of LD_122 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_121 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_121;

architecture SYN_BEHAVIORAL of LD_121 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_120 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_120;

architecture SYN_BEHAVIORAL of LD_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_119 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_119;

architecture SYN_BEHAVIORAL of LD_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_118 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_118;

architecture SYN_BEHAVIORAL of LD_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_117 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_117;

architecture SYN_BEHAVIORAL of LD_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_116 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_116;

architecture SYN_BEHAVIORAL of LD_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_115 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_115;

architecture SYN_BEHAVIORAL of LD_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_114 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_114;

architecture SYN_BEHAVIORAL of LD_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_113 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_113;

architecture SYN_BEHAVIORAL of LD_113 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_112 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_112;

architecture SYN_BEHAVIORAL of LD_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_111 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_111;

architecture SYN_BEHAVIORAL of LD_111 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_110 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_110;

architecture SYN_BEHAVIORAL of LD_110 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_109 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_109;

architecture SYN_BEHAVIORAL of LD_109 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_108 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_108;

architecture SYN_BEHAVIORAL of LD_108 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_107 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_107;

architecture SYN_BEHAVIORAL of LD_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_106 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_106;

architecture SYN_BEHAVIORAL of LD_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_105 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_105;

architecture SYN_BEHAVIORAL of LD_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_104 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_104;

architecture SYN_BEHAVIORAL of LD_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_103 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_103;

architecture SYN_BEHAVIORAL of LD_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_102 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_102;

architecture SYN_BEHAVIORAL of LD_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_101 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_101;

architecture SYN_BEHAVIORAL of LD_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_100 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_100;

architecture SYN_BEHAVIORAL of LD_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_99 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_99;

architecture SYN_BEHAVIORAL of LD_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_98 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_98;

architecture SYN_BEHAVIORAL of LD_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_97 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_97;

architecture SYN_BEHAVIORAL of LD_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_96 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_96;

architecture SYN_BEHAVIORAL of LD_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_95 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_95;

architecture SYN_BEHAVIORAL of LD_95 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_94 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_94;

architecture SYN_BEHAVIORAL of LD_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_93 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_93;

architecture SYN_BEHAVIORAL of LD_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_92 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_92;

architecture SYN_BEHAVIORAL of LD_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_91 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_91;

architecture SYN_BEHAVIORAL of LD_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_90 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_90;

architecture SYN_BEHAVIORAL of LD_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_89 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_89;

architecture SYN_BEHAVIORAL of LD_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_88 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_88;

architecture SYN_BEHAVIORAL of LD_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_87 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_87;

architecture SYN_BEHAVIORAL of LD_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_86 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_86;

architecture SYN_BEHAVIORAL of LD_86 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_85 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_85;

architecture SYN_BEHAVIORAL of LD_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_84 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_84;

architecture SYN_BEHAVIORAL of LD_84 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_83 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_83;

architecture SYN_BEHAVIORAL of LD_83 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_82 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_82;

architecture SYN_BEHAVIORAL of LD_82 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_81 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_81;

architecture SYN_BEHAVIORAL of LD_81 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_80 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_80;

architecture SYN_BEHAVIORAL of LD_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_79 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_79;

architecture SYN_BEHAVIORAL of LD_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_78 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_78;

architecture SYN_BEHAVIORAL of LD_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_77 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_77;

architecture SYN_BEHAVIORAL of LD_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_76 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_76;

architecture SYN_BEHAVIORAL of LD_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_75 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_75;

architecture SYN_BEHAVIORAL of LD_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_74 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_74;

architecture SYN_BEHAVIORAL of LD_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_73 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_73;

architecture SYN_BEHAVIORAL of LD_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_72 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_72;

architecture SYN_BEHAVIORAL of LD_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_71 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_71;

architecture SYN_BEHAVIORAL of LD_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_70 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_70;

architecture SYN_BEHAVIORAL of LD_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_69 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_69;

architecture SYN_BEHAVIORAL of LD_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_68 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_68;

architecture SYN_BEHAVIORAL of LD_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_67 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_67;

architecture SYN_BEHAVIORAL of LD_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_66 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_66;

architecture SYN_BEHAVIORAL of LD_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_65 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_65;

architecture SYN_BEHAVIORAL of LD_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_64 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_64;

architecture SYN_BEHAVIORAL of LD_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_63 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_63;

architecture SYN_BEHAVIORAL of LD_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_62 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_62;

architecture SYN_BEHAVIORAL of LD_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_61 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_61;

architecture SYN_BEHAVIORAL of LD_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_60 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_60;

architecture SYN_BEHAVIORAL of LD_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_59 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_59;

architecture SYN_BEHAVIORAL of LD_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_58 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_58;

architecture SYN_BEHAVIORAL of LD_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_57 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_57;

architecture SYN_BEHAVIORAL of LD_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_56 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_56;

architecture SYN_BEHAVIORAL of LD_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_55 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_55;

architecture SYN_BEHAVIORAL of LD_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_54 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_54;

architecture SYN_BEHAVIORAL of LD_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_53 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_53;

architecture SYN_BEHAVIORAL of LD_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_52 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_52;

architecture SYN_BEHAVIORAL of LD_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_51 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_51;

architecture SYN_BEHAVIORAL of LD_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_50 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_50;

architecture SYN_BEHAVIORAL of LD_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_49 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_49;

architecture SYN_BEHAVIORAL of LD_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_48 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_48;

architecture SYN_BEHAVIORAL of LD_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_47 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_47;

architecture SYN_BEHAVIORAL of LD_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_46 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_46;

architecture SYN_BEHAVIORAL of LD_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_45 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_45;

architecture SYN_BEHAVIORAL of LD_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_44 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_44;

architecture SYN_BEHAVIORAL of LD_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_43 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_43;

architecture SYN_BEHAVIORAL of LD_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_42 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_42;

architecture SYN_BEHAVIORAL of LD_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_41 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_41;

architecture SYN_BEHAVIORAL of LD_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_40 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_40;

architecture SYN_BEHAVIORAL of LD_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_39 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_39;

architecture SYN_BEHAVIORAL of LD_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_38 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_38;

architecture SYN_BEHAVIORAL of LD_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_37 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_37;

architecture SYN_BEHAVIORAL of LD_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_36 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_36;

architecture SYN_BEHAVIORAL of LD_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_35 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_35;

architecture SYN_BEHAVIORAL of LD_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_34 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_34;

architecture SYN_BEHAVIORAL of LD_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_33 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_33;

architecture SYN_BEHAVIORAL of LD_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_32 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_32;

architecture SYN_BEHAVIORAL of LD_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_31 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_31;

architecture SYN_BEHAVIORAL of LD_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_30 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_30;

architecture SYN_BEHAVIORAL of LD_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_29 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_29;

architecture SYN_BEHAVIORAL of LD_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_28 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_28;

architecture SYN_BEHAVIORAL of LD_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_27 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_27;

architecture SYN_BEHAVIORAL of LD_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_26 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_26;

architecture SYN_BEHAVIORAL of LD_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_25 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_25;

architecture SYN_BEHAVIORAL of LD_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_24 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_24;

architecture SYN_BEHAVIORAL of LD_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_23 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_23;

architecture SYN_BEHAVIORAL of LD_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_22 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_22;

architecture SYN_BEHAVIORAL of LD_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_21 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_21;

architecture SYN_BEHAVIORAL of LD_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_20 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_20;

architecture SYN_BEHAVIORAL of LD_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_19 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_19;

architecture SYN_BEHAVIORAL of LD_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_18 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_18;

architecture SYN_BEHAVIORAL of LD_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_17 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_17;

architecture SYN_BEHAVIORAL of LD_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_16 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_16;

architecture SYN_BEHAVIORAL of LD_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_15 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_15;

architecture SYN_BEHAVIORAL of LD_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_14 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_14;

architecture SYN_BEHAVIORAL of LD_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_13 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_13;

architecture SYN_BEHAVIORAL of LD_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_12 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_12;

architecture SYN_BEHAVIORAL of LD_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_11 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_11;

architecture SYN_BEHAVIORAL of LD_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_10 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_10;

architecture SYN_BEHAVIORAL of LD_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_9 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_9;

architecture SYN_BEHAVIORAL of LD_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_8 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_8;

architecture SYN_BEHAVIORAL of LD_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_7 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_7;

architecture SYN_BEHAVIORAL of LD_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_6 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_6;

architecture SYN_BEHAVIORAL of LD_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_5 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_5;

architecture SYN_BEHAVIORAL of LD_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_4 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_4;

architecture SYN_BEHAVIORAL of LD_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_3 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_3;

architecture SYN_BEHAVIORAL of LD_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_2 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_2;

architecture SYN_BEHAVIORAL of LD_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_1 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_1;

architecture SYN_BEHAVIORAL of LD_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_0 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_0;

architecture SYN_BEHAVIORAL of LD_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX41_N32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX41_N32_0;

architecture SYN_BEHAVIORAL of MUX41_N32_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n149, Z => n76);
   U2 : BUF_X1 port map( A => n148, Z => n72);
   U3 : BUF_X1 port map( A => n151, Z => n81);
   U4 : BUF_X1 port map( A => n150, Z => n77);
   U5 : INV_X1 port map( A => S(0), ZN => n85);
   U6 : BUF_X1 port map( A => n76, Z => n73);
   U7 : BUF_X1 port map( A => n76, Z => n74);
   U8 : BUF_X1 port map( A => n81, Z => n82);
   U9 : BUF_X1 port map( A => n81, Z => n83);
   U10 : BUF_X1 port map( A => n72, Z => n1);
   U11 : BUF_X1 port map( A => n72, Z => n70);
   U12 : BUF_X1 port map( A => n77, Z => n78);
   U13 : BUF_X1 port map( A => n77, Z => n79);
   U14 : BUF_X1 port map( A => n76, Z => n75);
   U15 : BUF_X1 port map( A => n81, Z => n84);
   U16 : BUF_X1 port map( A => n72, Z => n71);
   U17 : BUF_X1 port map( A => n77, Z => n80);
   U18 : NOR2_X1 port map( A1 => n85, A2 => S(1), ZN => n149);
   U19 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n148);
   U20 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n151);
   U21 : AND2_X1 port map( A1 => S(1), A2 => n85, ZN => n150);
   U22 : AOI22_X1 port map( A1 => B(0), A2 => n73, B1 => A(0), B2 => n1, ZN => 
                           n87);
   U23 : AOI22_X1 port map( A1 => B(1), A2 => n73, B1 => A(1), B2 => n1, ZN => 
                           n109);
   U24 : AOI22_X1 port map( A1 => B(2), A2 => n74, B1 => A(2), B2 => n70, ZN =>
                           n131);
   U25 : AOI22_X1 port map( A1 => B(3), A2 => n75, B1 => A(3), B2 => n71, ZN =>
                           n137);
   U26 : AOI22_X1 port map( A1 => B(4), A2 => n75, B1 => A(4), B2 => n71, ZN =>
                           n139);
   U27 : AOI22_X1 port map( A1 => B(5), A2 => n75, B1 => A(5), B2 => n71, ZN =>
                           n141);
   U28 : AOI22_X1 port map( A1 => B(6), A2 => n75, B1 => A(6), B2 => n71, ZN =>
                           n143);
   U29 : AOI22_X1 port map( A1 => B(7), A2 => n75, B1 => A(7), B2 => n71, ZN =>
                           n145);
   U30 : AOI22_X1 port map( A1 => B(8), A2 => n75, B1 => A(8), B2 => n71, ZN =>
                           n147);
   U31 : AOI22_X1 port map( A1 => B(9), A2 => n75, B1 => A(9), B2 => n71, ZN =>
                           n153);
   U32 : AOI22_X1 port map( A1 => B(10), A2 => n73, B1 => A(10), B2 => n1, ZN 
                           => n89);
   U33 : AOI22_X1 port map( A1 => B(11), A2 => n73, B1 => A(11), B2 => n1, ZN 
                           => n91);
   U34 : AOI22_X1 port map( A1 => B(12), A2 => n73, B1 => A(12), B2 => n1, ZN 
                           => n93);
   U35 : AOI22_X1 port map( A1 => B(13), A2 => n73, B1 => A(13), B2 => n1, ZN 
                           => n95);
   U36 : AOI22_X1 port map( A1 => B(14), A2 => n73, B1 => A(14), B2 => n1, ZN 
                           => n97);
   U37 : AOI22_X1 port map( A1 => B(15), A2 => n73, B1 => A(15), B2 => n1, ZN 
                           => n99);
   U38 : AOI22_X1 port map( A1 => B(16), A2 => n73, B1 => A(16), B2 => n1, ZN 
                           => n101);
   U39 : AOI22_X1 port map( A1 => B(17), A2 => n73, B1 => A(17), B2 => n1, ZN 
                           => n103);
   U40 : AOI22_X1 port map( A1 => B(18), A2 => n73, B1 => A(18), B2 => n1, ZN 
                           => n105);
   U41 : AOI22_X1 port map( A1 => B(19), A2 => n73, B1 => A(19), B2 => n1, ZN 
                           => n107);
   U42 : AOI22_X1 port map( A1 => B(20), A2 => n74, B1 => A(20), B2 => n70, ZN 
                           => n111);
   U43 : AOI22_X1 port map( A1 => B(21), A2 => n74, B1 => A(21), B2 => n70, ZN 
                           => n113);
   U44 : AOI22_X1 port map( A1 => B(22), A2 => n74, B1 => A(22), B2 => n70, ZN 
                           => n115);
   U45 : AOI22_X1 port map( A1 => B(23), A2 => n74, B1 => A(23), B2 => n70, ZN 
                           => n117);
   U46 : AOI22_X1 port map( A1 => B(24), A2 => n74, B1 => A(24), B2 => n70, ZN 
                           => n119);
   U47 : AOI22_X1 port map( A1 => B(25), A2 => n74, B1 => A(25), B2 => n70, ZN 
                           => n121);
   U48 : AOI22_X1 port map( A1 => B(26), A2 => n74, B1 => A(26), B2 => n70, ZN 
                           => n123);
   U49 : AOI22_X1 port map( A1 => B(27), A2 => n74, B1 => A(27), B2 => n70, ZN 
                           => n125);
   U50 : AOI22_X1 port map( A1 => B(28), A2 => n74, B1 => A(28), B2 => n70, ZN 
                           => n127);
   U51 : AOI22_X1 port map( A1 => B(29), A2 => n74, B1 => A(29), B2 => n70, ZN 
                           => n129);
   U52 : AOI22_X1 port map( A1 => B(30), A2 => n74, B1 => A(30), B2 => n70, ZN 
                           => n133);
   U53 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n71, ZN 
                           => n135);
   U54 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Y(0));
   U55 : AOI22_X1 port map( A1 => D(0), A2 => n82, B1 => C(0), B2 => n78, ZN =>
                           n86);
   U56 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Y(1));
   U57 : AOI22_X1 port map( A1 => D(1), A2 => n82, B1 => C(1), B2 => n78, ZN =>
                           n108);
   U58 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Y(2));
   U59 : AOI22_X1 port map( A1 => D(2), A2 => n83, B1 => C(2), B2 => n79, ZN =>
                           n130);
   U60 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Y(3));
   U61 : AOI22_X1 port map( A1 => D(3), A2 => n84, B1 => C(3), B2 => n80, ZN =>
                           n136);
   U62 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Y(4));
   U63 : AOI22_X1 port map( A1 => D(4), A2 => n84, B1 => C(4), B2 => n80, ZN =>
                           n138);
   U64 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Y(5));
   U65 : AOI22_X1 port map( A1 => D(5), A2 => n84, B1 => C(5), B2 => n80, ZN =>
                           n140);
   U66 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Y(6));
   U67 : AOI22_X1 port map( A1 => D(6), A2 => n84, B1 => C(6), B2 => n80, ZN =>
                           n142);
   U68 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Y(7));
   U69 : AOI22_X1 port map( A1 => D(7), A2 => n84, B1 => C(7), B2 => n80, ZN =>
                           n144);
   U70 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Y(8));
   U71 : AOI22_X1 port map( A1 => D(8), A2 => n84, B1 => C(8), B2 => n80, ZN =>
                           n146);
   U72 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Y(10));
   U73 : AOI22_X1 port map( A1 => D(10), A2 => n82, B1 => C(10), B2 => n78, ZN 
                           => n88);
   U74 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Y(11));
   U75 : AOI22_X1 port map( A1 => D(11), A2 => n82, B1 => C(11), B2 => n78, ZN 
                           => n90);
   U76 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Y(12));
   U77 : AOI22_X1 port map( A1 => D(12), A2 => n82, B1 => C(12), B2 => n78, ZN 
                           => n92);
   U78 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Y(13));
   U79 : AOI22_X1 port map( A1 => D(13), A2 => n82, B1 => C(13), B2 => n78, ZN 
                           => n94);
   U80 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Y(14));
   U81 : AOI22_X1 port map( A1 => D(14), A2 => n82, B1 => C(14), B2 => n78, ZN 
                           => n96);
   U82 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Y(15));
   U83 : AOI22_X1 port map( A1 => D(15), A2 => n82, B1 => C(15), B2 => n78, ZN 
                           => n98);
   U84 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Y(16));
   U85 : AOI22_X1 port map( A1 => D(16), A2 => n82, B1 => C(16), B2 => n78, ZN 
                           => n100);
   U86 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Y(17));
   U87 : AOI22_X1 port map( A1 => D(17), A2 => n82, B1 => C(17), B2 => n78, ZN 
                           => n102);
   U88 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Y(18));
   U89 : AOI22_X1 port map( A1 => D(18), A2 => n82, B1 => C(18), B2 => n78, ZN 
                           => n104);
   U90 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Y(19));
   U91 : AOI22_X1 port map( A1 => D(19), A2 => n82, B1 => C(19), B2 => n78, ZN 
                           => n106);
   U92 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Y(20));
   U93 : AOI22_X1 port map( A1 => D(20), A2 => n83, B1 => C(20), B2 => n79, ZN 
                           => n110);
   U94 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Y(21));
   U95 : AOI22_X1 port map( A1 => D(21), A2 => n83, B1 => C(21), B2 => n79, ZN 
                           => n112);
   U96 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Y(22));
   U97 : AOI22_X1 port map( A1 => D(22), A2 => n83, B1 => C(22), B2 => n79, ZN 
                           => n114);
   U98 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Y(23));
   U99 : AOI22_X1 port map( A1 => D(23), A2 => n83, B1 => C(23), B2 => n79, ZN 
                           => n116);
   U100 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Y(24));
   U101 : AOI22_X1 port map( A1 => D(24), A2 => n83, B1 => C(24), B2 => n79, ZN
                           => n118);
   U102 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Y(25));
   U103 : AOI22_X1 port map( A1 => D(25), A2 => n83, B1 => C(25), B2 => n79, ZN
                           => n120);
   U104 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Y(26));
   U105 : AOI22_X1 port map( A1 => D(26), A2 => n83, B1 => C(26), B2 => n79, ZN
                           => n122);
   U106 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Y(27));
   U107 : AOI22_X1 port map( A1 => D(27), A2 => n83, B1 => C(27), B2 => n79, ZN
                           => n124);
   U108 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Y(28));
   U109 : AOI22_X1 port map( A1 => D(28), A2 => n83, B1 => C(28), B2 => n79, ZN
                           => n126);
   U110 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Y(29));
   U111 : AOI22_X1 port map( A1 => D(29), A2 => n83, B1 => C(29), B2 => n79, ZN
                           => n128);
   U112 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Y(30));
   U113 : AOI22_X1 port map( A1 => D(30), A2 => n83, B1 => C(30), B2 => n79, ZN
                           => n132);
   U114 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Y(31));
   U115 : AOI22_X1 port map( A1 => D(31), A2 => n84, B1 => C(31), B2 => n80, ZN
                           => n134);
   U116 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Y(9));
   U117 : AOI22_X1 port map( A1 => D(9), A2 => n84, B1 => C(9), B2 => n80, ZN 
                           => n152);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_5 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_5;

architecture SYN_STRUCTURAL of LDR_N32_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_160
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_161
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_162
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_163
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_164
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_165
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_166
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_167
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_168
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_169
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_170
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_171
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_172
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_173
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_174
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_175
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_176
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_177
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_178
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_179
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_180
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_181
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_182
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_183
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_184
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_185
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_186
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_187
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_188
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_189
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_190
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_191
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_191 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_190 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_189 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_188 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_187 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_186 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_185 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_184 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_183 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_182 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_181 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_180 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_179 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_178 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_177 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_176 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_175 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_174 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_173 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_172 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_171 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_170 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_169 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9))
                           ;
   LDI_8 : LD_168 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8))
                           ;
   LDI_7 : LD_167 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7))
                           ;
   LDI_6 : LD_166 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6))
                           ;
   LDI_5 : LD_165 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5))
                           ;
   LDI_4 : LD_164 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4))
                           ;
   LDI_3 : LD_163 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3))
                           ;
   LDI_2 : LD_162 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2))
                           ;
   LDI_1 : LD_161 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1))
                           ;
   LDI_0 : LD_160 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0))
                           ;
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_4 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_4;

architecture SYN_STRUCTURAL of LDR_N32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_128
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_129
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_130
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_131
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_132
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_133
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_134
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_135
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_136
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_137
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_138
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_139
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_140
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_141
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_142
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_143
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_144
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_145
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_146
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_147
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_148
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_149
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_150
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_151
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_152
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_153
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_154
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_155
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_156
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_157
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_158
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_159
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_159 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_158 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_157 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_156 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_155 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_154 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_153 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_152 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_151 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_150 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_149 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_148 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_147 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_146 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_145 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_144 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_143 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_142 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_141 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_140 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_139 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_138 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_137 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9))
                           ;
   LDI_8 : LD_136 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8))
                           ;
   LDI_7 : LD_135 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7))
                           ;
   LDI_6 : LD_134 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6))
                           ;
   LDI_5 : LD_133 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5))
                           ;
   LDI_4 : LD_132 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4))
                           ;
   LDI_3 : LD_131 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3))
                           ;
   LDI_2 : LD_130 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2))
                           ;
   LDI_1 : LD_129 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1))
                           ;
   LDI_0 : LD_128 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0))
                           ;
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_3 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_3;

architecture SYN_STRUCTURAL of LDR_N32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_96
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_97
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_98
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_99
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_100
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_101
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_102
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_103
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_104
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_105
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_106
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_107
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_108
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_109
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_110
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_111
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_112
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_113
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_114
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_115
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_116
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_117
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_118
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_119
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_120
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_121
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_122
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_123
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_124
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_125
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_126
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_127
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_127 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_126 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_125 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_124 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_123 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_122 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_121 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_120 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_119 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_118 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_117 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_116 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_115 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_114 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_113 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_112 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_111 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_110 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_109 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_108 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_107 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_106 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_105 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9))
                           ;
   LDI_8 : LD_104 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8))
                           ;
   LDI_7 : LD_103 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7))
                           ;
   LDI_6 : LD_102 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6))
                           ;
   LDI_5 : LD_101 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5))
                           ;
   LDI_4 : LD_100 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4))
                           ;
   LDI_3 : LD_99 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3));
   LDI_2 : LD_98 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2));
   LDI_1 : LD_97 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1));
   LDI_0 : LD_96 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_2 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_2;

architecture SYN_STRUCTURAL of LDR_N32_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_64
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_65
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_66
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_67
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_68
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_69
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_70
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_71
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_72
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_73
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_74
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_75
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_76
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_77
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_78
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_79
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_80
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_81
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_82
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_83
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_84
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_85
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_86
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_87
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_88
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_89
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_90
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_91
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_92
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_93
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_94
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_95
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_95 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_94 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_93 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_92 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_91 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_90 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_89 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_88 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_87 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_86 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_85 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_84 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_83 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_82 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_81 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_80 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_79 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_78 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_77 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_76 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_75 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_74 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_73 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9));
   LDI_8 : LD_72 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8));
   LDI_7 : LD_71 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7));
   LDI_6 : LD_70 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6));
   LDI_5 : LD_69 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5));
   LDI_4 : LD_68 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4));
   LDI_3 : LD_67 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3));
   LDI_2 : LD_66 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2));
   LDI_1 : LD_65 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1));
   LDI_0 : LD_64 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_1 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_1;

architecture SYN_STRUCTURAL of LDR_N32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_32
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_33
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_34
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_35
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_36
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_37
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_38
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_39
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_40
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_41
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_42
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_43
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_44
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_45
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_46
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_47
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_48
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_49
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_50
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_51
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_52
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_53
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_54
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_55
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_56
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_57
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_58
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_59
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_60
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_61
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_62
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_63
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_63 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_62 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_61 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_60 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_59 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_58 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_57 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_56 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_55 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_54 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_53 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_52 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_51 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_50 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_49 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_48 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_47 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_46 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_45 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_44 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_43 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_42 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_41 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9));
   LDI_8 : LD_40 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8));
   LDI_7 : LD_39 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7));
   LDI_6 : LD_38 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6));
   LDI_5 : LD_37 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5));
   LDI_4 : LD_36 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4));
   LDI_3 : LD_35 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3));
   LDI_2 : LD_34 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2));
   LDI_1 : LD_33 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1));
   LDI_0 : LD_32 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_0 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_0;

architecture SYN_STRUCTURAL of LDR_N32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_0
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_1
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_2
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_3
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_4
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_5
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_6
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_7
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_8
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_9
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_10
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_11
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_12
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_13
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_14
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_15
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_16
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_17
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_18
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_19
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_20
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_21
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_22
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_23
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_24
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_25
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_26
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_27
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_28
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_29
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_30
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_31
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_31 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_30 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_29 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_28 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_27 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_26 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_25 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_24 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_23 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_22 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_21 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_20 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_19 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_18 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_17 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_16 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_15 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_14 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_13 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_12 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_11 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_10 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_9 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9));
   LDI_8 : LD_8 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8));
   LDI_7 : LD_7 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7));
   LDI_6 : LD_6 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6));
   LDI_5 : LD_5 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5));
   LDI_4 : LD_4 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4));
   LDI_3 : LD_3 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3));
   LDI_2 : LD_2 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2));
   LDI_1 : LD_1 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1));
   LDI_0 : LD_0 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_3;

architecture SYN_BEHAVIORAL of MUX21_N32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n69, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => n69
                           );
   U6 : INV_X1 port map( A => n80, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => n80
                           );
   U8 : INV_X1 port map( A => n91, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => n91
                           );
   U10 : INV_X1 port map( A => n94, ZN => Y(3));
   U11 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U12 : INV_X1 port map( A => n95, ZN => Y(4));
   U13 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U14 : INV_X1 port map( A => n96, ZN => Y(5));
   U15 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U16 : INV_X1 port map( A => n97, ZN => Y(6));
   U17 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U18 : INV_X1 port map( A => n98, ZN => Y(7));
   U19 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U20 : INV_X1 port map( A => n99, ZN => Y(8));
   U21 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U22 : INV_X1 port map( A => n70, ZN => Y(10));
   U23 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U24 : INV_X1 port map( A => n71, ZN => Y(11));
   U25 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U26 : INV_X1 port map( A => n72, ZN => Y(12));
   U27 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U28 : INV_X1 port map( A => n73, ZN => Y(13));
   U29 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U30 : INV_X1 port map( A => n74, ZN => Y(14));
   U31 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U32 : INV_X1 port map( A => n75, ZN => Y(15));
   U33 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U34 : INV_X1 port map( A => n76, ZN => Y(16));
   U35 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U36 : INV_X1 port map( A => n77, ZN => Y(17));
   U37 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U38 : INV_X1 port map( A => n78, ZN => Y(18));
   U39 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U40 : INV_X1 port map( A => n79, ZN => Y(19));
   U41 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U42 : INV_X1 port map( A => n81, ZN => Y(20));
   U43 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U44 : INV_X1 port map( A => n82, ZN => Y(21));
   U45 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U46 : INV_X1 port map( A => n83, ZN => Y(22));
   U47 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U48 : INV_X1 port map( A => n84, ZN => Y(23));
   U49 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U50 : INV_X1 port map( A => n85, ZN => Y(24));
   U51 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U52 : INV_X1 port map( A => n86, ZN => Y(25));
   U53 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U54 : INV_X1 port map( A => n87, ZN => Y(26));
   U55 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U56 : INV_X1 port map( A => n88, ZN => Y(27));
   U57 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U58 : INV_X1 port map( A => n89, ZN => Y(28));
   U59 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U60 : INV_X1 port map( A => n90, ZN => Y(29));
   U61 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U62 : INV_X1 port map( A => n92, ZN => Y(30));
   U63 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U64 : INV_X1 port map( A => n93, ZN => Y(31));
   U65 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U66 : INV_X1 port map( A => n100, ZN => Y(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_2;

architecture SYN_BEHAVIORAL of MUX21_N32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n69, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => n69
                           );
   U6 : INV_X1 port map( A => n80, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => n80
                           );
   U8 : INV_X1 port map( A => n91, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => n91
                           );
   U10 : INV_X1 port map( A => n94, ZN => Y(3));
   U11 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U12 : INV_X1 port map( A => n95, ZN => Y(4));
   U13 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U14 : INV_X1 port map( A => n96, ZN => Y(5));
   U15 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U16 : INV_X1 port map( A => n97, ZN => Y(6));
   U17 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U18 : INV_X1 port map( A => n98, ZN => Y(7));
   U19 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U20 : INV_X1 port map( A => n99, ZN => Y(8));
   U21 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U22 : INV_X1 port map( A => n70, ZN => Y(10));
   U23 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U24 : INV_X1 port map( A => n71, ZN => Y(11));
   U25 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U26 : INV_X1 port map( A => n72, ZN => Y(12));
   U27 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U28 : INV_X1 port map( A => n73, ZN => Y(13));
   U29 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U30 : INV_X1 port map( A => n74, ZN => Y(14));
   U31 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U32 : INV_X1 port map( A => n75, ZN => Y(15));
   U33 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U34 : INV_X1 port map( A => n76, ZN => Y(16));
   U35 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U36 : INV_X1 port map( A => n77, ZN => Y(17));
   U37 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U38 : INV_X1 port map( A => n78, ZN => Y(18));
   U39 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U40 : INV_X1 port map( A => n79, ZN => Y(19));
   U41 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U42 : INV_X1 port map( A => n81, ZN => Y(20));
   U43 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U44 : INV_X1 port map( A => n82, ZN => Y(21));
   U45 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U46 : INV_X1 port map( A => n83, ZN => Y(22));
   U47 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U48 : INV_X1 port map( A => n84, ZN => Y(23));
   U49 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U50 : INV_X1 port map( A => n85, ZN => Y(24));
   U51 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U52 : INV_X1 port map( A => n86, ZN => Y(25));
   U53 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U54 : INV_X1 port map( A => n87, ZN => Y(26));
   U55 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U56 : INV_X1 port map( A => n88, ZN => Y(27));
   U57 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U58 : INV_X1 port map( A => n89, ZN => Y(28));
   U59 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U60 : INV_X1 port map( A => n90, ZN => Y(29));
   U61 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U62 : INV_X1 port map( A => n92, ZN => Y(30));
   U63 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U64 : INV_X1 port map( A => n93, ZN => Y(31));
   U65 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U66 : INV_X1 port map( A => n100, ZN => Y(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_1;

architecture SYN_BEHAVIORAL of MUX21_N32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n93, ZN => Y(31));
   U5 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U6 : INV_X1 port map( A => n69, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => n69
                           );
   U8 : INV_X1 port map( A => n80, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => n80
                           );
   U10 : INV_X1 port map( A => n91, ZN => Y(2));
   U11 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U12 : INV_X1 port map( A => n94, ZN => Y(3));
   U13 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U14 : INV_X1 port map( A => n95, ZN => Y(4));
   U15 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U16 : INV_X1 port map( A => n96, ZN => Y(5));
   U17 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U18 : INV_X1 port map( A => n97, ZN => Y(6));
   U19 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U20 : INV_X1 port map( A => n98, ZN => Y(7));
   U21 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U22 : INV_X1 port map( A => n99, ZN => Y(8));
   U23 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U24 : INV_X1 port map( A => n70, ZN => Y(10));
   U25 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U26 : INV_X1 port map( A => n71, ZN => Y(11));
   U27 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U28 : INV_X1 port map( A => n72, ZN => Y(12));
   U29 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U30 : INV_X1 port map( A => n73, ZN => Y(13));
   U31 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U32 : INV_X1 port map( A => n74, ZN => Y(14));
   U33 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U34 : INV_X1 port map( A => n75, ZN => Y(15));
   U35 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U36 : INV_X1 port map( A => n76, ZN => Y(16));
   U37 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U38 : INV_X1 port map( A => n77, ZN => Y(17));
   U39 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U40 : INV_X1 port map( A => n78, ZN => Y(18));
   U41 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U42 : INV_X1 port map( A => n79, ZN => Y(19));
   U43 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U44 : INV_X1 port map( A => n81, ZN => Y(20));
   U45 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U46 : INV_X1 port map( A => n82, ZN => Y(21));
   U47 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U48 : INV_X1 port map( A => n83, ZN => Y(22));
   U49 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U50 : INV_X1 port map( A => n84, ZN => Y(23));
   U51 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U52 : INV_X1 port map( A => n85, ZN => Y(24));
   U53 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U54 : INV_X1 port map( A => n86, ZN => Y(25));
   U55 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U56 : INV_X1 port map( A => n87, ZN => Y(26));
   U57 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U58 : INV_X1 port map( A => n88, ZN => Y(27));
   U59 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U60 : INV_X1 port map( A => n89, ZN => Y(28));
   U61 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U62 : INV_X1 port map( A => n90, ZN => Y(29));
   U63 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U64 : INV_X1 port map( A => n92, ZN => Y(30));
   U65 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U66 : INV_X1 port map( A => n100, ZN => Y(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_0;

architecture SYN_BEHAVIORAL of MUX21_N32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n93, ZN => Y(31));
   U5 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U6 : INV_X1 port map( A => n69, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => n69
                           );
   U8 : INV_X1 port map( A => n80, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => n80
                           );
   U10 : INV_X1 port map( A => n91, ZN => Y(2));
   U11 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U12 : INV_X1 port map( A => n94, ZN => Y(3));
   U13 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U14 : INV_X1 port map( A => n95, ZN => Y(4));
   U15 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U16 : INV_X1 port map( A => n96, ZN => Y(5));
   U17 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U18 : INV_X1 port map( A => n97, ZN => Y(6));
   U19 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U20 : INV_X1 port map( A => n98, ZN => Y(7));
   U21 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U22 : INV_X1 port map( A => n99, ZN => Y(8));
   U23 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U24 : INV_X1 port map( A => n70, ZN => Y(10));
   U25 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U26 : INV_X1 port map( A => n71, ZN => Y(11));
   U27 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U28 : INV_X1 port map( A => n72, ZN => Y(12));
   U29 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U30 : INV_X1 port map( A => n73, ZN => Y(13));
   U31 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U32 : INV_X1 port map( A => n74, ZN => Y(14));
   U33 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U34 : INV_X1 port map( A => n75, ZN => Y(15));
   U35 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U36 : INV_X1 port map( A => n76, ZN => Y(16));
   U37 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U38 : INV_X1 port map( A => n77, ZN => Y(17));
   U39 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U40 : INV_X1 port map( A => n78, ZN => Y(18));
   U41 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U42 : INV_X1 port map( A => n79, ZN => Y(19));
   U43 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U44 : INV_X1 port map( A => n81, ZN => Y(20));
   U45 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U46 : INV_X1 port map( A => n82, ZN => Y(21));
   U47 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U48 : INV_X1 port map( A => n83, ZN => Y(22));
   U49 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U50 : INV_X1 port map( A => n84, ZN => Y(23));
   U51 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U52 : INV_X1 port map( A => n85, ZN => Y(24));
   U53 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U54 : INV_X1 port map( A => n86, ZN => Y(25));
   U55 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U56 : INV_X1 port map( A => n87, ZN => Y(26));
   U57 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U58 : INV_X1 port map( A => n88, ZN => Y(27));
   U59 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U60 : INV_X1 port map( A => n89, ZN => Y(28));
   U61 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U62 : INV_X1 port map( A => n90, ZN => Y(29));
   U63 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U64 : INV_X1 port map( A => n92, ZN => Y(30));
   U65 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U66 : INV_X1 port map( A => n100, ZN => Y(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_319 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_319;

architecture SYN_BEHAVIORAL of MUX21_L_319 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_318 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_318;

architecture SYN_BEHAVIORAL of MUX21_L_318 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_317 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_317;

architecture SYN_BEHAVIORAL of MUX21_L_317 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_316 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_316;

architecture SYN_BEHAVIORAL of MUX21_L_316 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_315 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_315;

architecture SYN_BEHAVIORAL of MUX21_L_315 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_314 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_314;

architecture SYN_BEHAVIORAL of MUX21_L_314 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_313 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_313;

architecture SYN_BEHAVIORAL of MUX21_L_313 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_312 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_312;

architecture SYN_BEHAVIORAL of MUX21_L_312 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_311 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_311;

architecture SYN_BEHAVIORAL of MUX21_L_311 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_310 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_310;

architecture SYN_BEHAVIORAL of MUX21_L_310 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_309 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_309;

architecture SYN_BEHAVIORAL of MUX21_L_309 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_308 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_308;

architecture SYN_BEHAVIORAL of MUX21_L_308 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_307 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_307;

architecture SYN_BEHAVIORAL of MUX21_L_307 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_306 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_306;

architecture SYN_BEHAVIORAL of MUX21_L_306 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_305 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_305;

architecture SYN_BEHAVIORAL of MUX21_L_305 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_304 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_304;

architecture SYN_BEHAVIORAL of MUX21_L_304 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_303 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_303;

architecture SYN_BEHAVIORAL of MUX21_L_303 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_302 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_302;

architecture SYN_BEHAVIORAL of MUX21_L_302 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_301 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_301;

architecture SYN_BEHAVIORAL of MUX21_L_301 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_300 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_300;

architecture SYN_BEHAVIORAL of MUX21_L_300 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_299 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_299;

architecture SYN_BEHAVIORAL of MUX21_L_299 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_298 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_298;

architecture SYN_BEHAVIORAL of MUX21_L_298 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_297 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_297;

architecture SYN_BEHAVIORAL of MUX21_L_297 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_296 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_296;

architecture SYN_BEHAVIORAL of MUX21_L_296 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_295 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_295;

architecture SYN_BEHAVIORAL of MUX21_L_295 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_294 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_294;

architecture SYN_BEHAVIORAL of MUX21_L_294 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_293 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_293;

architecture SYN_BEHAVIORAL of MUX21_L_293 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_292 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_292;

architecture SYN_BEHAVIORAL of MUX21_L_292 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_291 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_291;

architecture SYN_BEHAVIORAL of MUX21_L_291 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_290 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_290;

architecture SYN_BEHAVIORAL of MUX21_L_290 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_289 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_289;

architecture SYN_BEHAVIORAL of MUX21_L_289 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_288 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_288;

architecture SYN_BEHAVIORAL of MUX21_L_288 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_287 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_287;

architecture SYN_BEHAVIORAL of MUX21_L_287 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_286 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_286;

architecture SYN_BEHAVIORAL of MUX21_L_286 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_285 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_285;

architecture SYN_BEHAVIORAL of MUX21_L_285 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_284 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_284;

architecture SYN_BEHAVIORAL of MUX21_L_284 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_283 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_283;

architecture SYN_BEHAVIORAL of MUX21_L_283 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_282 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_282;

architecture SYN_BEHAVIORAL of MUX21_L_282 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_281 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_281;

architecture SYN_BEHAVIORAL of MUX21_L_281 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_280 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_280;

architecture SYN_BEHAVIORAL of MUX21_L_280 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_279 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_279;

architecture SYN_BEHAVIORAL of MUX21_L_279 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_278 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_278;

architecture SYN_BEHAVIORAL of MUX21_L_278 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_277 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_277;

architecture SYN_BEHAVIORAL of MUX21_L_277 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_276 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_276;

architecture SYN_BEHAVIORAL of MUX21_L_276 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_275 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_275;

architecture SYN_BEHAVIORAL of MUX21_L_275 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_274 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_274;

architecture SYN_BEHAVIORAL of MUX21_L_274 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_273 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_273;

architecture SYN_BEHAVIORAL of MUX21_L_273 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_272 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_272;

architecture SYN_BEHAVIORAL of MUX21_L_272 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_271 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_271;

architecture SYN_BEHAVIORAL of MUX21_L_271 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_270 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_270;

architecture SYN_BEHAVIORAL of MUX21_L_270 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_269 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_269;

architecture SYN_BEHAVIORAL of MUX21_L_269 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_268 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_268;

architecture SYN_BEHAVIORAL of MUX21_L_268 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_267 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_267;

architecture SYN_BEHAVIORAL of MUX21_L_267 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_266 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_266;

architecture SYN_BEHAVIORAL of MUX21_L_266 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_265 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_265;

architecture SYN_BEHAVIORAL of MUX21_L_265 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_264 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_264;

architecture SYN_BEHAVIORAL of MUX21_L_264 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_263 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_263;

architecture SYN_BEHAVIORAL of MUX21_L_263 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_262 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_262;

architecture SYN_BEHAVIORAL of MUX21_L_262 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_261 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_261;

architecture SYN_BEHAVIORAL of MUX21_L_261 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_260 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_260;

architecture SYN_BEHAVIORAL of MUX21_L_260 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_259 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_259;

architecture SYN_BEHAVIORAL of MUX21_L_259 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_258 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_258;

architecture SYN_BEHAVIORAL of MUX21_L_258 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_257 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_257;

architecture SYN_BEHAVIORAL of MUX21_L_257 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_256 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_256;

architecture SYN_BEHAVIORAL of MUX21_L_256 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_255 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_255;

architecture SYN_BEHAVIORAL of MUX21_L_255 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_254 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_254;

architecture SYN_BEHAVIORAL of MUX21_L_254 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_253 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_253;

architecture SYN_BEHAVIORAL of MUX21_L_253 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_252 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_252;

architecture SYN_BEHAVIORAL of MUX21_L_252 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_251 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_251;

architecture SYN_BEHAVIORAL of MUX21_L_251 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_250 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_250;

architecture SYN_BEHAVIORAL of MUX21_L_250 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_249 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_249;

architecture SYN_BEHAVIORAL of MUX21_L_249 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_248 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_248;

architecture SYN_BEHAVIORAL of MUX21_L_248 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_247 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_247;

architecture SYN_BEHAVIORAL of MUX21_L_247 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_246 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_246;

architecture SYN_BEHAVIORAL of MUX21_L_246 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_245 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_245;

architecture SYN_BEHAVIORAL of MUX21_L_245 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_244 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_244;

architecture SYN_BEHAVIORAL of MUX21_L_244 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_243 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_243;

architecture SYN_BEHAVIORAL of MUX21_L_243 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_242 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_242;

architecture SYN_BEHAVIORAL of MUX21_L_242 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_241 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_241;

architecture SYN_BEHAVIORAL of MUX21_L_241 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_240 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_240;

architecture SYN_BEHAVIORAL of MUX21_L_240 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_239 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_239;

architecture SYN_BEHAVIORAL of MUX21_L_239 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_238 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_238;

architecture SYN_BEHAVIORAL of MUX21_L_238 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_237 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_237;

architecture SYN_BEHAVIORAL of MUX21_L_237 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_236 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_236;

architecture SYN_BEHAVIORAL of MUX21_L_236 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_235 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_235;

architecture SYN_BEHAVIORAL of MUX21_L_235 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_234 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_234;

architecture SYN_BEHAVIORAL of MUX21_L_234 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_233 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_233;

architecture SYN_BEHAVIORAL of MUX21_L_233 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_232 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_232;

architecture SYN_BEHAVIORAL of MUX21_L_232 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_231 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_231;

architecture SYN_BEHAVIORAL of MUX21_L_231 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_230 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_230;

architecture SYN_BEHAVIORAL of MUX21_L_230 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_229 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_229;

architecture SYN_BEHAVIORAL of MUX21_L_229 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_228 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_228;

architecture SYN_BEHAVIORAL of MUX21_L_228 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_227 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_227;

architecture SYN_BEHAVIORAL of MUX21_L_227 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_226 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_226;

architecture SYN_BEHAVIORAL of MUX21_L_226 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_225 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_225;

architecture SYN_BEHAVIORAL of MUX21_L_225 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_224 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_224;

architecture SYN_BEHAVIORAL of MUX21_L_224 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_223 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_223;

architecture SYN_BEHAVIORAL of MUX21_L_223 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_222 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_222;

architecture SYN_BEHAVIORAL of MUX21_L_222 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_221 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_221;

architecture SYN_BEHAVIORAL of MUX21_L_221 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_220 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_220;

architecture SYN_BEHAVIORAL of MUX21_L_220 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_219 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_219;

architecture SYN_BEHAVIORAL of MUX21_L_219 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_218 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_218;

architecture SYN_BEHAVIORAL of MUX21_L_218 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_217 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_217;

architecture SYN_BEHAVIORAL of MUX21_L_217 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_216 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_216;

architecture SYN_BEHAVIORAL of MUX21_L_216 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_215 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_215;

architecture SYN_BEHAVIORAL of MUX21_L_215 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_214 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_214;

architecture SYN_BEHAVIORAL of MUX21_L_214 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_213 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_213;

architecture SYN_BEHAVIORAL of MUX21_L_213 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_212 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_212;

architecture SYN_BEHAVIORAL of MUX21_L_212 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_211 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_211;

architecture SYN_BEHAVIORAL of MUX21_L_211 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_210 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_210;

architecture SYN_BEHAVIORAL of MUX21_L_210 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_209 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_209;

architecture SYN_BEHAVIORAL of MUX21_L_209 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_208 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_208;

architecture SYN_BEHAVIORAL of MUX21_L_208 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_207 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_207;

architecture SYN_BEHAVIORAL of MUX21_L_207 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_206 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_206;

architecture SYN_BEHAVIORAL of MUX21_L_206 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_205 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_205;

architecture SYN_BEHAVIORAL of MUX21_L_205 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_204 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_204;

architecture SYN_BEHAVIORAL of MUX21_L_204 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_203 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_203;

architecture SYN_BEHAVIORAL of MUX21_L_203 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_202 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_202;

architecture SYN_BEHAVIORAL of MUX21_L_202 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_201 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_201;

architecture SYN_BEHAVIORAL of MUX21_L_201 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_200 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_200;

architecture SYN_BEHAVIORAL of MUX21_L_200 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_199 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_199;

architecture SYN_BEHAVIORAL of MUX21_L_199 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_198 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_198;

architecture SYN_BEHAVIORAL of MUX21_L_198 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_197 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_197;

architecture SYN_BEHAVIORAL of MUX21_L_197 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_196 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_196;

architecture SYN_BEHAVIORAL of MUX21_L_196 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_195 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_195;

architecture SYN_BEHAVIORAL of MUX21_L_195 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_194 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_194;

architecture SYN_BEHAVIORAL of MUX21_L_194 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_193 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_193;

architecture SYN_BEHAVIORAL of MUX21_L_193 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_192 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_192;

architecture SYN_BEHAVIORAL of MUX21_L_192 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_191 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_191;

architecture SYN_BEHAVIORAL of MUX21_L_191 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_190 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_190;

architecture SYN_BEHAVIORAL of MUX21_L_190 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_189 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_189;

architecture SYN_BEHAVIORAL of MUX21_L_189 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_188 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_188;

architecture SYN_BEHAVIORAL of MUX21_L_188 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_187 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_187;

architecture SYN_BEHAVIORAL of MUX21_L_187 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_186 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_186;

architecture SYN_BEHAVIORAL of MUX21_L_186 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_185 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_185;

architecture SYN_BEHAVIORAL of MUX21_L_185 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_184 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_184;

architecture SYN_BEHAVIORAL of MUX21_L_184 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_183 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_183;

architecture SYN_BEHAVIORAL of MUX21_L_183 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_182 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_182;

architecture SYN_BEHAVIORAL of MUX21_L_182 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_181 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_181;

architecture SYN_BEHAVIORAL of MUX21_L_181 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_180 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_180;

architecture SYN_BEHAVIORAL of MUX21_L_180 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_179 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_179;

architecture SYN_BEHAVIORAL of MUX21_L_179 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_178 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_178;

architecture SYN_BEHAVIORAL of MUX21_L_178 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_177 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_177;

architecture SYN_BEHAVIORAL of MUX21_L_177 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_176 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_176;

architecture SYN_BEHAVIORAL of MUX21_L_176 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_175 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_175;

architecture SYN_BEHAVIORAL of MUX21_L_175 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_174 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_174;

architecture SYN_BEHAVIORAL of MUX21_L_174 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_173 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_173;

architecture SYN_BEHAVIORAL of MUX21_L_173 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_172 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_172;

architecture SYN_BEHAVIORAL of MUX21_L_172 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_171 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_171;

architecture SYN_BEHAVIORAL of MUX21_L_171 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_170 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_170;

architecture SYN_BEHAVIORAL of MUX21_L_170 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_169 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_169;

architecture SYN_BEHAVIORAL of MUX21_L_169 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_168 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_168;

architecture SYN_BEHAVIORAL of MUX21_L_168 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_167 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_167;

architecture SYN_BEHAVIORAL of MUX21_L_167 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_166 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_166;

architecture SYN_BEHAVIORAL of MUX21_L_166 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_165 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_165;

architecture SYN_BEHAVIORAL of MUX21_L_165 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_164 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_164;

architecture SYN_BEHAVIORAL of MUX21_L_164 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_163 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_163;

architecture SYN_BEHAVIORAL of MUX21_L_163 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_162 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_162;

architecture SYN_BEHAVIORAL of MUX21_L_162 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_161 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_161;

architecture SYN_BEHAVIORAL of MUX21_L_161 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_160 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_160;

architecture SYN_BEHAVIORAL of MUX21_L_160 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_159 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_159;

architecture SYN_BEHAVIORAL of MUX21_L_159 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_158 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_158;

architecture SYN_BEHAVIORAL of MUX21_L_158 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_157 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_157;

architecture SYN_BEHAVIORAL of MUX21_L_157 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_156 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_156;

architecture SYN_BEHAVIORAL of MUX21_L_156 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_155 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_155;

architecture SYN_BEHAVIORAL of MUX21_L_155 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_154 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_154;

architecture SYN_BEHAVIORAL of MUX21_L_154 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_153 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_153;

architecture SYN_BEHAVIORAL of MUX21_L_153 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_152 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_152;

architecture SYN_BEHAVIORAL of MUX21_L_152 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_151 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_151;

architecture SYN_BEHAVIORAL of MUX21_L_151 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_150 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_150;

architecture SYN_BEHAVIORAL of MUX21_L_150 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_149 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_149;

architecture SYN_BEHAVIORAL of MUX21_L_149 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_148 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_148;

architecture SYN_BEHAVIORAL of MUX21_L_148 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_147 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_147;

architecture SYN_BEHAVIORAL of MUX21_L_147 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_146 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_146;

architecture SYN_BEHAVIORAL of MUX21_L_146 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_145 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_145;

architecture SYN_BEHAVIORAL of MUX21_L_145 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_144 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_144;

architecture SYN_BEHAVIORAL of MUX21_L_144 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_143 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_143;

architecture SYN_BEHAVIORAL of MUX21_L_143 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_142 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_142;

architecture SYN_BEHAVIORAL of MUX21_L_142 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_141 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_141;

architecture SYN_BEHAVIORAL of MUX21_L_141 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_140 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_140;

architecture SYN_BEHAVIORAL of MUX21_L_140 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_139 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_139;

architecture SYN_BEHAVIORAL of MUX21_L_139 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_138 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_138;

architecture SYN_BEHAVIORAL of MUX21_L_138 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_137 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_137;

architecture SYN_BEHAVIORAL of MUX21_L_137 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_136 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_136;

architecture SYN_BEHAVIORAL of MUX21_L_136 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_135 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_135;

architecture SYN_BEHAVIORAL of MUX21_L_135 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_134 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_134;

architecture SYN_BEHAVIORAL of MUX21_L_134 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_133 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_133;

architecture SYN_BEHAVIORAL of MUX21_L_133 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_132 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_132;

architecture SYN_BEHAVIORAL of MUX21_L_132 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_131 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_131;

architecture SYN_BEHAVIORAL of MUX21_L_131 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_130 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_130;

architecture SYN_BEHAVIORAL of MUX21_L_130 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_129 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_129;

architecture SYN_BEHAVIORAL of MUX21_L_129 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_128 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_128;

architecture SYN_BEHAVIORAL of MUX21_L_128 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_127 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_127;

architecture SYN_BEHAVIORAL of MUX21_L_127 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_126 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_126;

architecture SYN_BEHAVIORAL of MUX21_L_126 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_125 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_125;

architecture SYN_BEHAVIORAL of MUX21_L_125 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_124 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_124;

architecture SYN_BEHAVIORAL of MUX21_L_124 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_123 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_123;

architecture SYN_BEHAVIORAL of MUX21_L_123 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_122 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_122;

architecture SYN_BEHAVIORAL of MUX21_L_122 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_121 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_121;

architecture SYN_BEHAVIORAL of MUX21_L_121 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_120 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_120;

architecture SYN_BEHAVIORAL of MUX21_L_120 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_119 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_119;

architecture SYN_BEHAVIORAL of MUX21_L_119 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_118 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_118;

architecture SYN_BEHAVIORAL of MUX21_L_118 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_117 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_117;

architecture SYN_BEHAVIORAL of MUX21_L_117 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_116 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_116;

architecture SYN_BEHAVIORAL of MUX21_L_116 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_115 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_115;

architecture SYN_BEHAVIORAL of MUX21_L_115 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_114 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_114;

architecture SYN_BEHAVIORAL of MUX21_L_114 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_113 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_113;

architecture SYN_BEHAVIORAL of MUX21_L_113 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_112 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_112;

architecture SYN_BEHAVIORAL of MUX21_L_112 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_111 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_111;

architecture SYN_BEHAVIORAL of MUX21_L_111 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_110 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_110;

architecture SYN_BEHAVIORAL of MUX21_L_110 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_109 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_109;

architecture SYN_BEHAVIORAL of MUX21_L_109 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_108 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_108;

architecture SYN_BEHAVIORAL of MUX21_L_108 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_107 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_107;

architecture SYN_BEHAVIORAL of MUX21_L_107 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_106 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_106;

architecture SYN_BEHAVIORAL of MUX21_L_106 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_105 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_105;

architecture SYN_BEHAVIORAL of MUX21_L_105 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_104 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_104;

architecture SYN_BEHAVIORAL of MUX21_L_104 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_103 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_103;

architecture SYN_BEHAVIORAL of MUX21_L_103 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_102 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_102;

architecture SYN_BEHAVIORAL of MUX21_L_102 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_101 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_101;

architecture SYN_BEHAVIORAL of MUX21_L_101 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_100 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_100;

architecture SYN_BEHAVIORAL of MUX21_L_100 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_99 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_99;

architecture SYN_BEHAVIORAL of MUX21_L_99 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_98 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_98;

architecture SYN_BEHAVIORAL of MUX21_L_98 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_97 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_97;

architecture SYN_BEHAVIORAL of MUX21_L_97 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_96 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_96;

architecture SYN_BEHAVIORAL of MUX21_L_96 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_95 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_95;

architecture SYN_BEHAVIORAL of MUX21_L_95 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_94 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_94;

architecture SYN_BEHAVIORAL of MUX21_L_94 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_93 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_93;

architecture SYN_BEHAVIORAL of MUX21_L_93 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_92 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_92;

architecture SYN_BEHAVIORAL of MUX21_L_92 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_91 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_91;

architecture SYN_BEHAVIORAL of MUX21_L_91 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_90 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_90;

architecture SYN_BEHAVIORAL of MUX21_L_90 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_89 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_89;

architecture SYN_BEHAVIORAL of MUX21_L_89 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_88 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_88;

architecture SYN_BEHAVIORAL of MUX21_L_88 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_87 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_87;

architecture SYN_BEHAVIORAL of MUX21_L_87 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_86 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_86;

architecture SYN_BEHAVIORAL of MUX21_L_86 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_85 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_85;

architecture SYN_BEHAVIORAL of MUX21_L_85 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_84 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_84;

architecture SYN_BEHAVIORAL of MUX21_L_84 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_83 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_83;

architecture SYN_BEHAVIORAL of MUX21_L_83 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_82 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_82;

architecture SYN_BEHAVIORAL of MUX21_L_82 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_81 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_81;

architecture SYN_BEHAVIORAL of MUX21_L_81 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_80 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_80;

architecture SYN_BEHAVIORAL of MUX21_L_80 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_79 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_79;

architecture SYN_BEHAVIORAL of MUX21_L_79 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_78 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_78;

architecture SYN_BEHAVIORAL of MUX21_L_78 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_77 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_77;

architecture SYN_BEHAVIORAL of MUX21_L_77 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_76 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_76;

architecture SYN_BEHAVIORAL of MUX21_L_76 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_75 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_75;

architecture SYN_BEHAVIORAL of MUX21_L_75 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_74 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_74;

architecture SYN_BEHAVIORAL of MUX21_L_74 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_73 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_73;

architecture SYN_BEHAVIORAL of MUX21_L_73 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_72 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_72;

architecture SYN_BEHAVIORAL of MUX21_L_72 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_71 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_71;

architecture SYN_BEHAVIORAL of MUX21_L_71 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_70 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_70;

architecture SYN_BEHAVIORAL of MUX21_L_70 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_69 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_69;

architecture SYN_BEHAVIORAL of MUX21_L_69 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_68 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_68;

architecture SYN_BEHAVIORAL of MUX21_L_68 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_67 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_67;

architecture SYN_BEHAVIORAL of MUX21_L_67 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_66 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_66;

architecture SYN_BEHAVIORAL of MUX21_L_66 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_65 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_65;

architecture SYN_BEHAVIORAL of MUX21_L_65 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_64 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_64;

architecture SYN_BEHAVIORAL of MUX21_L_64 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_63 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_63;

architecture SYN_BEHAVIORAL of MUX21_L_63 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_62 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_62;

architecture SYN_BEHAVIORAL of MUX21_L_62 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_61 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_61;

architecture SYN_BEHAVIORAL of MUX21_L_61 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_60 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_60;

architecture SYN_BEHAVIORAL of MUX21_L_60 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_59 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_59;

architecture SYN_BEHAVIORAL of MUX21_L_59 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_58 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_58;

architecture SYN_BEHAVIORAL of MUX21_L_58 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_57 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_57;

architecture SYN_BEHAVIORAL of MUX21_L_57 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_56 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_56;

architecture SYN_BEHAVIORAL of MUX21_L_56 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_55 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_55;

architecture SYN_BEHAVIORAL of MUX21_L_55 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_54 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_54;

architecture SYN_BEHAVIORAL of MUX21_L_54 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_53 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_53;

architecture SYN_BEHAVIORAL of MUX21_L_53 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_52 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_52;

architecture SYN_BEHAVIORAL of MUX21_L_52 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_51 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_51;

architecture SYN_BEHAVIORAL of MUX21_L_51 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_50 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_50;

architecture SYN_BEHAVIORAL of MUX21_L_50 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_49 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_49;

architecture SYN_BEHAVIORAL of MUX21_L_49 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_48 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_48;

architecture SYN_BEHAVIORAL of MUX21_L_48 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_47 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_47;

architecture SYN_BEHAVIORAL of MUX21_L_47 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_46 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_46;

architecture SYN_BEHAVIORAL of MUX21_L_46 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_45 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_45;

architecture SYN_BEHAVIORAL of MUX21_L_45 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_44 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_44;

architecture SYN_BEHAVIORAL of MUX21_L_44 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_43 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_43;

architecture SYN_BEHAVIORAL of MUX21_L_43 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_42 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_42;

architecture SYN_BEHAVIORAL of MUX21_L_42 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_41 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_41;

architecture SYN_BEHAVIORAL of MUX21_L_41 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_40 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_40;

architecture SYN_BEHAVIORAL of MUX21_L_40 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_39 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_39;

architecture SYN_BEHAVIORAL of MUX21_L_39 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_38 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_38;

architecture SYN_BEHAVIORAL of MUX21_L_38 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_37 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_37;

architecture SYN_BEHAVIORAL of MUX21_L_37 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_36 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_36;

architecture SYN_BEHAVIORAL of MUX21_L_36 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_35 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_35;

architecture SYN_BEHAVIORAL of MUX21_L_35 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_34 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_34;

architecture SYN_BEHAVIORAL of MUX21_L_34 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_33 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_33;

architecture SYN_BEHAVIORAL of MUX21_L_33 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_32 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_32;

architecture SYN_BEHAVIORAL of MUX21_L_32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_31;

architecture SYN_BEHAVIORAL of MUX21_L_31 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_30;

architecture SYN_BEHAVIORAL of MUX21_L_30 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_29;

architecture SYN_BEHAVIORAL of MUX21_L_29 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_28;

architecture SYN_BEHAVIORAL of MUX21_L_28 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_27;

architecture SYN_BEHAVIORAL of MUX21_L_27 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_26;

architecture SYN_BEHAVIORAL of MUX21_L_26 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_25;

architecture SYN_BEHAVIORAL of MUX21_L_25 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_24;

architecture SYN_BEHAVIORAL of MUX21_L_24 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_23;

architecture SYN_BEHAVIORAL of MUX21_L_23 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_22;

architecture SYN_BEHAVIORAL of MUX21_L_22 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_21;

architecture SYN_BEHAVIORAL of MUX21_L_21 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_20;

architecture SYN_BEHAVIORAL of MUX21_L_20 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_19;

architecture SYN_BEHAVIORAL of MUX21_L_19 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_18;

architecture SYN_BEHAVIORAL of MUX21_L_18 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_17;

architecture SYN_BEHAVIORAL of MUX21_L_17 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_16;

architecture SYN_BEHAVIORAL of MUX21_L_16 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_15;

architecture SYN_BEHAVIORAL of MUX21_L_15 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_14;

architecture SYN_BEHAVIORAL of MUX21_L_14 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_13;

architecture SYN_BEHAVIORAL of MUX21_L_13 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_12;

architecture SYN_BEHAVIORAL of MUX21_L_12 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_11;

architecture SYN_BEHAVIORAL of MUX21_L_11 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_10;

architecture SYN_BEHAVIORAL of MUX21_L_10 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_9;

architecture SYN_BEHAVIORAL of MUX21_L_9 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_8;

architecture SYN_BEHAVIORAL of MUX21_L_8 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_7;

architecture SYN_BEHAVIORAL of MUX21_L_7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_6;

architecture SYN_BEHAVIORAL of MUX21_L_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_5;

architecture SYN_BEHAVIORAL of MUX21_L_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_4;

architecture SYN_BEHAVIORAL of MUX21_L_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_3;

architecture SYN_BEHAVIORAL of MUX21_L_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_2;

architecture SYN_BEHAVIORAL of MUX21_L_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_1;

architecture SYN_BEHAVIORAL of MUX21_L_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_0;

architecture SYN_BEHAVIORAL of MUX21_L_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => n1, B2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : BUF_X1 port map( A => S, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_7;

architecture SYN_BEHAVIORAL of MUX21_N4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n5);
   U2 : INV_X1 port map( A => n6, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => S, B2 => B(3), ZN => n6)
                           ;
   U4 : INV_X1 port map( A => n9, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n5, B1 => B(0), B2 => S, ZN => n9)
                           ;
   U6 : INV_X1 port map( A => n8, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n5, B1 => B(1), B2 => S, ZN => n8)
                           ;
   U8 : INV_X1 port map( A => n7, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => S, ZN => n7)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_BEHAVIORAL of RCA_N4_15 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n1, n2, n3, n4, n5
      , n17, n18 : std_logic;

begin
   
   U15 : XOR2_X1 port map( A => n2, B => n5, Z => n7);
   U16 : XOR2_X1 port map( A => n18, B => n8, Z => S(2));
   U17 : XOR2_X1 port map( A => B(2), B => A(2), Z => n8);
   U18 : XOR2_X1 port map( A => n9, B => n10, Z => S(1));
   U19 : XOR2_X1 port map( A => B(1), B => A(1), Z => n10);
   U20 : XOR2_X1 port map( A => A(0), B => n11, Z => S(0));
   U21 : XOR2_X1 port map( A => Ci, B => B(0), Z => n11);
   U1 : INV_X1 port map( A => B(0), ZN => n1);
   U2 : INV_X1 port map( A => A(0), ZN => n4);
   U3 : INV_X1 port map( A => n5, ZN => n17);
   U4 : INV_X1 port map( A => n2, ZN => n3);
   U5 : OAI22_X1 port map( A1 => n6, A2 => n17, B1 => n12, B2 => n3, ZN => Co);
   U6 : AND2_X1 port map( A1 => n17, A2 => n6, ZN => n12);
   U7 : BUF_X1 port map( A => A(3), Z => n5);
   U8 : BUF_X1 port map( A => B(3), Z => n2);
   U9 : AOI22_X1 port map( A1 => n18, A2 => A(2), B1 => n13, B2 => B(2), ZN => 
                           n6);
   U10 : OR2_X1 port map( A1 => A(2), A2 => n18, ZN => n13);
   U11 : INV_X1 port map( A => n14, ZN => n18);
   U12 : AOI22_X1 port map( A1 => n9, A2 => A(1), B1 => n15, B2 => B(1), ZN => 
                           n14);
   U13 : OR2_X1 port map( A1 => A(1), A2 => n9, ZN => n15);
   U14 : OAI21_X1 port map( B1 => n4, B2 => n1, A => n16, ZN => n9);
   U22 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n16);
   U23 : XNOR2_X1 port map( A => n6, B => n7, ZN => S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_7 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_7;

architecture SYN_BEHAVIORAL of ENCODER_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n1, n2, n6 : std_logic;

begin
   
   U10 : XOR2_X1 port map( A => B(0), B => B(1), Z => n4);
   U3 : NOR3_X1 port map( A1 => n2, A2 => n3, A3 => n4, ZN => Y(2));
   U4 : OAI21_X1 port map( B1 => n1, B2 => n6, A => n5, ZN => Y(0));
   U5 : OAI21_X1 port map( B1 => n6, B2 => n2, A => n5, ZN => Y(1));
   U6 : INV_X1 port map( A => n1, ZN => n2);
   U7 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => n5);
   U8 : INV_X1 port map( A => n4, ZN => n6);
   U9 : BUF_X1 port map( A => B(2), Z => n1);
   U11 : AND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_6;

architecture SYN_STRUCTURAL of CSB_N4_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n1, n2, 
      n3, n_1246, n_1247 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_13 port map( A(3) => n3, A(2) => A(2), A(1) => A(1), A(0) => 
                           n2, B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0) 
                           => n1, Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1246);
   RCA1 : RCA_N4_12 port map( A(3) => n3, A(2) => A(2), A(1) => A(1), A(0) => 
                           n2, B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0) 
                           => n1, Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1247);
   MUX : MUX21_N4_6 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : BUF_X1 port map( A => A(0), Z => n2);
   U4 : BUF_X1 port map( A => B(0), Z => n1);
   U5 : BUF_X1 port map( A => A(3), Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_7;

architecture SYN_STRUCTURAL of CSB_N4_7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n1, n2, 
      n3, n4, n_1248, n_1249 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_15 port map( A(3) => n4, A(2) => A(2), A(1) => A(1), A(0) => 
                           n3, B(3) => n2, B(2) => B(2), B(1) => B(1), B(0) => 
                           n1, Ci => X_Logic0_port, S(3) => SUM0_3_port, S(2) 
                           => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1248);
   RCA1 : RCA_N4_14 port map( A(3) => n4, A(2) => A(2), A(1) => A(1), A(0) => 
                           n3, B(3) => n2, B(2) => B(2), B(1) => B(1), B(0) => 
                           n1, Ci => X_Logic1_port, S(3) => SUM1_3_port, S(2) 
                           => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1249);
   MUX : MUX21_N4_7 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : BUF_X1 port map( A => B(0), Z => n1);
   U4 : BUF_X1 port map( A => A(0), Z => n3);
   U5 : BUF_X1 port map( A => B(3), Z => n2);
   U6 : BUF_X1 port map( A => A(3), Z => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_33 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_33;

architecture SYN_BEHAVIORAL of PG_BLOCK_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gkj, B2 => Pik, A => Gik, ZN => n2);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_8 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_8;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_ROW_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  P, G : 
         out std_logic_vector (31 downto 0));

end PG_ROW_N32;

architecture SYN_BEHAVIORAL of PG_ROW_N32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n1, n2, n4 : std_logic;

begin
   
   U37 : XOR2_X1 port map( A => B(9), B => A(9), Z => P(9));
   U38 : XOR2_X1 port map( A => B(8), B => A(8), Z => P(8));
   U39 : XOR2_X1 port map( A => B(7), B => A(7), Z => P(7));
   U40 : XOR2_X1 port map( A => B(6), B => A(6), Z => P(6));
   U41 : XOR2_X1 port map( A => B(5), B => A(5), Z => P(5));
   U42 : XOR2_X1 port map( A => B(4), B => A(4), Z => P(4));
   U43 : XOR2_X1 port map( A => B(3), B => A(3), Z => P(3));
   U44 : XOR2_X1 port map( A => B(31), B => A(31), Z => P(31));
   U45 : XOR2_X1 port map( A => B(30), B => A(30), Z => P(30));
   U46 : XOR2_X1 port map( A => B(2), B => A(2), Z => P(2));
   U47 : XOR2_X1 port map( A => B(29), B => A(29), Z => P(29));
   U48 : XOR2_X1 port map( A => B(28), B => A(28), Z => P(28));
   U49 : XOR2_X1 port map( A => B(27), B => A(27), Z => P(27));
   U50 : XOR2_X1 port map( A => B(26), B => A(26), Z => P(26));
   U51 : XOR2_X1 port map( A => B(25), B => A(25), Z => P(25));
   U52 : XOR2_X1 port map( A => B(24), B => A(24), Z => P(24));
   U53 : XOR2_X1 port map( A => B(23), B => A(23), Z => P(23));
   U54 : XOR2_X1 port map( A => B(22), B => A(22), Z => P(22));
   U55 : XOR2_X1 port map( A => B(21), B => A(21), Z => P(21));
   U56 : XOR2_X1 port map( A => B(20), B => A(20), Z => P(20));
   U57 : XOR2_X1 port map( A => B(1), B => A(1), Z => P(1));
   U58 : XOR2_X1 port map( A => B(19), B => A(19), Z => P(19));
   U59 : XOR2_X1 port map( A => B(18), B => A(18), Z => P(18));
   U60 : XOR2_X1 port map( A => B(17), B => A(17), Z => P(17));
   U61 : XOR2_X1 port map( A => B(16), B => A(16), Z => P(16));
   U62 : XOR2_X1 port map( A => B(15), B => A(15), Z => P(15));
   U63 : XOR2_X1 port map( A => B(14), B => A(14), Z => P(14));
   U64 : XOR2_X1 port map( A => B(13), B => A(13), Z => P(13));
   U65 : XOR2_X1 port map( A => B(12), B => A(12), Z => P(12));
   U66 : XOR2_X1 port map( A => B(11), B => A(11), Z => P(11));
   U67 : XOR2_X1 port map( A => B(10), B => A(10), Z => P(10));
   U1 : XNOR2_X1 port map( A => n2, B => A(0), ZN => P(0));
   U2 : INV_X1 port map( A => n1, ZN => n2);
   U3 : BUF_X1 port map( A => B(0), Z => n1);
   U4 : INV_X1 port map( A => A(0), ZN => n4);
   U5 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => G(1));
   U6 : OAI21_X1 port map( B1 => n2, B2 => n4, A => n3, ZN => G(0));
   U7 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => G(2));
   U8 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => G(3));
   U9 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => G(4));
   U10 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => G(5));
   U11 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => G(8));
   U12 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => G(9));
   U13 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => G(6));
   U14 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => G(7));
   U15 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => G(10));
   U16 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => G(11));
   U17 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => G(17));
   U18 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => G(16));
   U19 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => G(25));
   U20 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => G(24));
   U21 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => G(29));
   U22 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => G(28));
   U23 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => G(19));
   U24 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => G(18));
   U25 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => G(27));
   U26 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => G(26));
   U27 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => G(31));
   U28 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => G(30));
   U29 : OAI21_X1 port map( B1 => A(0), B2 => n1, A => Ci, ZN => n3);
   U30 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => G(21));
   U31 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => G(20));
   U32 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => G(23));
   U33 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => G(22));
   U34 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => G(14));
   U35 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => G(15));
   U36 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => G(12));
   U68 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => G(13));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_N32_2;

architecture SYN_BEHAVIORAL of RCA_N32_2 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, 
      n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104
      , n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47 : std_logic;

begin
   
   U129 : XOR2_X1 port map( A => n48, B => n49, Z => S(9));
   U130 : XOR2_X1 port map( A => B(9), B => A(9), Z => n49);
   U131 : XOR2_X1 port map( A => B(8), B => A(8), Z => n51);
   U132 : XOR2_X1 port map( A => n52, B => n53, Z => S(7));
   U133 : XOR2_X1 port map( A => B(7), B => A(7), Z => n53);
   U134 : XOR2_X1 port map( A => B(6), B => A(6), Z => n55);
   U135 : XOR2_X1 port map( A => n56, B => n57, Z => S(5));
   U136 : XOR2_X1 port map( A => B(5), B => A(5), Z => n57);
   U137 : XOR2_X1 port map( A => B(4), B => A(4), Z => n59);
   U138 : XOR2_X1 port map( A => B(3), B => A(3), Z => n61);
   U139 : XOR2_X1 port map( A => n2, B => n62, Z => S(31));
   U140 : XOR2_X1 port map( A => B(31), B => A(31), Z => n62);
   U141 : XOR2_X1 port map( A => n63, B => n64, Z => S(30));
   U142 : XOR2_X1 port map( A => B(30), B => A(30), Z => n64);
   U143 : XOR2_X1 port map( A => B(2), B => A(2), Z => n66);
   U144 : XOR2_X1 port map( A => B(28), B => A(28), Z => n69);
   U145 : XOR2_X1 port map( A => n70, B => n71, Z => S(27));
   U146 : XOR2_X1 port map( A => B(27), B => A(27), Z => n71);
   U147 : XOR2_X1 port map( A => B(26), B => A(26), Z => n73);
   U148 : XOR2_X1 port map( A => n74, B => n75, Z => S(25));
   U149 : XOR2_X1 port map( A => B(25), B => A(25), Z => n75);
   U150 : XOR2_X1 port map( A => B(24), B => A(24), Z => n77);
   U151 : XOR2_X1 port map( A => n78, B => n79, Z => S(23));
   U152 : XOR2_X1 port map( A => B(23), B => A(23), Z => n79);
   U153 : XOR2_X1 port map( A => B(22), B => A(22), Z => n81);
   U154 : XOR2_X1 port map( A => n82, B => n83, Z => S(21));
   U155 : XOR2_X1 port map( A => B(21), B => A(21), Z => n83);
   U156 : XOR2_X1 port map( A => B(20), B => A(20), Z => n85);
   U157 : XOR2_X1 port map( A => B(1), B => A(1), Z => n87);
   U158 : XOR2_X1 port map( A => n88, B => n89, Z => S(19));
   U159 : XOR2_X1 port map( A => B(19), B => A(19), Z => n89);
   U160 : XOR2_X1 port map( A => B(18), B => A(18), Z => n91);
   U161 : XOR2_X1 port map( A => n92, B => n93, Z => S(17));
   U162 : XOR2_X1 port map( A => B(17), B => A(17), Z => n93);
   U163 : XOR2_X1 port map( A => B(16), B => A(16), Z => n95);
   U164 : XOR2_X1 port map( A => n96, B => n97, Z => S(15));
   U165 : XOR2_X1 port map( A => B(15), B => A(15), Z => n97);
   U166 : XOR2_X1 port map( A => B(14), B => A(14), Z => n99);
   U167 : XOR2_X1 port map( A => n100, B => n101, Z => S(13));
   U168 : XOR2_X1 port map( A => B(13), B => A(13), Z => n101);
   U169 : XOR2_X1 port map( A => B(12), B => A(12), Z => n103);
   U170 : XOR2_X1 port map( A => n104, B => n105, Z => S(11));
   U171 : XOR2_X1 port map( A => B(11), B => A(11), Z => n105);
   U172 : XOR2_X1 port map( A => n34, B => n106, Z => S(10));
   U173 : XOR2_X1 port map( A => B(10), B => A(10), Z => n106);
   U174 : XOR2_X1 port map( A => A(0), B => n107, Z => S(0));
   U175 : XOR2_X1 port map( A => Ci, B => B(0), Z => n107);
   U1 : INV_X1 port map( A => n112, ZN => n5);
   U2 : OAI21_X1 port map( B1 => n108, B2 => n1, A => n109, ZN => Co);
   U3 : INV_X1 port map( A => n131, ZN => n34);
   U4 : INV_X1 port map( A => n108, ZN => n2);
   U5 : AOI22_X1 port map( A1 => n44, A2 => A(3), B1 => n139, B2 => B(3), ZN =>
                           n58);
   U6 : OR2_X1 port map( A1 => A(3), A2 => n44, ZN => n139);
   U7 : INV_X1 port map( A => n60, ZN => n44);
   U8 : AOI21_X1 port map( B1 => n56, B2 => A(5), A => n41, ZN => n54);
   U9 : INV_X1 port map( A => n137, ZN => n41);
   U10 : OAI21_X1 port map( B1 => A(5), B2 => n56, A => B(5), ZN => n137);
   U11 : AOI21_X1 port map( B1 => n52, B2 => A(7), A => n38, ZN => n50);
   U12 : INV_X1 port map( A => n135, ZN => n38);
   U13 : OAI21_X1 port map( B1 => A(7), B2 => n52, A => B(7), ZN => n135);
   U14 : AOI21_X1 port map( B1 => n104, B2 => A(11), A => n32, ZN => n102);
   U15 : INV_X1 port map( A => n130, ZN => n32);
   U16 : OAI21_X1 port map( B1 => A(11), B2 => n104, A => B(11), ZN => n130);
   U17 : AOI21_X1 port map( B1 => n100, B2 => A(13), A => n29, ZN => n98);
   U18 : INV_X1 port map( A => n128, ZN => n29);
   U19 : OAI21_X1 port map( B1 => A(13), B2 => n100, A => B(13), ZN => n128);
   U20 : AOI21_X1 port map( B1 => n96, B2 => A(15), A => n26, ZN => n94);
   U21 : INV_X1 port map( A => n126, ZN => n26);
   U22 : OAI21_X1 port map( B1 => A(15), B2 => n96, A => B(15), ZN => n126);
   U23 : AOI21_X1 port map( B1 => n92, B2 => A(17), A => n23, ZN => n90);
   U24 : INV_X1 port map( A => n124, ZN => n23);
   U25 : OAI21_X1 port map( B1 => A(17), B2 => n92, A => B(17), ZN => n124);
   U26 : AOI21_X1 port map( B1 => n88, B2 => A(19), A => n20, ZN => n84);
   U27 : INV_X1 port map( A => n122, ZN => n20);
   U28 : OAI21_X1 port map( B1 => A(19), B2 => n88, A => B(19), ZN => n122);
   U29 : AOI21_X1 port map( B1 => n82, B2 => A(21), A => n17, ZN => n80);
   U30 : INV_X1 port map( A => n120, ZN => n17);
   U31 : OAI21_X1 port map( B1 => A(21), B2 => n82, A => B(21), ZN => n120);
   U32 : AOI21_X1 port map( B1 => n78, B2 => A(23), A => n14, ZN => n76);
   U33 : INV_X1 port map( A => n118, ZN => n14);
   U34 : OAI21_X1 port map( B1 => A(23), B2 => n78, A => B(23), ZN => n118);
   U35 : AOI21_X1 port map( B1 => n74, B2 => A(25), A => n11, ZN => n72);
   U36 : INV_X1 port map( A => n116, ZN => n11);
   U37 : OAI21_X1 port map( B1 => A(25), B2 => n74, A => B(25), ZN => n116);
   U38 : AOI21_X1 port map( B1 => n70, B2 => A(27), A => n8, ZN => n68);
   U39 : INV_X1 port map( A => n114, ZN => n8);
   U40 : OAI21_X1 port map( B1 => A(27), B2 => n70, A => B(27), ZN => n114);
   U41 : OAI21_X1 port map( B1 => n58, B2 => n42, A => n138, ZN => n56);
   U42 : INV_X1 port map( A => A(4), ZN => n42);
   U43 : OAI21_X1 port map( B1 => A(4), B2 => n43, A => B(4), ZN => n138);
   U44 : INV_X1 port map( A => n58, ZN => n43);
   U45 : OAI21_X1 port map( B1 => n54, B2 => n39, A => n136, ZN => n52);
   U46 : INV_X1 port map( A => A(6), ZN => n39);
   U47 : OAI21_X1 port map( B1 => A(6), B2 => n40, A => B(6), ZN => n136);
   U48 : INV_X1 port map( A => n54, ZN => n40);
   U49 : OAI21_X1 port map( B1 => n50, B2 => n36, A => n134, ZN => n48);
   U50 : INV_X1 port map( A => A(8), ZN => n36);
   U51 : OAI21_X1 port map( B1 => A(8), B2 => n37, A => B(8), ZN => n134);
   U52 : INV_X1 port map( A => n50, ZN => n37);
   U53 : OAI21_X1 port map( B1 => n102, B2 => n30, A => n129, ZN => n100);
   U54 : INV_X1 port map( A => A(12), ZN => n30);
   U55 : OAI21_X1 port map( B1 => A(12), B2 => n31, A => B(12), ZN => n129);
   U56 : INV_X1 port map( A => n102, ZN => n31);
   U57 : OAI21_X1 port map( B1 => n98, B2 => n27, A => n127, ZN => n96);
   U58 : INV_X1 port map( A => A(14), ZN => n27);
   U59 : OAI21_X1 port map( B1 => A(14), B2 => n28, A => B(14), ZN => n127);
   U60 : INV_X1 port map( A => n98, ZN => n28);
   U61 : OAI21_X1 port map( B1 => n94, B2 => n24, A => n125, ZN => n92);
   U62 : INV_X1 port map( A => A(16), ZN => n24);
   U63 : OAI21_X1 port map( B1 => A(16), B2 => n25, A => B(16), ZN => n125);
   U64 : INV_X1 port map( A => n94, ZN => n25);
   U65 : OAI21_X1 port map( B1 => n90, B2 => n21, A => n123, ZN => n88);
   U66 : INV_X1 port map( A => A(18), ZN => n21);
   U67 : OAI21_X1 port map( B1 => A(18), B2 => n22, A => B(18), ZN => n123);
   U68 : INV_X1 port map( A => n90, ZN => n22);
   U69 : OAI21_X1 port map( B1 => n84, B2 => n18, A => n121, ZN => n82);
   U70 : INV_X1 port map( A => A(20), ZN => n18);
   U71 : OAI21_X1 port map( B1 => A(20), B2 => n19, A => B(20), ZN => n121);
   U72 : INV_X1 port map( A => n84, ZN => n19);
   U73 : OAI21_X1 port map( B1 => n80, B2 => n15, A => n119, ZN => n78);
   U74 : INV_X1 port map( A => A(22), ZN => n15);
   U75 : OAI21_X1 port map( B1 => A(22), B2 => n16, A => B(22), ZN => n119);
   U76 : INV_X1 port map( A => n80, ZN => n16);
   U77 : OAI21_X1 port map( B1 => n76, B2 => n12, A => n117, ZN => n74);
   U78 : INV_X1 port map( A => A(24), ZN => n12);
   U79 : OAI21_X1 port map( B1 => A(24), B2 => n13, A => B(24), ZN => n117);
   U80 : INV_X1 port map( A => n76, ZN => n13);
   U81 : OAI21_X1 port map( B1 => n72, B2 => n9, A => n115, ZN => n70);
   U82 : INV_X1 port map( A => A(26), ZN => n9);
   U83 : OAI21_X1 port map( B1 => A(26), B2 => n10, A => B(26), ZN => n115);
   U84 : INV_X1 port map( A => n72, ZN => n10);
   U85 : OAI21_X1 port map( B1 => n131, B2 => n33, A => n132, ZN => n104);
   U86 : INV_X1 port map( A => A(10), ZN => n33);
   U87 : OAI21_X1 port map( B1 => A(10), B2 => n34, A => B(10), ZN => n132);
   U88 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n111, ZN => n63);
   U89 : OAI21_X1 port map( B1 => A(29), B2 => n112, A => B(29), ZN => n111);
   U90 : AOI22_X1 port map( A1 => n45, A2 => A(2), B1 => n140, B2 => B(2), ZN 
                           => n60);
   U91 : OR2_X1 port map( A1 => A(2), A2 => n45, ZN => n140);
   U92 : INV_X1 port map( A => n65, ZN => n45);
   U93 : AOI21_X1 port map( B1 => n48, B2 => A(9), A => n35, ZN => n131);
   U94 : INV_X1 port map( A => n133, ZN => n35);
   U95 : OAI21_X1 port map( B1 => A(9), B2 => n48, A => B(9), ZN => n133);
   U96 : AOI21_X1 port map( B1 => n63, B2 => A(30), A => n3, ZN => n108);
   U97 : INV_X1 port map( A => n110, ZN => n3);
   U98 : OAI21_X1 port map( B1 => A(30), B2 => n63, A => B(30), ZN => n110);
   U99 : XNOR2_X1 port map( A => n5, B => n67, ZN => S(29));
   U100 : XNOR2_X1 port map( A => B(29), B => n4, ZN => n67);
   U101 : OAI21_X1 port map( B1 => n68, B2 => n6, A => n113, ZN => n112);
   U102 : INV_X1 port map( A => A(28), ZN => n6);
   U103 : OAI21_X1 port map( B1 => A(28), B2 => n7, A => B(28), ZN => n113);
   U104 : INV_X1 port map( A => n68, ZN => n7);
   U105 : XNOR2_X1 port map( A => n60, B => n61, ZN => S(3));
   U106 : XNOR2_X1 port map( A => n58, B => n59, ZN => S(4));
   U107 : XNOR2_X1 port map( A => n54, B => n55, ZN => S(6));
   U108 : XNOR2_X1 port map( A => n50, B => n51, ZN => S(8));
   U109 : XNOR2_X1 port map( A => n102, B => n103, ZN => S(12));
   U110 : XNOR2_X1 port map( A => n98, B => n99, ZN => S(14));
   U111 : XNOR2_X1 port map( A => n94, B => n95, ZN => S(16));
   U112 : XNOR2_X1 port map( A => n90, B => n91, ZN => S(18));
   U113 : XNOR2_X1 port map( A => n84, B => n85, ZN => S(20));
   U114 : XNOR2_X1 port map( A => n80, B => n81, ZN => S(22));
   U115 : XNOR2_X1 port map( A => n76, B => n77, ZN => S(24));
   U116 : XNOR2_X1 port map( A => n72, B => n73, ZN => S(26));
   U117 : XNOR2_X1 port map( A => n68, B => n69, ZN => S(28));
   U118 : AOI22_X1 port map( A1 => n46, A2 => A(1), B1 => n141, B2 => B(1), ZN 
                           => n65);
   U119 : OR2_X1 port map( A1 => A(1), A2 => n46, ZN => n141);
   U120 : INV_X1 port map( A => n86, ZN => n46);
   U121 : OAI21_X1 port map( B1 => A(31), B2 => n2, A => B(31), ZN => n109);
   U122 : XNOR2_X1 port map( A => n86, B => n87, ZN => S(1));
   U123 : XNOR2_X1 port map( A => n65, B => n66, ZN => S(2));
   U124 : INV_X1 port map( A => A(29), ZN => n4);
   U125 : INV_X1 port map( A => A(31), ZN => n1);
   U126 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n47, ZN => n86);
   U127 : INV_X1 port map( A => n142, ZN => n47);
   U128 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n142);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX81_N32_3 is

   port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX81_N32_3;

architecture SYN_BEHAVIORAL of MUX81_N32_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n1, n2,
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n11, Z => n152);
   U2 : BUF_X1 port map( A => n12, Z => n148);
   U3 : BUF_X1 port map( A => n13, Z => n144);
   U4 : BUF_X1 port map( A => n14, Z => n140);
   U5 : BUF_X1 port map( A => n9, Z => n157);
   U6 : BUF_X1 port map( A => n10, Z => n153);
   U7 : BUF_X1 port map( A => n7, Z => n165);
   U8 : BUF_X1 port map( A => n8, Z => n161);
   U9 : AOI22_X1 port map( A1 => D(16), A2 => n149, B1 => C(16), B2 => n145, ZN
                           => n108);
   U10 : AOI22_X1 port map( A1 => D(1), A2 => n149, B1 => C(1), B2 => n145, ZN 
                           => n92);
   U11 : AOI22_X1 port map( A1 => D(2), A2 => n150, B1 => C(2), B2 => n146, ZN 
                           => n48);
   U12 : AOI22_X1 port map( A1 => D(3), A2 => n151, B1 => C(3), B2 => n147, ZN 
                           => n36);
   U13 : AOI22_X1 port map( A1 => D(4), A2 => n151, B1 => C(4), B2 => n147, ZN 
                           => n32);
   U14 : AOI22_X1 port map( A1 => D(5), A2 => n151, B1 => C(5), B2 => n147, ZN 
                           => n28);
   U15 : AOI22_X1 port map( A1 => D(6), A2 => n151, B1 => C(6), B2 => n147, ZN 
                           => n24);
   U16 : AOI22_X1 port map( A1 => D(7), A2 => n151, B1 => C(7), B2 => n147, ZN 
                           => n20);
   U17 : AOI22_X1 port map( A1 => D(8), A2 => n151, B1 => C(8), B2 => n147, ZN 
                           => n16);
   U18 : AOI22_X1 port map( A1 => D(9), A2 => n151, B1 => C(9), B2 => n147, ZN 
                           => n4);
   U19 : AOI22_X1 port map( A1 => D(10), A2 => n149, B1 => C(10), B2 => n145, 
                           ZN => n132);
   U20 : AOI22_X1 port map( A1 => D(11), A2 => n149, B1 => C(11), B2 => n145, 
                           ZN => n128);
   U21 : AOI22_X1 port map( A1 => D(12), A2 => n149, B1 => C(12), B2 => n145, 
                           ZN => n124);
   U22 : AOI22_X1 port map( A1 => D(13), A2 => n149, B1 => C(13), B2 => n145, 
                           ZN => n120);
   U23 : AOI22_X1 port map( A1 => D(14), A2 => n149, B1 => C(14), B2 => n145, 
                           ZN => n116);
   U24 : AOI22_X1 port map( A1 => D(15), A2 => n149, B1 => C(15), B2 => n145, 
                           ZN => n112);
   U25 : INV_X1 port map( A => S(1), ZN => n170);
   U26 : INV_X1 port map( A => S(0), ZN => n169);
   U27 : BUF_X1 port map( A => n152, Z => n149);
   U28 : BUF_X1 port map( A => n144, Z => n141);
   U29 : BUF_X1 port map( A => n152, Z => n150);
   U30 : BUF_X1 port map( A => n144, Z => n142);
   U31 : BUF_X1 port map( A => n157, Z => n158);
   U32 : BUF_X1 port map( A => n165, Z => n166);
   U33 : BUF_X1 port map( A => n157, Z => n159);
   U34 : BUF_X1 port map( A => n165, Z => n167);
   U35 : BUF_X1 port map( A => n148, Z => n145);
   U36 : BUF_X1 port map( A => n140, Z => n1);
   U37 : BUF_X1 port map( A => n148, Z => n146);
   U38 : BUF_X1 port map( A => n140, Z => n2);
   U39 : BUF_X1 port map( A => n153, Z => n154);
   U40 : BUF_X1 port map( A => n161, Z => n162);
   U41 : BUF_X1 port map( A => n153, Z => n155);
   U42 : BUF_X1 port map( A => n161, Z => n163);
   U43 : BUF_X1 port map( A => n152, Z => n151);
   U44 : BUF_X1 port map( A => n144, Z => n143);
   U45 : BUF_X1 port map( A => n148, Z => n147);
   U46 : BUF_X1 port map( A => n140, Z => n139);
   U47 : BUF_X1 port map( A => n157, Z => n160);
   U48 : BUF_X1 port map( A => n165, Z => n168);
   U49 : BUF_X1 port map( A => n153, Z => n156);
   U50 : BUF_X1 port map( A => n161, Z => n164);
   U51 : NOR3_X1 port map( A1 => n169, A2 => S(2), A3 => n170, ZN => n11);
   U52 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n170, ZN => n12);
   U53 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n169, ZN => n13);
   U54 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => S(0), ZN => n14);
   U55 : AND3_X1 port map( A1 => S(0), A2 => n170, A3 => S(2), ZN => n9);
   U56 : AND3_X1 port map( A1 => n169, A2 => n170, A3 => S(2), ZN => n10);
   U57 : AND3_X1 port map( A1 => S(1), A2 => S(0), A3 => S(2), ZN => n7);
   U58 : AND3_X1 port map( A1 => S(1), A2 => n169, A3 => S(2), ZN => n8);
   U59 : AOI22_X1 port map( A1 => F(17), A2 => n158, B1 => E(17), B2 => n154, 
                           ZN => n105);
   U60 : AOI22_X1 port map( A1 => F(18), A2 => n158, B1 => E(18), B2 => n154, 
                           ZN => n101);
   U61 : AOI22_X1 port map( A1 => F(19), A2 => n158, B1 => E(19), B2 => n154, 
                           ZN => n97);
   U62 : AOI22_X1 port map( A1 => F(20), A2 => n159, B1 => E(20), B2 => n155, 
                           ZN => n89);
   U63 : AOI22_X1 port map( A1 => F(21), A2 => n159, B1 => E(21), B2 => n155, 
                           ZN => n85);
   U64 : AOI22_X1 port map( A1 => F(22), A2 => n159, B1 => E(22), B2 => n155, 
                           ZN => n81);
   U65 : AOI22_X1 port map( A1 => F(23), A2 => n159, B1 => E(23), B2 => n155, 
                           ZN => n77);
   U66 : AOI22_X1 port map( A1 => F(24), A2 => n159, B1 => E(24), B2 => n155, 
                           ZN => n73);
   U67 : AOI22_X1 port map( A1 => F(25), A2 => n159, B1 => E(25), B2 => n155, 
                           ZN => n69);
   U68 : AOI22_X1 port map( A1 => F(26), A2 => n159, B1 => E(26), B2 => n155, 
                           ZN => n65);
   U69 : AOI22_X1 port map( A1 => F(27), A2 => n159, B1 => E(27), B2 => n155, 
                           ZN => n61);
   U70 : AOI22_X1 port map( A1 => F(28), A2 => n159, B1 => E(28), B2 => n155, 
                           ZN => n57);
   U71 : AOI22_X1 port map( A1 => F(29), A2 => n159, B1 => E(29), B2 => n155, 
                           ZN => n53);
   U72 : AOI22_X1 port map( A1 => F(30), A2 => n159, B1 => E(30), B2 => n155, 
                           ZN => n45);
   U73 : AOI22_X1 port map( A1 => F(31), A2 => n160, B1 => E(31), B2 => n156, 
                           ZN => n41);
   U74 : NAND4_X1 port map( A1 => n135, A2 => n136, A3 => n137, A4 => n138, ZN 
                           => Y(0));
   U75 : AOI22_X1 port map( A1 => F(0), A2 => n158, B1 => E(0), B2 => n154, ZN 
                           => n137);
   U76 : AOI22_X1 port map( A1 => H(0), A2 => n166, B1 => G(0), B2 => n162, ZN 
                           => n138);
   U77 : AOI22_X1 port map( A1 => B(0), A2 => n141, B1 => A(0), B2 => n1, ZN =>
                           n135);
   U78 : NAND4_X1 port map( A1 => n51, A2 => n52, A3 => n53, A4 => n54, ZN => 
                           Y(29));
   U79 : AOI22_X1 port map( A1 => H(29), A2 => n167, B1 => G(29), B2 => n163, 
                           ZN => n54);
   U80 : AOI22_X1 port map( A1 => B(29), A2 => n142, B1 => A(29), B2 => n2, ZN 
                           => n51);
   U81 : AOI22_X1 port map( A1 => D(29), A2 => n150, B1 => C(29), B2 => n146, 
                           ZN => n52);
   U82 : NAND4_X1 port map( A1 => n103, A2 => n104, A3 => n105, A4 => n106, ZN 
                           => Y(17));
   U83 : AOI22_X1 port map( A1 => H(17), A2 => n166, B1 => G(17), B2 => n162, 
                           ZN => n106);
   U84 : AOI22_X1 port map( A1 => B(17), A2 => n141, B1 => A(17), B2 => n1, ZN 
                           => n103);
   U85 : AOI22_X1 port map( A1 => D(17), A2 => n149, B1 => C(17), B2 => n145, 
                           ZN => n104);
   U86 : NAND4_X1 port map( A1 => n99, A2 => n100, A3 => n101, A4 => n102, ZN 
                           => Y(18));
   U87 : AOI22_X1 port map( A1 => H(18), A2 => n166, B1 => G(18), B2 => n162, 
                           ZN => n102);
   U88 : AOI22_X1 port map( A1 => B(18), A2 => n141, B1 => A(18), B2 => n1, ZN 
                           => n99);
   U89 : AOI22_X1 port map( A1 => D(18), A2 => n149, B1 => C(18), B2 => n145, 
                           ZN => n100);
   U90 : NAND4_X1 port map( A1 => n95, A2 => n96, A3 => n97, A4 => n98, ZN => 
                           Y(19));
   U91 : AOI22_X1 port map( A1 => H(19), A2 => n166, B1 => G(19), B2 => n162, 
                           ZN => n98);
   U92 : AOI22_X1 port map( A1 => B(19), A2 => n141, B1 => A(19), B2 => n1, ZN 
                           => n95);
   U93 : AOI22_X1 port map( A1 => D(19), A2 => n149, B1 => C(19), B2 => n145, 
                           ZN => n96);
   U94 : NAND4_X1 port map( A1 => n87, A2 => n88, A3 => n89, A4 => n90, ZN => 
                           Y(20));
   U95 : AOI22_X1 port map( A1 => H(20), A2 => n167, B1 => G(20), B2 => n163, 
                           ZN => n90);
   U96 : AOI22_X1 port map( A1 => B(20), A2 => n142, B1 => A(20), B2 => n2, ZN 
                           => n87);
   U97 : AOI22_X1 port map( A1 => D(20), A2 => n150, B1 => C(20), B2 => n146, 
                           ZN => n88);
   U98 : NAND4_X1 port map( A1 => n83, A2 => n84, A3 => n85, A4 => n86, ZN => 
                           Y(21));
   U99 : AOI22_X1 port map( A1 => H(21), A2 => n167, B1 => G(21), B2 => n163, 
                           ZN => n86);
   U100 : AOI22_X1 port map( A1 => B(21), A2 => n142, B1 => A(21), B2 => n2, ZN
                           => n83);
   U101 : AOI22_X1 port map( A1 => D(21), A2 => n150, B1 => C(21), B2 => n146, 
                           ZN => n84);
   U102 : NAND4_X1 port map( A1 => n79, A2 => n80, A3 => n81, A4 => n82, ZN => 
                           Y(22));
   U103 : AOI22_X1 port map( A1 => H(22), A2 => n167, B1 => G(22), B2 => n163, 
                           ZN => n82);
   U104 : AOI22_X1 port map( A1 => B(22), A2 => n142, B1 => A(22), B2 => n2, ZN
                           => n79);
   U105 : AOI22_X1 port map( A1 => D(22), A2 => n150, B1 => C(22), B2 => n146, 
                           ZN => n80);
   U106 : NAND4_X1 port map( A1 => n75, A2 => n76, A3 => n77, A4 => n78, ZN => 
                           Y(23));
   U107 : AOI22_X1 port map( A1 => H(23), A2 => n167, B1 => G(23), B2 => n163, 
                           ZN => n78);
   U108 : AOI22_X1 port map( A1 => B(23), A2 => n142, B1 => A(23), B2 => n2, ZN
                           => n75);
   U109 : AOI22_X1 port map( A1 => D(23), A2 => n150, B1 => C(23), B2 => n146, 
                           ZN => n76);
   U110 : NAND4_X1 port map( A1 => n71, A2 => n72, A3 => n73, A4 => n74, ZN => 
                           Y(24));
   U111 : AOI22_X1 port map( A1 => H(24), A2 => n167, B1 => G(24), B2 => n163, 
                           ZN => n74);
   U112 : AOI22_X1 port map( A1 => B(24), A2 => n142, B1 => A(24), B2 => n2, ZN
                           => n71);
   U113 : AOI22_X1 port map( A1 => D(24), A2 => n150, B1 => C(24), B2 => n146, 
                           ZN => n72);
   U114 : NAND4_X1 port map( A1 => n67, A2 => n68, A3 => n69, A4 => n70, ZN => 
                           Y(25));
   U115 : AOI22_X1 port map( A1 => H(25), A2 => n167, B1 => G(25), B2 => n163, 
                           ZN => n70);
   U116 : AOI22_X1 port map( A1 => B(25), A2 => n142, B1 => A(25), B2 => n2, ZN
                           => n67);
   U117 : AOI22_X1 port map( A1 => D(25), A2 => n150, B1 => C(25), B2 => n146, 
                           ZN => n68);
   U118 : NAND4_X1 port map( A1 => n63, A2 => n64, A3 => n65, A4 => n66, ZN => 
                           Y(26));
   U119 : AOI22_X1 port map( A1 => H(26), A2 => n167, B1 => G(26), B2 => n163, 
                           ZN => n66);
   U120 : AOI22_X1 port map( A1 => B(26), A2 => n142, B1 => A(26), B2 => n2, ZN
                           => n63);
   U121 : AOI22_X1 port map( A1 => D(26), A2 => n150, B1 => C(26), B2 => n146, 
                           ZN => n64);
   U122 : NAND4_X1 port map( A1 => n59, A2 => n60, A3 => n61, A4 => n62, ZN => 
                           Y(27));
   U123 : AOI22_X1 port map( A1 => H(27), A2 => n167, B1 => G(27), B2 => n163, 
                           ZN => n62);
   U124 : AOI22_X1 port map( A1 => B(27), A2 => n142, B1 => A(27), B2 => n2, ZN
                           => n59);
   U125 : AOI22_X1 port map( A1 => D(27), A2 => n150, B1 => C(27), B2 => n146, 
                           ZN => n60);
   U126 : NAND4_X1 port map( A1 => n55, A2 => n56, A3 => n57, A4 => n58, ZN => 
                           Y(28));
   U127 : AOI22_X1 port map( A1 => H(28), A2 => n167, B1 => G(28), B2 => n163, 
                           ZN => n58);
   U128 : AOI22_X1 port map( A1 => B(28), A2 => n142, B1 => A(28), B2 => n2, ZN
                           => n55);
   U129 : AOI22_X1 port map( A1 => D(28), A2 => n150, B1 => C(28), B2 => n146, 
                           ZN => n56);
   U130 : NAND4_X1 port map( A1 => n43, A2 => n44, A3 => n45, A4 => n46, ZN => 
                           Y(30));
   U131 : AOI22_X1 port map( A1 => H(30), A2 => n167, B1 => G(30), B2 => n163, 
                           ZN => n46);
   U132 : AOI22_X1 port map( A1 => B(30), A2 => n142, B1 => A(30), B2 => n2, ZN
                           => n43);
   U133 : AOI22_X1 port map( A1 => D(30), A2 => n150, B1 => C(30), B2 => n146, 
                           ZN => n44);
   U134 : NAND4_X1 port map( A1 => n39, A2 => n40, A3 => n41, A4 => n42, ZN => 
                           Y(31));
   U135 : AOI22_X1 port map( A1 => H(31), A2 => n168, B1 => G(31), B2 => n164, 
                           ZN => n42);
   U136 : AOI22_X1 port map( A1 => B(31), A2 => n143, B1 => A(31), B2 => n139, 
                           ZN => n39);
   U137 : AOI22_X1 port map( A1 => D(31), A2 => n151, B1 => C(31), B2 => n147, 
                           ZN => n40);
   U138 : AOI22_X1 port map( A1 => D(0), A2 => n149, B1 => C(0), B2 => n145, ZN
                           => n136);
   U139 : NAND4_X1 port map( A1 => n91, A2 => n92, A3 => n93, A4 => n94, ZN => 
                           Y(1));
   U140 : AOI22_X1 port map( A1 => H(1), A2 => n166, B1 => G(1), B2 => n162, ZN
                           => n94);
   U141 : AOI22_X1 port map( A1 => B(1), A2 => n141, B1 => A(1), B2 => n1, ZN 
                           => n91);
   U142 : AOI22_X1 port map( A1 => F(1), A2 => n158, B1 => E(1), B2 => n154, ZN
                           => n93);
   U143 : NAND4_X1 port map( A1 => n47, A2 => n48, A3 => n49, A4 => n50, ZN => 
                           Y(2));
   U144 : AOI22_X1 port map( A1 => H(2), A2 => n167, B1 => G(2), B2 => n163, ZN
                           => n50);
   U145 : AOI22_X1 port map( A1 => B(2), A2 => n142, B1 => A(2), B2 => n2, ZN 
                           => n47);
   U146 : AOI22_X1 port map( A1 => F(2), A2 => n159, B1 => E(2), B2 => n155, ZN
                           => n49);
   U147 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           Y(3));
   U148 : AOI22_X1 port map( A1 => H(3), A2 => n168, B1 => G(3), B2 => n164, ZN
                           => n38);
   U149 : AOI22_X1 port map( A1 => B(3), A2 => n143, B1 => A(3), B2 => n139, ZN
                           => n35);
   U150 : AOI22_X1 port map( A1 => F(3), A2 => n160, B1 => E(3), B2 => n156, ZN
                           => n37);
   U151 : NAND4_X1 port map( A1 => n31, A2 => n32, A3 => n33, A4 => n34, ZN => 
                           Y(4));
   U152 : AOI22_X1 port map( A1 => H(4), A2 => n168, B1 => G(4), B2 => n164, ZN
                           => n34);
   U153 : AOI22_X1 port map( A1 => B(4), A2 => n143, B1 => A(4), B2 => n139, ZN
                           => n31);
   U154 : AOI22_X1 port map( A1 => F(4), A2 => n160, B1 => E(4), B2 => n156, ZN
                           => n33);
   U155 : NAND4_X1 port map( A1 => n27, A2 => n28, A3 => n29, A4 => n30, ZN => 
                           Y(5));
   U156 : AOI22_X1 port map( A1 => H(5), A2 => n168, B1 => G(5), B2 => n164, ZN
                           => n30);
   U157 : AOI22_X1 port map( A1 => B(5), A2 => n143, B1 => A(5), B2 => n139, ZN
                           => n27);
   U158 : AOI22_X1 port map( A1 => F(5), A2 => n160, B1 => E(5), B2 => n156, ZN
                           => n29);
   U159 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           Y(6));
   U160 : AOI22_X1 port map( A1 => H(6), A2 => n168, B1 => G(6), B2 => n164, ZN
                           => n26);
   U161 : AOI22_X1 port map( A1 => B(6), A2 => n143, B1 => A(6), B2 => n139, ZN
                           => n23);
   U162 : AOI22_X1 port map( A1 => F(6), A2 => n160, B1 => E(6), B2 => n156, ZN
                           => n25);
   U163 : NAND4_X1 port map( A1 => n19, A2 => n20, A3 => n21, A4 => n22, ZN => 
                           Y(7));
   U164 : AOI22_X1 port map( A1 => H(7), A2 => n168, B1 => G(7), B2 => n164, ZN
                           => n22);
   U165 : AOI22_X1 port map( A1 => B(7), A2 => n143, B1 => A(7), B2 => n139, ZN
                           => n19);
   U166 : AOI22_X1 port map( A1 => F(7), A2 => n160, B1 => E(7), B2 => n156, ZN
                           => n21);
   U167 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           Y(8));
   U168 : AOI22_X1 port map( A1 => H(8), A2 => n168, B1 => G(8), B2 => n164, ZN
                           => n18);
   U169 : AOI22_X1 port map( A1 => B(8), A2 => n143, B1 => A(8), B2 => n139, ZN
                           => n15);
   U170 : AOI22_X1 port map( A1 => F(8), A2 => n160, B1 => E(8), B2 => n156, ZN
                           => n17);
   U171 : NAND4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => Y(9)
                           );
   U172 : AOI22_X1 port map( A1 => H(9), A2 => n168, B1 => G(9), B2 => n164, ZN
                           => n6);
   U173 : AOI22_X1 port map( A1 => B(9), A2 => n143, B1 => A(9), B2 => n139, ZN
                           => n3);
   U174 : AOI22_X1 port map( A1 => F(9), A2 => n160, B1 => E(9), B2 => n156, ZN
                           => n5);
   U175 : NAND4_X1 port map( A1 => n131, A2 => n132, A3 => n133, A4 => n134, ZN
                           => Y(10));
   U176 : AOI22_X1 port map( A1 => H(10), A2 => n166, B1 => G(10), B2 => n162, 
                           ZN => n134);
   U177 : AOI22_X1 port map( A1 => B(10), A2 => n141, B1 => A(10), B2 => n1, ZN
                           => n131);
   U178 : AOI22_X1 port map( A1 => F(10), A2 => n158, B1 => E(10), B2 => n154, 
                           ZN => n133);
   U179 : NAND4_X1 port map( A1 => n127, A2 => n128, A3 => n129, A4 => n130, ZN
                           => Y(11));
   U180 : AOI22_X1 port map( A1 => H(11), A2 => n166, B1 => G(11), B2 => n162, 
                           ZN => n130);
   U181 : AOI22_X1 port map( A1 => B(11), A2 => n141, B1 => A(11), B2 => n1, ZN
                           => n127);
   U182 : AOI22_X1 port map( A1 => F(11), A2 => n158, B1 => E(11), B2 => n154, 
                           ZN => n129);
   U183 : NAND4_X1 port map( A1 => n123, A2 => n124, A3 => n125, A4 => n126, ZN
                           => Y(12));
   U184 : AOI22_X1 port map( A1 => H(12), A2 => n166, B1 => G(12), B2 => n162, 
                           ZN => n126);
   U185 : AOI22_X1 port map( A1 => B(12), A2 => n141, B1 => A(12), B2 => n1, ZN
                           => n123);
   U186 : AOI22_X1 port map( A1 => F(12), A2 => n158, B1 => E(12), B2 => n154, 
                           ZN => n125);
   U187 : NAND4_X1 port map( A1 => n119, A2 => n120, A3 => n121, A4 => n122, ZN
                           => Y(13));
   U188 : AOI22_X1 port map( A1 => H(13), A2 => n166, B1 => G(13), B2 => n162, 
                           ZN => n122);
   U189 : AOI22_X1 port map( A1 => B(13), A2 => n141, B1 => A(13), B2 => n1, ZN
                           => n119);
   U190 : AOI22_X1 port map( A1 => F(13), A2 => n158, B1 => E(13), B2 => n154, 
                           ZN => n121);
   U191 : NAND4_X1 port map( A1 => n115, A2 => n116, A3 => n117, A4 => n118, ZN
                           => Y(14));
   U192 : AOI22_X1 port map( A1 => H(14), A2 => n166, B1 => G(14), B2 => n162, 
                           ZN => n118);
   U193 : AOI22_X1 port map( A1 => B(14), A2 => n141, B1 => A(14), B2 => n1, ZN
                           => n115);
   U194 : AOI22_X1 port map( A1 => F(14), A2 => n158, B1 => E(14), B2 => n154, 
                           ZN => n117);
   U195 : NAND4_X1 port map( A1 => n111, A2 => n112, A3 => n113, A4 => n114, ZN
                           => Y(15));
   U196 : AOI22_X1 port map( A1 => H(15), A2 => n166, B1 => G(15), B2 => n162, 
                           ZN => n114);
   U197 : AOI22_X1 port map( A1 => B(15), A2 => n141, B1 => A(15), B2 => n1, ZN
                           => n111);
   U198 : AOI22_X1 port map( A1 => F(15), A2 => n158, B1 => E(15), B2 => n154, 
                           ZN => n113);
   U199 : NAND4_X1 port map( A1 => n107, A2 => n108, A3 => n109, A4 => n110, ZN
                           => Y(16));
   U200 : AOI22_X1 port map( A1 => H(16), A2 => n166, B1 => G(16), B2 => n162, 
                           ZN => n110);
   U201 : AOI22_X1 port map( A1 => B(16), A2 => n141, B1 => A(16), B2 => n1, ZN
                           => n107);
   U202 : AOI22_X1 port map( A1 => F(16), A2 => n158, B1 => E(16), B2 => n154, 
                           ZN => n109);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BOOTH_ENCODER_N16 is

   port( B : in std_logic_vector (15 downto 0);  Bo : out std_logic_vector (23 
         downto 0));

end BOOTH_ENCODER_N16;

architecture SYN_STRUCTURAL of BOOTH_ENCODER_N16 is

   component ENCODER_0
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_1
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_2
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_3
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_4
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_5
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_6
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_7
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   ENC_0 : ENCODER_7 port map( B(2) => B(1), B(1) => B(0), B(0) => 
                           X_Logic0_port, Y(2) => Bo(2), Y(1) => Bo(1), Y(0) =>
                           Bo(0));
   ENC_1 : ENCODER_6 port map( B(2) => B(3), B(1) => B(2), B(0) => B(1), Y(2) 
                           => Bo(5), Y(1) => Bo(4), Y(0) => Bo(3));
   ENC_2 : ENCODER_5 port map( B(2) => B(5), B(1) => B(4), B(0) => B(3), Y(2) 
                           => Bo(8), Y(1) => Bo(7), Y(0) => Bo(6));
   ENC_3 : ENCODER_4 port map( B(2) => B(7), B(1) => B(6), B(0) => B(5), Y(2) 
                           => Bo(11), Y(1) => Bo(10), Y(0) => Bo(9));
   ENC_4 : ENCODER_3 port map( B(2) => B(9), B(1) => B(8), B(0) => B(7), Y(2) 
                           => Bo(14), Y(1) => Bo(13), Y(0) => Bo(12));
   ENC_5 : ENCODER_2 port map( B(2) => B(11), B(1) => B(10), B(0) => B(9), Y(2)
                           => Bo(17), Y(1) => Bo(16), Y(0) => Bo(15));
   ENC_6 : ENCODER_1 port map( B(2) => B(13), B(1) => B(12), B(0) => B(11), 
                           Y(2) => Bo(20), Y(1) => Bo(19), Y(0) => Bo(18));
   ENC_7 : ENCODER_0 port map( B(2) => B(15), B(1) => B(14), B(0) => B(13), 
                           Y(2) => Bo(23), Y(1) => Bo(22), Y(0) => Bo(21));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GENERATOR_N32_NB8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_N32_NB8;

architecture SYN_STRUCTURAL of SUM_GENERATOR_N32_NB8 is

   component CSB_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_1 : CSB_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => Ci(0), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   CSBI_2 : CSB_N4_6 port map( A(3) => A(7), A(2) => A(6), A(1) => A(5), A(0) 
                           => A(4), B(3) => B(7), B(2) => B(6), B(1) => B(5), 
                           B(0) => B(4), Ci => Ci(1), S(3) => S(7), S(2) => 
                           S(6), S(1) => S(5), S(0) => S(4));
   CSBI_3 : CSB_N4_5 port map( A(3) => A(11), A(2) => A(10), A(1) => A(9), A(0)
                           => A(8), B(3) => B(11), B(2) => B(10), B(1) => B(9),
                           B(0) => B(8), Ci => Ci(2), S(3) => S(11), S(2) => 
                           S(10), S(1) => S(9), S(0) => S(8));
   CSBI_4 : CSB_N4_4 port map( A(3) => A(15), A(2) => A(14), A(1) => A(13), 
                           A(0) => A(12), B(3) => B(15), B(2) => B(14), B(1) =>
                           B(13), B(0) => B(12), Ci => Ci(3), S(3) => S(15), 
                           S(2) => S(14), S(1) => S(13), S(0) => S(12));
   CSBI_5 : CSB_N4_3 port map( A(3) => A(19), A(2) => A(18), A(1) => A(17), 
                           A(0) => A(16), B(3) => B(19), B(2) => B(18), B(1) =>
                           B(17), B(0) => B(16), Ci => Ci(4), S(3) => S(19), 
                           S(2) => S(18), S(1) => S(17), S(0) => S(16));
   CSBI_6 : CSB_N4_2 port map( A(3) => A(23), A(2) => A(22), A(1) => A(21), 
                           A(0) => A(20), B(3) => B(23), B(2) => B(22), B(1) =>
                           B(21), B(0) => B(20), Ci => Ci(5), S(3) => S(23), 
                           S(2) => S(22), S(1) => S(21), S(0) => S(20));
   CSBI_7 : CSB_N4_1 port map( A(3) => A(27), A(2) => A(26), A(1) => A(25), 
                           A(0) => A(24), B(3) => B(27), B(2) => B(26), B(1) =>
                           B(25), B(0) => B(24), Ci => Ci(6), S(3) => S(27), 
                           S(2) => S(26), S(1) => S(25), S(0) => S(24));
   CSBI_8 : CSB_N4_0 port map( A(3) => A(31), A(2) => A(30), A(1) => A(29), 
                           A(0) => A(28), B(3) => B(31), B(2) => B(30), B(1) =>
                           B(29), B(0) => B(28), Ci => Ci(7), S(3) => S(31), 
                           S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_N32_NB8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_N32_NB8;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_N32_NB8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component PG_BLOCK_0
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_0
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_1
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_1
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_2
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_2
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_3
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_3
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_4
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_5
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_6
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_4
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_7
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_5
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_8
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_9
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_10
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_11
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_6
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_12
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_13
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_14
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_15
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_16
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_17
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_18
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_7
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_19
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_20
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_21
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_22
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_23
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_24
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_25
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_26
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_27
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_28
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_29
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_30
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_31
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_32
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_33
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_8
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_ROW_N32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  P, G
            : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port,
      Co_2_port, Co_1_port, Co_0_port, G_4_31_port, G_4_27_port, G_4_23_port, 
      G_3_31_port, G_3_27_port, G_3_19_port, G_3_15_port, G_3_11_port, 
      G_2_31_port, G_2_23_port, G_2_15_port, G_2_7_port, G_1_31_port, 
      G_1_29_port, G_1_27_port, G_1_25_port, G_1_23_port, G_1_21_port, 
      G_1_19_port, G_1_17_port, G_1_15_port, G_1_13_port, G_1_11_port, 
      G_1_9_port, G_1_7_port, G_1_5_port, G_1_3_port, G_1_1_port, G_0_31_port, 
      G_0_30_port, G_0_29_port, G_0_28_port, G_0_27_port, G_0_26_port, 
      G_0_25_port, G_0_24_port, G_0_23_port, G_0_22_port, G_0_21_port, 
      G_0_20_port, G_0_19_port, G_0_18_port, G_0_17_port, G_0_16_port, 
      G_0_15_port, G_0_14_port, G_0_13_port, G_0_12_port, G_0_11_port, 
      G_0_10_port, G_0_9_port, G_0_8_port, G_0_7_port, G_0_6_port, G_0_5_port, 
      G_0_4_port, G_0_3_port, G_0_2_port, G_0_1_port, G_0_0_port, P_5_15_port, 
      P_4_31_port, P_4_27_port, P_4_23_port, P_4_7_port, P_3_31_port, 
      P_3_27_port, P_3_19_port, P_3_15_port, P_3_11_port, P_2_31_port, 
      P_2_23_port, P_2_15_port, P_2_7_port, P_1_31_port, P_1_29_port, 
      P_1_27_port, P_1_25_port, P_1_23_port, P_1_21_port, P_1_19_port, 
      P_1_17_port, P_1_15_port, P_1_13_port, P_1_11_port, P_1_9_port, 
      P_1_7_port, P_1_5_port, P_1_3_port, P_0_31_port, P_0_30_port, P_0_29_port
      , P_0_28_port, P_0_27_port, P_0_26_port, P_0_25_port, P_0_24_port, 
      P_0_23_port, P_0_22_port, P_0_21_port, P_0_20_port, P_0_19_port, 
      P_0_18_port, P_0_17_port, P_0_16_port, P_0_15_port, P_0_14_port, 
      P_0_13_port, P_0_12_port, P_0_11_port, P_0_10_port, P_0_9_port, 
      P_0_8_port, P_0_7_port, P_0_6_port, P_0_5_port, P_0_4_port, P_0_3_port, 
      P_0_2_port, P_0_1_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12
      , n13, n14, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   X_Logic0_port <= '0';
   PG_ROW_INSTANCE : PG_ROW_N32 port map( A(31) => A(31), A(30) => A(30), A(29)
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => Ci, P(31) => P_0_31_port, P(30) => 
                           P_0_30_port, P(29) => P_0_29_port, P(28) => 
                           P_0_28_port, P(27) => P_0_27_port, P(26) => 
                           P_0_26_port, P(25) => P_0_25_port, P(24) => 
                           P_0_24_port, P(23) => P_0_23_port, P(22) => 
                           P_0_22_port, P(21) => P_0_21_port, P(20) => 
                           P_0_20_port, P(19) => P_0_19_port, P(18) => 
                           P_0_18_port, P(17) => P_0_17_port, P(16) => 
                           P_0_16_port, P(15) => P_0_15_port, P(14) => 
                           P_0_14_port, P(13) => P_0_13_port, P(12) => 
                           P_0_12_port, P(11) => P_0_11_port, P(10) => 
                           P_0_10_port, P(9) => P_0_9_port, P(8) => P_0_8_port,
                           P(7) => P_0_7_port, P(6) => P_0_6_port, P(5) => 
                           P_0_5_port, P(4) => P_0_4_port, P(3) => P_0_3_port, 
                           P(2) => P_0_2_port, P(1) => P_0_1_port, P(0) => 
                           n_1250, G(31) => G_0_31_port, G(30) => G_0_30_port, 
                           G(29) => G_0_29_port, G(28) => G_0_28_port, G(27) =>
                           G_0_27_port, G(26) => G_0_26_port, G(25) => 
                           G_0_25_port, G(24) => G_0_24_port, G(23) => 
                           G_0_23_port, G(22) => G_0_22_port, G(21) => 
                           G_0_21_port, G(20) => G_0_20_port, G(19) => 
                           G_0_19_port, G(18) => G_0_18_port, G(17) => 
                           G_0_17_port, G(16) => G_0_16_port, G(15) => 
                           G_0_15_port, G(14) => G_0_14_port, G(13) => 
                           G_0_13_port, G(12) => G_0_12_port, G(11) => 
                           G_0_11_port, G(10) => G_0_10_port, G(9) => 
                           G_0_9_port, G(8) => G_0_8_port, G(7) => G_0_7_port, 
                           G(6) => G_0_6_port, G(5) => G_0_5_port, G(4) => 
                           G_0_4_port, G(3) => G_0_3_port, G(2) => G_0_2_port, 
                           G(1) => G_0_1_port, G(0) => G_0_0_port);
   G_BLOCK_INSTANCE_1_1 : GENERATE_BLOCK_8 port map( Gik => G_0_1_port, Gkj => 
                           G_0_0_port, Pik => P_0_1_port, Gij => G_1_1_port);
   PG_BLOCK_REG_INSTANCE_1_3 : PG_BLOCK_33 port map( Gik => G_0_3_port, Gkj => 
                           G_0_2_port, Pik => P_0_3_port, Pkj => P_0_2_port, 
                           Gij => G_1_3_port, Pij => P_1_3_port);
   PG_BLOCK_REG_INSTANCE_1_5 : PG_BLOCK_32 port map( Gik => G_0_5_port, Gkj => 
                           G_0_4_port, Pik => P_0_5_port, Pkj => P_0_4_port, 
                           Gij => G_1_5_port, Pij => P_1_5_port);
   PG_BLOCK_REG_INSTANCE_1_7 : PG_BLOCK_31 port map( Gik => G_0_7_port, Gkj => 
                           G_0_6_port, Pik => P_0_7_port, Pkj => P_0_6_port, 
                           Gij => G_1_7_port, Pij => P_1_7_port);
   PG_BLOCK_REG_INSTANCE_1_9 : PG_BLOCK_30 port map( Gik => G_0_9_port, Gkj => 
                           G_0_8_port, Pik => P_0_9_port, Pkj => P_0_8_port, 
                           Gij => G_1_9_port, Pij => P_1_9_port);
   PG_BLOCK_REG_INSTANCE_1_11 : PG_BLOCK_29 port map( Gik => G_0_11_port, Gkj 
                           => G_0_10_port, Pik => P_0_11_port, Pkj => 
                           P_0_10_port, Gij => G_1_11_port, Pij => P_1_11_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_13 : PG_BLOCK_28 port map( Gik => G_0_13_port, Gkj 
                           => G_0_12_port, Pik => P_0_13_port, Pkj => 
                           P_0_12_port, Gij => G_1_13_port, Pij => P_1_13_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_15 : PG_BLOCK_27 port map( Gik => G_0_15_port, Gkj 
                           => G_0_14_port, Pik => P_0_15_port, Pkj => 
                           P_0_14_port, Gij => G_1_15_port, Pij => P_1_15_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_17 : PG_BLOCK_26 port map( Gik => G_0_17_port, Gkj 
                           => G_0_16_port, Pik => P_0_17_port, Pkj => 
                           P_0_16_port, Gij => G_1_17_port, Pij => P_1_17_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_19 : PG_BLOCK_25 port map( Gik => G_0_19_port, Gkj 
                           => G_0_18_port, Pik => P_0_19_port, Pkj => 
                           P_0_18_port, Gij => G_1_19_port, Pij => P_1_19_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_21 : PG_BLOCK_24 port map( Gik => G_0_21_port, Gkj 
                           => G_0_20_port, Pik => P_0_21_port, Pkj => 
                           P_0_20_port, Gij => G_1_21_port, Pij => P_1_21_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_23 : PG_BLOCK_23 port map( Gik => G_0_23_port, Gkj 
                           => G_0_22_port, Pik => P_0_23_port, Pkj => 
                           P_0_22_port, Gij => G_1_23_port, Pij => P_1_23_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_25 : PG_BLOCK_22 port map( Gik => G_0_25_port, Gkj 
                           => G_0_24_port, Pik => P_0_25_port, Pkj => 
                           P_0_24_port, Gij => G_1_25_port, Pij => P_1_25_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_27 : PG_BLOCK_21 port map( Gik => G_0_27_port, Gkj 
                           => G_0_26_port, Pik => P_0_27_port, Pkj => 
                           P_0_26_port, Gij => G_1_27_port, Pij => P_1_27_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_29 : PG_BLOCK_20 port map( Gik => G_0_29_port, Gkj 
                           => G_0_28_port, Pik => P_0_29_port, Pkj => 
                           P_0_28_port, Gij => G_1_29_port, Pij => P_1_29_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_31 : PG_BLOCK_19 port map( Gik => G_0_31_port, Gkj 
                           => G_0_30_port, Pik => P_0_31_port, Pkj => 
                           P_0_30_port, Gij => G_1_31_port, Pij => P_1_31_port)
                           ;
   G_BLOCK_INSTANCE_2_3 : GENERATE_BLOCK_7 port map( Gik => G_1_3_port, Gkj => 
                           G_1_1_port, Pik => P_1_3_port, Gij => Co_0_port);
   PG_BLOCK_REG_INSTANCE_2_7 : PG_BLOCK_18 port map( Gik => G_1_7_port, Gkj => 
                           G_1_5_port, Pik => P_1_7_port, Pkj => P_1_5_port, 
                           Gij => G_2_7_port, Pij => P_2_7_port);
   PG_BLOCK_REG_INSTANCE_2_11 : PG_BLOCK_17 port map( Gik => G_1_11_port, Gkj 
                           => G_1_9_port, Pik => P_1_11_port, Pkj => P_1_9_port
                           , Gij => G_3_11_port, Pij => P_3_11_port);
   PG_BLOCK_REG_INSTANCE_2_15 : PG_BLOCK_16 port map( Gik => G_1_15_port, Gkj 
                           => G_1_13_port, Pik => P_1_15_port, Pkj => 
                           P_1_13_port, Gij => G_2_15_port, Pij => P_2_15_port)
                           ;
   PG_BLOCK_REG_INSTANCE_2_19 : PG_BLOCK_15 port map( Gik => G_1_19_port, Gkj 
                           => G_1_17_port, Pik => P_1_19_port, Pkj => 
                           P_1_17_port, Gij => G_3_19_port, Pij => P_3_19_port)
                           ;
   PG_BLOCK_REG_INSTANCE_2_23 : PG_BLOCK_14 port map( Gik => G_1_23_port, Gkj 
                           => G_1_21_port, Pik => P_1_23_port, Pkj => 
                           P_1_21_port, Gij => G_2_23_port, Pij => P_2_23_port)
                           ;
   PG_BLOCK_REG_INSTANCE_2_27 : PG_BLOCK_13 port map( Gik => G_1_27_port, Gkj 
                           => G_1_25_port, Pik => P_1_27_port, Pkj => 
                           P_1_25_port, Gij => G_3_27_port, Pij => P_3_27_port)
                           ;
   PG_BLOCK_REG_INSTANCE_2_31 : PG_BLOCK_12 port map( Gik => G_1_31_port, Gkj 
                           => G_1_29_port, Pik => P_1_31_port, Pkj => 
                           P_1_29_port, Gij => G_2_31_port, Pij => P_2_31_port)
                           ;
   G_BLOCK_INSTANCE_3_7 : GENERATE_BLOCK_6 port map( Gik => G_2_7_port, Gkj => 
                           Co_0_port, Pik => P_2_7_port, Gij => n1);
   PG_BLOCK_REG_INSTANCE_3_7 : PG_BLOCK_11 port map( Gik => G_2_7_port, Gkj => 
                           Co_0_port, Pik => P_2_7_port, Pkj => X_Logic0_port, 
                           Gij => n2, Pij => P_4_7_port);
   PG_BLOCK_REG_INSTANCE_3_15 : PG_BLOCK_10 port map( Gik => G_2_15_port, Gkj 
                           => G_3_11_port, Pik => P_2_15_port, Pkj => 
                           P_3_11_port, Gij => G_3_15_port, Pij => P_3_15_port)
                           ;
   PG_BLOCK_REG_INSTANCE_3_23 : PG_BLOCK_9 port map( Gik => G_2_23_port, Gkj =>
                           G_3_19_port, Pik => P_2_23_port, Pkj => P_3_19_port,
                           Gij => G_4_23_port, Pij => P_4_23_port);
   PG_BLOCK_REG_INSTANCE_3_31 : PG_BLOCK_8 port map( Gik => G_2_31_port, Gkj =>
                           G_3_27_port, Pik => P_2_31_port, Pkj => P_3_27_port,
                           Gij => G_3_31_port, Pij => P_3_31_port);
   G_BLOCK_INSTANCE_4_11 : GENERATE_BLOCK_5 port map( Gik => G_3_11_port, Gkj 
                           => Co_1_port, Pik => P_3_11_port, Gij => n3);
   PG_BLOCK_REG_INSTANCE_4_11 : PG_BLOCK_7 port map( Gik => G_3_11_port, Gkj =>
                           Co_1_port, Pik => P_3_11_port, Pkj => P_4_7_port, 
                           Gij => n4, Pij => n_1251);
   G_BLOCK_INSTANCE_4_15 : GENERATE_BLOCK_4 port map( Gik => G_3_15_port, Gkj 
                           => Co_1_port, Pik => P_3_15_port, Gij => n5);
   PG_BLOCK_REG_INSTANCE_4_15 : PG_BLOCK_6 port map( Gik => G_3_15_port, Gkj =>
                           Co_1_port, Pik => P_3_15_port, Pkj => P_4_7_port, 
                           Gij => n6, Pij => P_5_15_port);
   PG_BLOCK_REG_INSTANCE_4_27 : PG_BLOCK_5 port map( Gik => G_3_27_port, Gkj =>
                           G_4_23_port, Pik => P_3_27_port, Pkj => P_4_23_port,
                           Gij => G_4_27_port, Pij => P_4_27_port);
   PG_BLOCK_REG_INSTANCE_4_31 : PG_BLOCK_4 port map( Gik => G_3_31_port, Gkj =>
                           G_4_23_port, Pik => P_3_31_port, Pkj => P_4_23_port,
                           Gij => G_4_31_port, Pij => P_4_31_port);
   G_BLOCK_INSTANCE_5_19 : GENERATE_BLOCK_3 port map( Gik => G_3_19_port, Gkj 
                           => Co_3_port, Pik => P_3_19_port, Gij => n7);
   PG_BLOCK_REG_INSTANCE_5_19 : PG_BLOCK_3 port map( Gik => G_3_19_port, Gkj =>
                           Co_3_port, Pik => P_3_19_port, Pkj => P_5_15_port, 
                           Gij => n8, Pij => n_1252);
   G_BLOCK_INSTANCE_5_23 : GENERATE_BLOCK_2 port map( Gik => G_4_23_port, Gkj 
                           => Co_3_port, Pik => P_4_23_port, Gij => n9);
   PG_BLOCK_REG_INSTANCE_5_23 : PG_BLOCK_2 port map( Gik => G_4_23_port, Gkj =>
                           Co_3_port, Pik => P_4_23_port, Pkj => P_5_15_port, 
                           Gij => n10, Pij => n_1253);
   G_BLOCK_INSTANCE_5_27 : GENERATE_BLOCK_1 port map( Gik => G_4_27_port, Gkj 
                           => Co_3_port, Pik => P_4_27_port, Gij => n11);
   PG_BLOCK_REG_INSTANCE_5_27 : PG_BLOCK_1 port map( Gik => G_4_27_port, Gkj =>
                           Co_3_port, Pik => P_4_27_port, Pkj => P_5_15_port, 
                           Gij => n12, Pij => n_1254);
   G_BLOCK_INSTANCE_5_31 : GENERATE_BLOCK_0 port map( Gik => G_4_31_port, Gkj 
                           => Co_3_port, Pik => P_4_31_port, Gij => n13);
   PG_BLOCK_REG_INSTANCE_5_31 : PG_BLOCK_0 port map( Gik => G_4_31_port, Gkj =>
                           Co_3_port, Pik => P_4_31_port, Pkj => P_5_15_port, 
                           Gij => n14, Pij => n_1255);
   U2 : AND2_X1 port map( A1 => n5, A2 => n6, ZN => Co_3_port);
   U3 : AND2_X1 port map( A1 => n13, A2 => n14, ZN => Co_7_port);
   U4 : AND2_X1 port map( A1 => n11, A2 => n12, ZN => Co_6_port);
   U5 : AND2_X1 port map( A1 => n9, A2 => n10, ZN => Co_5_port);
   U6 : AND2_X1 port map( A1 => n7, A2 => n8, ZN => Co_4_port);
   U7 : AND2_X1 port map( A1 => n3, A2 => n4, ZN => Co_2_port);
   U8 : AND2_X1 port map( A1 => n1, A2 => n2, ZN => Co_1_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_61;

architecture SYN_BEHAVIORAL of AND2_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_63;

architecture SYN_BEHAVIORAL of XNOR2_63 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ZERO_DETECTOR_N32_0 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic);

end ZERO_DETECTOR_N32_0;

architecture SYN_STRUCTURAL of ZERO_DETECTOR_N32_0 is

   component AND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, M_4_1_port, M_4_0_port, M_3_3_port, M_3_2_port, 
      M_3_1_port, M_3_0_port, M_2_7_port, M_2_6_port, M_2_5_port, M_2_4_port, 
      M_2_3_port, M_2_2_port, M_2_1_port, M_2_0_port, M_1_15_port, M_1_14_port,
      M_1_13_port, M_1_12_port, M_1_11_port, M_1_10_port, M_1_9_port, 
      M_1_8_port, M_1_7_port, M_1_6_port, M_1_5_port, M_1_4_port, M_1_3_port, 
      M_1_2_port, M_1_1_port, M_1_0_port, M_0_31_port, M_0_30_port, M_0_29_port
      , M_0_28_port, M_0_27_port, M_0_26_port, M_0_25_port, M_0_24_port, 
      M_0_23_port, M_0_22_port, M_0_21_port, M_0_20_port, M_0_19_port, 
      M_0_18_port, M_0_17_port, M_0_16_port, M_0_15_port, M_0_14_port, 
      M_0_13_port, M_0_12_port, M_0_11_port, M_0_10_port, M_0_9_port, 
      M_0_8_port, M_0_7_port, M_0_6_port, M_0_5_port, M_0_4_port, M_0_3_port, 
      M_0_2_port, M_0_1_port, M_0_0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   XOR0_i_0_0 : XNOR2_31 port map( A => A(0), B => X_Logic0_port, Y => 
                           M_0_0_port);
   XOR0_i_0_1 : XNOR2_30 port map( A => A(1), B => X_Logic0_port, Y => 
                           M_0_1_port);
   XOR0_i_0_2 : XNOR2_29 port map( A => A(2), B => X_Logic0_port, Y => 
                           M_0_2_port);
   XOR0_i_0_3 : XNOR2_28 port map( A => A(3), B => X_Logic0_port, Y => 
                           M_0_3_port);
   XOR0_i_0_4 : XNOR2_27 port map( A => A(4), B => X_Logic0_port, Y => 
                           M_0_4_port);
   XOR0_i_0_5 : XNOR2_26 port map( A => A(5), B => X_Logic0_port, Y => 
                           M_0_5_port);
   XOR0_i_0_6 : XNOR2_25 port map( A => A(6), B => X_Logic0_port, Y => 
                           M_0_6_port);
   XOR0_i_0_7 : XNOR2_24 port map( A => A(7), B => X_Logic0_port, Y => 
                           M_0_7_port);
   XOR0_i_0_8 : XNOR2_23 port map( A => A(8), B => X_Logic0_port, Y => 
                           M_0_8_port);
   XOR0_i_0_9 : XNOR2_22 port map( A => A(9), B => X_Logic0_port, Y => 
                           M_0_9_port);
   XOR0_i_0_10 : XNOR2_21 port map( A => A(10), B => X_Logic0_port, Y => 
                           M_0_10_port);
   XOR0_i_0_11 : XNOR2_20 port map( A => A(11), B => X_Logic0_port, Y => 
                           M_0_11_port);
   XOR0_i_0_12 : XNOR2_19 port map( A => A(12), B => X_Logic0_port, Y => 
                           M_0_12_port);
   XOR0_i_0_13 : XNOR2_18 port map( A => A(13), B => X_Logic0_port, Y => 
                           M_0_13_port);
   XOR0_i_0_14 : XNOR2_17 port map( A => A(14), B => X_Logic0_port, Y => 
                           M_0_14_port);
   XOR0_i_0_15 : XNOR2_16 port map( A => A(15), B => X_Logic0_port, Y => 
                           M_0_15_port);
   XOR0_i_0_16 : XNOR2_15 port map( A => A(16), B => X_Logic0_port, Y => 
                           M_0_16_port);
   XOR0_i_0_17 : XNOR2_14 port map( A => A(17), B => X_Logic0_port, Y => 
                           M_0_17_port);
   XOR0_i_0_18 : XNOR2_13 port map( A => A(18), B => X_Logic0_port, Y => 
                           M_0_18_port);
   XOR0_i_0_19 : XNOR2_12 port map( A => A(19), B => X_Logic0_port, Y => 
                           M_0_19_port);
   XOR0_i_0_20 : XNOR2_11 port map( A => A(20), B => X_Logic0_port, Y => 
                           M_0_20_port);
   XOR0_i_0_21 : XNOR2_10 port map( A => A(21), B => X_Logic0_port, Y => 
                           M_0_21_port);
   XOR0_i_0_22 : XNOR2_9 port map( A => A(22), B => X_Logic0_port, Y => 
                           M_0_22_port);
   XOR0_i_0_23 : XNOR2_8 port map( A => A(23), B => X_Logic0_port, Y => 
                           M_0_23_port);
   XOR0_i_0_24 : XNOR2_7 port map( A => A(24), B => X_Logic0_port, Y => 
                           M_0_24_port);
   XOR0_i_0_25 : XNOR2_6 port map( A => A(25), B => X_Logic0_port, Y => 
                           M_0_25_port);
   XOR0_i_0_26 : XNOR2_5 port map( A => A(26), B => X_Logic0_port, Y => 
                           M_0_26_port);
   XOR0_i_0_27 : XNOR2_4 port map( A => A(27), B => X_Logic0_port, Y => 
                           M_0_27_port);
   XOR0_i_0_28 : XNOR2_3 port map( A => A(28), B => X_Logic0_port, Y => 
                           M_0_28_port);
   XOR0_i_0_29 : XNOR2_2 port map( A => A(29), B => X_Logic0_port, Y => 
                           M_0_29_port);
   XOR0_i_0_30 : XNOR2_1 port map( A => A(30), B => X_Logic0_port, Y => 
                           M_0_30_port);
   XOR0_i_0_31 : XNOR2_0 port map( A => A(31), B => X_Logic0_port, Y => 
                           M_0_31_port);
   AND_i_1_0 : AND2_30 port map( A => M_0_0_port, B => M_0_1_port, Y => 
                           M_1_0_port);
   AND_i_1_1 : AND2_29 port map( A => M_0_2_port, B => M_0_3_port, Y => 
                           M_1_1_port);
   AND_i_1_2 : AND2_28 port map( A => M_0_4_port, B => M_0_5_port, Y => 
                           M_1_2_port);
   AND_i_1_3 : AND2_27 port map( A => M_0_6_port, B => M_0_7_port, Y => 
                           M_1_3_port);
   AND_i_1_4 : AND2_26 port map( A => M_0_8_port, B => M_0_9_port, Y => 
                           M_1_4_port);
   AND_i_1_5 : AND2_25 port map( A => M_0_10_port, B => M_0_11_port, Y => 
                           M_1_5_port);
   AND_i_1_6 : AND2_24 port map( A => M_0_12_port, B => M_0_13_port, Y => 
                           M_1_6_port);
   AND_i_1_7 : AND2_23 port map( A => M_0_14_port, B => M_0_15_port, Y => 
                           M_1_7_port);
   AND_i_1_8 : AND2_22 port map( A => M_0_16_port, B => M_0_17_port, Y => 
                           M_1_8_port);
   AND_i_1_9 : AND2_21 port map( A => M_0_18_port, B => M_0_19_port, Y => 
                           M_1_9_port);
   AND_i_1_10 : AND2_20 port map( A => M_0_20_port, B => M_0_21_port, Y => 
                           M_1_10_port);
   AND_i_1_11 : AND2_19 port map( A => M_0_22_port, B => M_0_23_port, Y => 
                           M_1_11_port);
   AND_i_1_12 : AND2_18 port map( A => M_0_24_port, B => M_0_25_port, Y => 
                           M_1_12_port);
   AND_i_1_13 : AND2_17 port map( A => M_0_26_port, B => M_0_27_port, Y => 
                           M_1_13_port);
   AND_i_1_14 : AND2_16 port map( A => M_0_28_port, B => M_0_29_port, Y => 
                           M_1_14_port);
   AND_i_1_15 : AND2_15 port map( A => M_0_30_port, B => M_0_31_port, Y => 
                           M_1_15_port);
   AND_i_2_0 : AND2_14 port map( A => M_1_0_port, B => M_1_1_port, Y => 
                           M_2_0_port);
   AND_i_2_1 : AND2_13 port map( A => M_1_2_port, B => M_1_3_port, Y => 
                           M_2_1_port);
   AND_i_2_2 : AND2_12 port map( A => M_1_4_port, B => M_1_5_port, Y => 
                           M_2_2_port);
   AND_i_2_3 : AND2_11 port map( A => M_1_6_port, B => M_1_7_port, Y => 
                           M_2_3_port);
   AND_i_2_4 : AND2_10 port map( A => M_1_8_port, B => M_1_9_port, Y => 
                           M_2_4_port);
   AND_i_2_5 : AND2_9 port map( A => M_1_10_port, B => M_1_11_port, Y => 
                           M_2_5_port);
   AND_i_2_6 : AND2_8 port map( A => M_1_12_port, B => M_1_13_port, Y => 
                           M_2_6_port);
   AND_i_2_7 : AND2_7 port map( A => M_1_14_port, B => M_1_15_port, Y => 
                           M_2_7_port);
   AND_i_3_0 : AND2_6 port map( A => M_2_0_port, B => M_2_1_port, Y => 
                           M_3_0_port);
   AND_i_3_1 : AND2_5 port map( A => M_2_2_port, B => M_2_3_port, Y => 
                           M_3_1_port);
   AND_i_3_2 : AND2_4 port map( A => M_2_4_port, B => M_2_5_port, Y => 
                           M_3_2_port);
   AND_i_3_3 : AND2_3 port map( A => M_2_6_port, B => M_2_7_port, Y => 
                           M_3_3_port);
   AND_i_4_0 : AND2_2 port map( A => M_3_0_port, B => M_3_1_port, Y => 
                           M_4_0_port);
   AND_i_4_1 : AND2_1 port map( A => M_3_2_port, B => M_3_3_port, Y => 
                           M_4_1_port);
   AND_i_5_0 : AND2_0 port map( A => M_4_0_port, B => M_4_1_port, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity COMPARATOR_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic_vector (3 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end COMPARATOR_N32;

architecture SYN_BEHAVIORAL of COMPARATOR_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal X_Logic0_port, Y_0_port, N46, N47, N48, N49, N50, N51, N52, N53, N54,
      N55, n17, n18, n23, n24, n25, n26, n27, n28, n29, n30, n31, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20, n21,
      n22, n32, n33, n34, n35, n_1256, n_1257 : std_logic;

begin
   Y <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, Y_0_port );
   
   X_Logic0_port <= '0';
   n17 <= '1';
   n18 <= '0';
   r71 : COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4 port map( A(31) => A(31), A(30)
                           => A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => n22,
                           A(14) => n21, A(13) => n20, A(12) => n19, A(11) => 
                           n16, A(10) => n15, A(9) => n14, A(8) => n13, A(7) =>
                           n12, A(6) => n11, A(5) => n10, A(4) => n9, A(3) => 
                           n8, A(2) => n7, A(1) => A(1), A(0) => n6, B(31) => 
                           B(31), B(30) => B(30), B(29) => B(29), B(28) => 
                           B(28), B(27) => B(27), B(26) => B(26), B(25) => 
                           B(25), B(24) => B(24), B(23) => B(23), B(22) => 
                           B(22), B(21) => B(21), B(20) => B(20), B(19) => 
                           B(19), B(18) => B(18), B(17) => B(17), B(16) => 
                           B(16), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => n5, B(3) => n4, 
                           B(2) => n3, B(1) => n2, B(0) => n1, TC => n17, LT =>
                           N48, GT => N50, EQ => n_1256, LE => N52, GE => N54, 
                           NE => n_1257);
   r70 : COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5 port map( A(31) => A(31), A(30)
                           => A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => n22,
                           A(14) => n21, A(13) => n20, A(12) => n19, A(11) => 
                           n16, A(10) => n15, A(9) => n14, A(8) => n13, A(7) =>
                           n12, A(6) => n11, A(5) => n10, A(4) => n9, A(3) => 
                           n8, A(2) => n7, A(1) => A(1), A(0) => n6, B(31) => 
                           B(31), B(30) => B(30), B(29) => B(29), B(28) => 
                           B(28), B(27) => B(27), B(26) => B(26), B(25) => 
                           B(25), B(24) => B(24), B(23) => B(23), B(22) => 
                           B(22), B(21) => B(21), B(20) => B(20), B(19) => 
                           B(19), B(18) => B(18), B(17) => B(17), B(16) => 
                           B(16), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => n5, B(3) => n4, 
                           B(2) => n3, B(1) => n2, B(0) => n1, TC => n18, LT =>
                           N49, GT => N51, EQ => N46, LE => N53, GE => N55, NE 
                           => N47);
   U4 : BUF_X1 port map( A => B(3), Z => n4);
   U5 : BUF_X1 port map( A => B(1), Z => n2);
   U6 : BUF_X1 port map( A => B(0), Z => n1);
   U7 : BUF_X1 port map( A => A(2), Z => n7);
   U8 : BUF_X1 port map( A => A(6), Z => n11);
   U9 : BUF_X1 port map( A => A(10), Z => n15);
   U10 : BUF_X1 port map( A => A(0), Z => n6);
   U11 : BUF_X1 port map( A => A(14), Z => n21);
   U12 : BUF_X1 port map( A => B(4), Z => n5);
   U13 : BUF_X1 port map( A => B(2), Z => n3);
   U14 : BUF_X1 port map( A => A(4), Z => n9);
   U15 : BUF_X1 port map( A => A(5), Z => n10);
   U16 : BUF_X1 port map( A => A(8), Z => n13);
   U17 : BUF_X1 port map( A => A(9), Z => n14);
   U18 : BUF_X1 port map( A => A(12), Z => n19);
   U19 : BUF_X1 port map( A => A(13), Z => n20);
   U20 : BUF_X1 port map( A => A(3), Z => n8);
   U21 : BUF_X1 port map( A => A(7), Z => n12);
   U22 : BUF_X1 port map( A => A(11), Z => n16);
   U23 : BUF_X1 port map( A => A(15), Z => n22);
   U24 : OAI22_X1 port map( A1 => n28, A2 => n33, B1 => S(1), B2 => n29, ZN => 
                           n27);
   U25 : AOI22_X1 port map( A1 => N52, A2 => n35, B1 => N53, B2 => S(0), ZN => 
                           n28);
   U26 : AOI22_X1 port map( A1 => N50, A2 => n35, B1 => N51, B2 => S(0), ZN => 
                           n29);
   U27 : OAI22_X1 port map( A1 => n30, A2 => n33, B1 => S(1), B2 => n31, ZN => 
                           n26);
   U28 : AOI22_X1 port map( A1 => N48, A2 => n35, B1 => N49, B2 => S(0), ZN => 
                           n30);
   U29 : AOI22_X1 port map( A1 => N46, A2 => n35, B1 => N47, B2 => S(0), ZN => 
                           n31);
   U30 : INV_X1 port map( A => S(0), ZN => n35);
   U31 : AOI22_X1 port map( A1 => N54, A2 => n35, B1 => S(0), B2 => N55, ZN => 
                           n25);
   U32 : OAI21_X1 port map( B1 => S(3), B2 => n23, A => n24, ZN => Y_0_port);
   U33 : NAND4_X1 port map( A1 => n34, A2 => S(3), A3 => n32, A4 => n33, ZN => 
                           n24);
   U34 : AOI22_X1 port map( A1 => n26, A2 => n32, B1 => S(2), B2 => n27, ZN => 
                           n23);
   U35 : INV_X1 port map( A => n25, ZN => n34);
   U36 : INV_X1 port map( A => S(1), ZN => n33);
   U37 : INV_X1 port map( A => S(2), ZN => n32);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LOGIC_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic_vector (1 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end LOGIC_N32;

architecture SYN_BEHAVIORAL of LOGIC_N32 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n132, n133, n134, n135, n136, n137, n138, n139
      , n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => n69, Z => n11);
   U3 : BUF_X1 port map( A => n69, Z => n10);
   U4 : BUF_X1 port map( A => n20, Z => n19);
   U5 : BUF_X1 port map( A => n20, Z => n18);
   U6 : BUF_X1 port map( A => n11, Z => n4);
   U7 : BUF_X1 port map( A => n11, Z => n5);
   U8 : BUF_X1 port map( A => n10, Z => n8);
   U9 : BUF_X1 port map( A => n10, Z => n7);
   U10 : BUF_X1 port map( A => n11, Z => n6);
   U11 : BUF_X1 port map( A => n18, Z => n16);
   U12 : BUF_X1 port map( A => n18, Z => n15);
   U13 : BUF_X1 port map( A => n19, Z => n12);
   U14 : BUF_X1 port map( A => n19, Z => n13);
   U15 : BUF_X1 port map( A => n19, Z => n14);
   U16 : BUF_X1 port map( A => n18, Z => n17);
   U17 : BUF_X1 port map( A => n10, Z => n9);
   U18 : INV_X1 port map( A => n26, ZN => n27);
   U19 : INV_X1 port map( A => n28, ZN => n29);
   U20 : INV_X1 port map( A => n30, ZN => n31);
   U21 : INV_X1 port map( A => n32, ZN => n33);
   U22 : INV_X1 port map( A => n34, ZN => n35);
   U23 : INV_X1 port map( A => n36, ZN => n37);
   U24 : INV_X1 port map( A => n38, ZN => n39);
   U25 : INV_X1 port map( A => n40, ZN => n41);
   U26 : INV_X1 port map( A => n42, ZN => n43);
   U27 : INV_X1 port map( A => n44, ZN => n45);
   U28 : INV_X1 port map( A => n46, ZN => n47);
   U29 : INV_X1 port map( A => n48, ZN => n49);
   U30 : INV_X1 port map( A => n50, ZN => n51);
   U31 : INV_X1 port map( A => n52, ZN => n53);
   U32 : INV_X1 port map( A => n54, ZN => n55);
   U33 : INV_X1 port map( A => n56, ZN => n57);
   U34 : OAI22_X1 port map( A1 => n130, A2 => n21, B1 => n131, B2 => n27, ZN =>
                           Y(0));
   U35 : AOI21_X1 port map( B1 => n14, B2 => n21, A => n6, ZN => n131);
   U36 : AOI221_X1 port map( B1 => n26, B2 => n3, C1 => n12, C2 => n27, A => n4
                           , ZN => n130);
   U37 : INV_X1 port map( A => B(0), ZN => n21);
   U38 : OAI22_X1 port map( A1 => n108, A2 => n22, B1 => n109, B2 => n29, ZN =>
                           Y(1));
   U39 : AOI21_X1 port map( B1 => n16, B2 => n22, A => n8, ZN => n109);
   U40 : AOI221_X1 port map( B1 => n28, B2 => n2, C1 => n13, C2 => n29, A => n5
                           , ZN => n108);
   U41 : INV_X1 port map( A => B(1), ZN => n22);
   U42 : OAI22_X1 port map( A1 => n86, A2 => n23, B1 => n87, B2 => n31, ZN => 
                           Y(2));
   U43 : AOI21_X1 port map( B1 => n15, B2 => n23, A => n7, ZN => n87);
   U44 : AOI221_X1 port map( B1 => n30, B2 => n1, C1 => n14, C2 => n31, A => n6
                           , ZN => n86);
   U45 : INV_X1 port map( A => B(2), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n80, A2 => n24, B1 => n81, B2 => n33, ZN => 
                           Y(3));
   U47 : AOI21_X1 port map( B1 => n15, B2 => n24, A => n7, ZN => n81);
   U48 : AOI221_X1 port map( B1 => n32, B2 => n1, C1 => n13, C2 => n33, A => n5
                           , ZN => n80);
   U49 : INV_X1 port map( A => B(3), ZN => n24);
   U50 : OAI22_X1 port map( A1 => n78, A2 => n25, B1 => n79, B2 => n35, ZN => 
                           Y(4));
   U51 : AOI21_X1 port map( B1 => n15, B2 => n25, A => n7, ZN => n79);
   U52 : AOI221_X1 port map( B1 => n34, B2 => n1, C1 => n13, C2 => n35, A => n5
                           , ZN => n78);
   U53 : INV_X1 port map( A => B(4), ZN => n25);
   U54 : BUF_X1 port map( A => A(1), Z => n28);
   U55 : BUF_X1 port map( A => A(3), Z => n32);
   U56 : BUF_X1 port map( A => A(4), Z => n34);
   U57 : BUF_X1 port map( A => A(7), Z => n40);
   U58 : BUF_X1 port map( A => A(8), Z => n42);
   U59 : BUF_X1 port map( A => A(11), Z => n48);
   U60 : BUF_X1 port map( A => A(12), Z => n50);
   U61 : BUF_X1 port map( A => A(15), Z => n56);
   U62 : BUF_X1 port map( A => A(0), Z => n26);
   U63 : BUF_X1 port map( A => A(2), Z => n30);
   U64 : BUF_X1 port map( A => A(5), Z => n36);
   U65 : BUF_X1 port map( A => A(6), Z => n38);
   U66 : BUF_X1 port map( A => A(9), Z => n44);
   U67 : BUF_X1 port map( A => A(10), Z => n46);
   U68 : BUF_X1 port map( A => A(13), Z => n52);
   U69 : BUF_X1 port map( A => A(14), Z => n54);
   U70 : BUF_X1 port map( A => n167, Z => n1);
   U71 : BUF_X1 port map( A => n167, Z => n2);
   U72 : BUF_X1 port map( A => n167, Z => n3);
   U73 : AND2_X1 port map( A1 => S(0), A2 => n3, ZN => n69);
   U74 : OAI22_X1 port map( A1 => n84, A2 => n141, B1 => n85, B2 => n59, ZN => 
                           Y(30));
   U75 : AOI21_X1 port map( B1 => n15, B2 => n141, A => n7, ZN => n85);
   U76 : AOI221_X1 port map( B1 => A(30), B2 => n1, C1 => n14, C2 => n59, A => 
                           n6, ZN => n84);
   U77 : INV_X1 port map( A => B(30), ZN => n141);
   U78 : OAI22_X1 port map( A1 => n116, A2 => n155, B1 => n117, B2 => n139, ZN 
                           => Y(16));
   U79 : AOI21_X1 port map( B1 => n17, B2 => n155, A => n8, ZN => n117);
   U80 : AOI221_X1 port map( B1 => A(16), B2 => n3, C1 => n13, C2 => n139, A =>
                           n4, ZN => n116);
   U81 : INV_X1 port map( A => B(16), ZN => n155);
   U82 : OAI22_X1 port map( A1 => n106, A2 => n151, B1 => n107, B2 => n135, ZN 
                           => Y(20));
   U83 : AOI21_X1 port map( B1 => n16, B2 => n151, A => n8, ZN => n107);
   U84 : AOI221_X1 port map( B1 => A(20), B2 => n2, C1 => n13, C2 => n135, A =>
                           n5, ZN => n106);
   U85 : INV_X1 port map( A => B(20), ZN => n151);
   U86 : OAI22_X1 port map( A1 => n98, A2 => n147, B1 => n99, B2 => n65, ZN => 
                           Y(24));
   U87 : AOI21_X1 port map( B1 => n16, B2 => n147, A => n7, ZN => n99);
   U88 : AOI221_X1 port map( B1 => A(24), B2 => n2, C1 => n14, C2 => n65, A => 
                           n6, ZN => n98);
   U89 : INV_X1 port map( A => B(24), ZN => n147);
   U90 : OAI22_X1 port map( A1 => n90, A2 => n143, B1 => n91, B2 => n61, ZN => 
                           Y(28));
   U91 : AOI21_X1 port map( B1 => n15, B2 => n143, A => n7, ZN => n91);
   U92 : AOI221_X1 port map( B1 => A(28), B2 => n1, C1 => n14, C2 => n61, A => 
                           n6, ZN => n90);
   U93 : INV_X1 port map( A => B(28), ZN => n143);
   U94 : OAI22_X1 port map( A1 => n112, A2 => n153, B1 => n113, B2 => n137, ZN 
                           => Y(18));
   U95 : AOI21_X1 port map( B1 => n16, B2 => n153, A => n8, ZN => n113);
   U96 : AOI221_X1 port map( B1 => A(18), B2 => n2, C1 => n13, C2 => n137, A =>
                           n5, ZN => n112);
   U97 : INV_X1 port map( A => B(18), ZN => n153);
   U98 : OAI22_X1 port map( A1 => n102, A2 => n149, B1 => n103, B2 => n133, ZN 
                           => Y(22));
   U99 : AOI21_X1 port map( B1 => n16, B2 => n149, A => n8, ZN => n103);
   U100 : AOI221_X1 port map( B1 => A(22), B2 => n2, C1 => n14, C2 => n133, A 
                           => n5, ZN => n102);
   U101 : INV_X1 port map( A => B(22), ZN => n149);
   U102 : OAI22_X1 port map( A1 => n94, A2 => n145, B1 => n95, B2 => n63, ZN =>
                           Y(26));
   U103 : AOI21_X1 port map( B1 => n16, B2 => n145, A => n7, ZN => n95);
   U104 : AOI221_X1 port map( B1 => A(26), B2 => n2, C1 => n14, C2 => n63, A =>
                           n5, ZN => n94);
   U105 : INV_X1 port map( A => B(26), ZN => n145);
   U106 : OAI22_X1 port map( A1 => n114, A2 => n154, B1 => n115, B2 => n138, ZN
                           => Y(17));
   U107 : AOI21_X1 port map( B1 => n16, B2 => n154, A => n8, ZN => n115);
   U108 : AOI221_X1 port map( B1 => A(17), B2 => n3, C1 => n13, C2 => n138, A 
                           => n5, ZN => n114);
   U109 : INV_X1 port map( A => B(17), ZN => n154);
   U110 : OAI22_X1 port map( A1 => n104, A2 => n150, B1 => n105, B2 => n134, ZN
                           => Y(21));
   U111 : AOI21_X1 port map( B1 => n16, B2 => n150, A => n8, ZN => n105);
   U112 : AOI221_X1 port map( B1 => A(21), B2 => n2, C1 => n13, C2 => n134, A 
                           => n5, ZN => n104);
   U113 : INV_X1 port map( A => B(21), ZN => n150);
   U114 : OAI22_X1 port map( A1 => n96, A2 => n146, B1 => n97, B2 => n64, ZN =>
                           Y(25));
   U115 : AOI21_X1 port map( B1 => n16, B2 => n146, A => n7, ZN => n97);
   U116 : AOI221_X1 port map( B1 => A(25), B2 => n2, C1 => n14, C2 => n64, A =>
                           n6, ZN => n96);
   U117 : INV_X1 port map( A => B(25), ZN => n146);
   U118 : OAI22_X1 port map( A1 => n88, A2 => n142, B1 => n89, B2 => n60, ZN =>
                           Y(29));
   U119 : AOI21_X1 port map( B1 => n15, B2 => n142, A => n7, ZN => n89);
   U120 : AOI221_X1 port map( B1 => A(29), B2 => n1, C1 => n14, C2 => n60, A =>
                           n6, ZN => n88);
   U121 : INV_X1 port map( A => B(29), ZN => n142);
   U122 : OAI22_X1 port map( A1 => n110, A2 => n152, B1 => n111, B2 => n136, ZN
                           => Y(19));
   U123 : AOI21_X1 port map( B1 => n16, B2 => n152, A => n8, ZN => n111);
   U124 : AOI221_X1 port map( B1 => A(19), B2 => n2, C1 => n13, C2 => n136, A 
                           => n5, ZN => n110);
   U125 : INV_X1 port map( A => B(19), ZN => n152);
   U126 : OAI22_X1 port map( A1 => n100, A2 => n148, B1 => n101, B2 => n132, ZN
                           => Y(23));
   U127 : AOI21_X1 port map( B1 => n16, B2 => n148, A => n8, ZN => n101);
   U128 : AOI221_X1 port map( B1 => A(23), B2 => n2, C1 => n13, C2 => n132, A 
                           => n5, ZN => n100);
   U129 : INV_X1 port map( A => B(23), ZN => n148);
   U130 : OAI22_X1 port map( A1 => n92, A2 => n144, B1 => n93, B2 => n62, ZN =>
                           Y(27));
   U131 : AOI21_X1 port map( B1 => n16, B2 => n144, A => n7, ZN => n93);
   U132 : AOI221_X1 port map( B1 => A(27), B2 => n2, C1 => n14, C2 => n62, A =>
                           n6, ZN => n92);
   U133 : INV_X1 port map( A => B(27), ZN => n144);
   U134 : OAI22_X1 port map( A1 => n82, A2 => n140, B1 => n83, B2 => n58, ZN =>
                           Y(31));
   U135 : AOI21_X1 port map( B1 => n15, B2 => n140, A => n7, ZN => n83);
   U136 : AOI221_X1 port map( B1 => A(31), B2 => n1, C1 => n14, C2 => n58, A =>
                           n6, ZN => n82);
   U137 : INV_X1 port map( A => B(31), ZN => n140);
   U138 : INV_X1 port map( A => A(30), ZN => n59);
   U139 : OAI22_X1 port map( A1 => n76, A2 => n166, B1 => n77, B2 => n37, ZN =>
                           Y(5));
   U140 : AOI21_X1 port map( B1 => n15, B2 => n166, A => n6, ZN => n77);
   U141 : INV_X1 port map( A => B(5), ZN => n166);
   U142 : AOI221_X1 port map( B1 => n36, B2 => n1, C1 => n13, C2 => n37, A => 
                           n5, ZN => n76);
   U143 : OAI22_X1 port map( A1 => n74, A2 => n165, B1 => n75, B2 => n39, ZN =>
                           Y(6));
   U144 : AOI21_X1 port map( B1 => n15, B2 => n165, A => n6, ZN => n75);
   U145 : AOI221_X1 port map( B1 => n38, B2 => n1, C1 => n12, C2 => n39, A => 
                           n4, ZN => n74);
   U146 : INV_X1 port map( A => B(6), ZN => n165);
   U147 : OAI22_X1 port map( A1 => n72, A2 => n164, B1 => n73, B2 => n41, ZN =>
                           Y(7));
   U148 : AOI21_X1 port map( B1 => n15, B2 => n164, A => n7, ZN => n73);
   U149 : INV_X1 port map( A => B(7), ZN => n164);
   U150 : AOI221_X1 port map( B1 => n40, B2 => n1, C1 => n12, C2 => n41, A => 
                           n4, ZN => n72);
   U151 : OAI22_X1 port map( A1 => n70, A2 => n163, B1 => n71, B2 => n43, ZN =>
                           Y(8));
   U152 : AOI21_X1 port map( B1 => n15, B2 => n163, A => n6, ZN => n71);
   U153 : INV_X1 port map( A => B(8), ZN => n163);
   U154 : AOI221_X1 port map( B1 => n42, B2 => n1, C1 => n12, C2 => n43, A => 
                           n4, ZN => n70);
   U155 : OAI22_X1 port map( A1 => n66, A2 => n162, B1 => n67, B2 => n45, ZN =>
                           Y(9));
   U156 : AOI21_X1 port map( B1 => n15, B2 => n162, A => n7, ZN => n67);
   U157 : INV_X1 port map( A => B(9), ZN => n162);
   U158 : AOI221_X1 port map( B1 => n44, B2 => n2, C1 => n12, C2 => n45, A => 
                           n4, ZN => n66);
   U159 : OAI22_X1 port map( A1 => n128, A2 => n161, B1 => n129, B2 => n47, ZN 
                           => Y(10));
   U160 : AOI21_X1 port map( B1 => n17, B2 => n161, A => n9, ZN => n129);
   U161 : AOI221_X1 port map( B1 => n46, B2 => n3, C1 => n12, C2 => n47, A => 
                           n4, ZN => n128);
   U162 : INV_X1 port map( A => B(10), ZN => n161);
   U163 : OAI22_X1 port map( A1 => n126, A2 => n160, B1 => n127, B2 => n49, ZN 
                           => Y(11));
   U164 : AOI21_X1 port map( B1 => n17, B2 => n160, A => n9, ZN => n127);
   U165 : INV_X1 port map( A => B(11), ZN => n160);
   U166 : AOI221_X1 port map( B1 => n48, B2 => n3, C1 => n12, C2 => n49, A => 
                           n4, ZN => n126);
   U167 : OAI22_X1 port map( A1 => n124, A2 => n159, B1 => n125, B2 => n51, ZN 
                           => Y(12));
   U168 : AOI21_X1 port map( B1 => n17, B2 => n159, A => n8, ZN => n125);
   U169 : INV_X1 port map( A => B(12), ZN => n159);
   U170 : AOI221_X1 port map( B1 => n50, B2 => n3, C1 => n12, C2 => n51, A => 
                           n4, ZN => n124);
   U171 : OAI22_X1 port map( A1 => n122, A2 => n158, B1 => n123, B2 => n53, ZN 
                           => Y(13));
   U172 : AOI21_X1 port map( B1 => n17, B2 => n158, A => n8, ZN => n123);
   U173 : INV_X1 port map( A => B(13), ZN => n158);
   U174 : AOI221_X1 port map( B1 => n52, B2 => n3, C1 => n12, C2 => n53, A => 
                           n4, ZN => n122);
   U175 : OAI22_X1 port map( A1 => n120, A2 => n157, B1 => n121, B2 => n55, ZN 
                           => Y(14));
   U176 : AOI21_X1 port map( B1 => n17, B2 => n157, A => n8, ZN => n121);
   U177 : AOI221_X1 port map( B1 => n54, B2 => n3, C1 => n12, C2 => n55, A => 
                           n4, ZN => n120);
   U178 : INV_X1 port map( A => B(14), ZN => n157);
   U179 : OAI22_X1 port map( A1 => n118, A2 => n156, B1 => n119, B2 => n57, ZN 
                           => Y(15));
   U180 : AOI21_X1 port map( B1 => n17, B2 => n156, A => n8, ZN => n119);
   U181 : AOI221_X1 port map( B1 => n56, B2 => n3, C1 => n12, C2 => n57, A => 
                           n4, ZN => n118);
   U182 : INV_X1 port map( A => B(15), ZN => n156);
   U183 : INV_X1 port map( A => A(16), ZN => n139);
   U184 : INV_X1 port map( A => A(20), ZN => n135);
   U185 : INV_X1 port map( A => A(24), ZN => n65);
   U186 : INV_X1 port map( A => A(28), ZN => n61);
   U187 : INV_X1 port map( A => A(18), ZN => n137);
   U188 : INV_X1 port map( A => A(22), ZN => n133);
   U189 : INV_X1 port map( A => A(26), ZN => n63);
   U190 : INV_X1 port map( A => A(17), ZN => n138);
   U191 : INV_X1 port map( A => A(21), ZN => n134);
   U192 : INV_X1 port map( A => A(25), ZN => n64);
   U193 : INV_X1 port map( A => A(29), ZN => n60);
   U194 : INV_X1 port map( A => A(19), ZN => n136);
   U195 : INV_X1 port map( A => A(23), ZN => n132);
   U196 : INV_X1 port map( A => A(27), ZN => n62);
   U197 : INV_X1 port map( A => A(31), ZN => n58);
   U198 : INV_X1 port map( A => S(1), ZN => n167);
   U199 : BUF_X1 port map( A => n68, Z => n20);
   U200 : NOR2_X1 port map( A1 => n1, A2 => S(0), ZN => n68);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BARREL_SHIFTER_RIGHT_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end BARREL_SHIFTER_RIGHT_N32;

architecture SYN_STRUCTURAL of BARREL_SHIFTER_RIGHT_N32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_L_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_32
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_33
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_34
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_35
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_36
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_37
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_38
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_39
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_40
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_41
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_42
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_43
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_44
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_45
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_46
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_47
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_48
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_49
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_50
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_51
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_52
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_53
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_54
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_55
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_56
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_57
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_58
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_59
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_60
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_61
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_62
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_63
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_64
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_65
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_66
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_67
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_68
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_69
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_70
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_71
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_72
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_73
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_74
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_75
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_76
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_77
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_78
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_79
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_80
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_81
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_82
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_83
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_84
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_85
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_86
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_87
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_88
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_89
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_90
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_91
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_92
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_93
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_94
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_95
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_96
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_97
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_98
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_99
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_100
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_101
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_102
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_103
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_104
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_105
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_106
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_107
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_108
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_109
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_110
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_111
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_112
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_113
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_114
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_115
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_116
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_117
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_118
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_119
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_120
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_121
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_122
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_123
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_124
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_125
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_126
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_127
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_128
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_129
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_130
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_131
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_132
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_133
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_134
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_135
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_136
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_137
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_138
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_139
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_140
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_141
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_142
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_143
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_144
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_145
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_146
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_147
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_148
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_149
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_150
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_151
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_152
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_153
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_154
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_155
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_156
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_157
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_158
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_159
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal TMP_4_31_port, TMP_4_30_port, TMP_4_29_port, TMP_4_28_port, 
      TMP_4_27_port, TMP_4_26_port, TMP_4_25_port, TMP_4_24_port, TMP_4_23_port
      , TMP_4_22_port, TMP_4_21_port, TMP_4_20_port, TMP_4_19_port, 
      TMP_4_18_port, TMP_4_17_port, TMP_4_16_port, TMP_4_15_port, TMP_4_14_port
      , TMP_4_13_port, TMP_4_12_port, TMP_4_11_port, TMP_4_10_port, 
      TMP_4_9_port, TMP_4_8_port, TMP_4_7_port, TMP_4_6_port, TMP_4_5_port, 
      TMP_4_4_port, TMP_4_3_port, TMP_4_2_port, TMP_4_1_port, TMP_4_0_port, 
      TMP_3_31_port, TMP_3_30_port, TMP_3_29_port, TMP_3_28_port, TMP_3_27_port
      , TMP_3_26_port, TMP_3_25_port, TMP_3_24_port, TMP_3_23_port, 
      TMP_3_22_port, TMP_3_21_port, TMP_3_20_port, TMP_3_19_port, TMP_3_18_port
      , TMP_3_17_port, TMP_3_16_port, TMP_3_15_port, TMP_3_14_port, 
      TMP_3_13_port, TMP_3_12_port, TMP_3_11_port, TMP_3_10_port, TMP_3_9_port,
      TMP_3_8_port, TMP_3_7_port, TMP_3_6_port, TMP_3_5_port, TMP_3_4_port, 
      TMP_3_3_port, TMP_3_2_port, TMP_3_1_port, TMP_3_0_port, TMP_2_31_port, 
      TMP_2_30_port, TMP_2_29_port, TMP_2_28_port, TMP_2_27_port, TMP_2_26_port
      , TMP_2_25_port, TMP_2_24_port, TMP_2_23_port, TMP_2_22_port, 
      TMP_2_21_port, TMP_2_20_port, TMP_2_19_port, TMP_2_18_port, TMP_2_17_port
      , TMP_2_16_port, TMP_2_15_port, TMP_2_14_port, TMP_2_13_port, 
      TMP_2_12_port, TMP_2_11_port, TMP_2_10_port, TMP_2_9_port, TMP_2_8_port, 
      TMP_2_7_port, TMP_2_6_port, TMP_2_5_port, TMP_2_4_port, TMP_2_3_port, 
      TMP_2_2_port, TMP_2_1_port, TMP_2_0_port, TMP_1_31_port, TMP_1_30_port, 
      TMP_1_29_port, TMP_1_28_port, TMP_1_27_port, TMP_1_26_port, TMP_1_25_port
      , TMP_1_24_port, TMP_1_23_port, TMP_1_22_port, TMP_1_21_port, 
      TMP_1_20_port, TMP_1_19_port, TMP_1_18_port, TMP_1_17_port, TMP_1_16_port
      , TMP_1_15_port, TMP_1_14_port, TMP_1_13_port, TMP_1_12_port, 
      TMP_1_11_port, TMP_1_10_port, TMP_1_9_port, TMP_1_8_port, TMP_1_7_port, 
      TMP_1_6_port, TMP_1_5_port, TMP_1_4_port, TMP_1_3_port, TMP_1_2_port, 
      TMP_1_1_port, TMP_1_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24 : 
      std_logic;

begin
   
   MUX21_K_0_0 : MUX21_L_159 port map( A => A(0), B => A(1), S => n5, Y => 
                           TMP_1_0_port);
   MUX21_K_0_1 : MUX21_L_158 port map( A => A(1), B => A(2), S => n5, Y => 
                           TMP_1_1_port);
   MUX21_K_0_2 : MUX21_L_157 port map( A => A(2), B => A(3), S => n5, Y => 
                           TMP_1_2_port);
   MUX21_K_0_3 : MUX21_L_156 port map( A => A(3), B => A(4), S => n5, Y => 
                           TMP_1_3_port);
   MUX21_K_0_4 : MUX21_L_155 port map( A => A(4), B => A(5), S => n5, Y => 
                           TMP_1_4_port);
   MUX21_K_0_5 : MUX21_L_154 port map( A => A(5), B => A(6), S => n5, Y => 
                           TMP_1_5_port);
   MUX21_K_0_6 : MUX21_L_153 port map( A => A(6), B => A(7), S => n5, Y => 
                           TMP_1_6_port);
   MUX21_K_0_7 : MUX21_L_152 port map( A => A(7), B => A(8), S => n5, Y => 
                           TMP_1_7_port);
   MUX21_K_0_8 : MUX21_L_151 port map( A => A(8), B => A(9), S => n5, Y => 
                           TMP_1_8_port);
   MUX21_K_0_9 : MUX21_L_150 port map( A => A(9), B => A(10), S => n5, Y => 
                           TMP_1_9_port);
   MUX21_K_0_10 : MUX21_L_149 port map( A => A(10), B => A(11), S => n5, Y => 
                           TMP_1_10_port);
   MUX21_K_0_11 : MUX21_L_148 port map( A => A(11), B => A(12), S => n5, Y => 
                           TMP_1_11_port);
   MUX21_K_0_12 : MUX21_L_147 port map( A => A(12), B => A(13), S => n6, Y => 
                           TMP_1_12_port);
   MUX21_K_0_13 : MUX21_L_146 port map( A => A(13), B => A(14), S => n6, Y => 
                           TMP_1_13_port);
   MUX21_K_0_14 : MUX21_L_145 port map( A => A(14), B => A(15), S => n6, Y => 
                           TMP_1_14_port);
   MUX21_K_0_15 : MUX21_L_144 port map( A => A(15), B => A(16), S => n6, Y => 
                           TMP_1_15_port);
   MUX21_K_0_16 : MUX21_L_143 port map( A => A(16), B => A(17), S => n6, Y => 
                           TMP_1_16_port);
   MUX21_K_0_17 : MUX21_L_142 port map( A => A(17), B => A(18), S => n6, Y => 
                           TMP_1_17_port);
   MUX21_K_0_18 : MUX21_L_141 port map( A => A(18), B => A(19), S => n6, Y => 
                           TMP_1_18_port);
   MUX21_K_0_19 : MUX21_L_140 port map( A => A(19), B => A(20), S => n6, Y => 
                           TMP_1_19_port);
   MUX21_K_0_20 : MUX21_L_139 port map( A => A(20), B => A(21), S => n6, Y => 
                           TMP_1_20_port);
   MUX21_K_0_21 : MUX21_L_138 port map( A => A(21), B => A(22), S => n6, Y => 
                           TMP_1_21_port);
   MUX21_K_0_22 : MUX21_L_137 port map( A => A(22), B => A(23), S => n6, Y => 
                           TMP_1_22_port);
   MUX21_K_0_23 : MUX21_L_136 port map( A => A(23), B => A(24), S => n6, Y => 
                           TMP_1_23_port);
   MUX21_K_0_24 : MUX21_L_135 port map( A => A(24), B => A(25), S => n7, Y => 
                           TMP_1_24_port);
   MUX21_K_0_25 : MUX21_L_134 port map( A => A(25), B => A(26), S => n7, Y => 
                           TMP_1_25_port);
   MUX21_K_0_26 : MUX21_L_133 port map( A => A(26), B => A(27), S => n7, Y => 
                           TMP_1_26_port);
   MUX21_K_0_27 : MUX21_L_132 port map( A => A(27), B => A(28), S => n7, Y => 
                           TMP_1_27_port);
   MUX21_K_0_28 : MUX21_L_131 port map( A => A(28), B => A(29), S => n7, Y => 
                           TMP_1_28_port);
   MUX21_K_0_29 : MUX21_L_130 port map( A => A(29), B => A(30), S => n7, Y => 
                           TMP_1_29_port);
   MUX21_K_0_30 : MUX21_L_129 port map( A => A(30), B => A(31), S => n7, Y => 
                           TMP_1_30_port);
   MUX21_J_0_0 : MUX21_L_128 port map( A => A(31), B => n1, S => n7, Y => 
                           TMP_1_31_port);
   MUX21_K_1_0 : MUX21_L_127 port map( A => TMP_1_0_port, B => TMP_1_2_port, S 
                           => n9, Y => TMP_2_0_port);
   MUX21_K_1_1 : MUX21_L_126 port map( A => TMP_1_1_port, B => TMP_1_3_port, S 
                           => n9, Y => TMP_2_1_port);
   MUX21_K_1_2 : MUX21_L_125 port map( A => TMP_1_2_port, B => TMP_1_4_port, S 
                           => n9, Y => TMP_2_2_port);
   MUX21_K_1_3 : MUX21_L_124 port map( A => TMP_1_3_port, B => TMP_1_5_port, S 
                           => n9, Y => TMP_2_3_port);
   MUX21_K_1_4 : MUX21_L_123 port map( A => TMP_1_4_port, B => TMP_1_6_port, S 
                           => n9, Y => TMP_2_4_port);
   MUX21_K_1_5 : MUX21_L_122 port map( A => TMP_1_5_port, B => TMP_1_7_port, S 
                           => n9, Y => TMP_2_5_port);
   MUX21_K_1_6 : MUX21_L_121 port map( A => TMP_1_6_port, B => TMP_1_8_port, S 
                           => n9, Y => TMP_2_6_port);
   MUX21_K_1_7 : MUX21_L_120 port map( A => TMP_1_7_port, B => TMP_1_9_port, S 
                           => n9, Y => TMP_2_7_port);
   MUX21_K_1_8 : MUX21_L_119 port map( A => TMP_1_8_port, B => TMP_1_10_port, S
                           => n9, Y => TMP_2_8_port);
   MUX21_K_1_9 : MUX21_L_118 port map( A => TMP_1_9_port, B => TMP_1_11_port, S
                           => n9, Y => TMP_2_9_port);
   MUX21_K_1_10 : MUX21_L_117 port map( A => TMP_1_10_port, B => TMP_1_12_port,
                           S => n9, Y => TMP_2_10_port);
   MUX21_K_1_11 : MUX21_L_116 port map( A => TMP_1_11_port, B => TMP_1_13_port,
                           S => n9, Y => TMP_2_11_port);
   MUX21_K_1_12 : MUX21_L_115 port map( A => TMP_1_12_port, B => TMP_1_14_port,
                           S => n10, Y => TMP_2_12_port);
   MUX21_K_1_13 : MUX21_L_114 port map( A => TMP_1_13_port, B => TMP_1_15_port,
                           S => n10, Y => TMP_2_13_port);
   MUX21_K_1_14 : MUX21_L_113 port map( A => TMP_1_14_port, B => TMP_1_16_port,
                           S => n10, Y => TMP_2_14_port);
   MUX21_K_1_15 : MUX21_L_112 port map( A => TMP_1_15_port, B => TMP_1_17_port,
                           S => n10, Y => TMP_2_15_port);
   MUX21_K_1_16 : MUX21_L_111 port map( A => TMP_1_16_port, B => TMP_1_18_port,
                           S => n10, Y => TMP_2_16_port);
   MUX21_K_1_17 : MUX21_L_110 port map( A => TMP_1_17_port, B => TMP_1_19_port,
                           S => n10, Y => TMP_2_17_port);
   MUX21_K_1_18 : MUX21_L_109 port map( A => TMP_1_18_port, B => TMP_1_20_port,
                           S => n10, Y => TMP_2_18_port);
   MUX21_K_1_19 : MUX21_L_108 port map( A => TMP_1_19_port, B => TMP_1_21_port,
                           S => n10, Y => TMP_2_19_port);
   MUX21_K_1_20 : MUX21_L_107 port map( A => TMP_1_20_port, B => TMP_1_22_port,
                           S => n10, Y => TMP_2_20_port);
   MUX21_K_1_21 : MUX21_L_106 port map( A => TMP_1_21_port, B => TMP_1_23_port,
                           S => n10, Y => TMP_2_21_port);
   MUX21_K_1_22 : MUX21_L_105 port map( A => TMP_1_22_port, B => TMP_1_24_port,
                           S => n10, Y => TMP_2_22_port);
   MUX21_K_1_23 : MUX21_L_104 port map( A => TMP_1_23_port, B => TMP_1_25_port,
                           S => n10, Y => TMP_2_23_port);
   MUX21_K_1_24 : MUX21_L_103 port map( A => TMP_1_24_port, B => TMP_1_26_port,
                           S => n11, Y => TMP_2_24_port);
   MUX21_K_1_25 : MUX21_L_102 port map( A => TMP_1_25_port, B => TMP_1_27_port,
                           S => n11, Y => TMP_2_25_port);
   MUX21_K_1_26 : MUX21_L_101 port map( A => TMP_1_26_port, B => TMP_1_28_port,
                           S => n11, Y => TMP_2_26_port);
   MUX21_K_1_27 : MUX21_L_100 port map( A => TMP_1_27_port, B => TMP_1_29_port,
                           S => n11, Y => TMP_2_27_port);
   MUX21_K_1_28 : MUX21_L_99 port map( A => TMP_1_28_port, B => TMP_1_30_port, 
                           S => n11, Y => TMP_2_28_port);
   MUX21_K_1_29 : MUX21_L_98 port map( A => TMP_1_29_port, B => TMP_1_31_port, 
                           S => n11, Y => TMP_2_29_port);
   MUX21_J_1_0 : MUX21_L_97 port map( A => TMP_1_30_port, B => n1, S => n11, Y 
                           => TMP_2_30_port);
   MUX21_J_1_1 : MUX21_L_96 port map( A => TMP_1_31_port, B => n1, S => n11, Y 
                           => TMP_2_31_port);
   MUX21_K_2_0 : MUX21_L_95 port map( A => TMP_2_0_port, B => TMP_2_4_port, S 
                           => n13, Y => TMP_3_0_port);
   MUX21_K_2_1 : MUX21_L_94 port map( A => TMP_2_1_port, B => TMP_2_5_port, S 
                           => n13, Y => TMP_3_1_port);
   MUX21_K_2_2 : MUX21_L_93 port map( A => TMP_2_2_port, B => TMP_2_6_port, S 
                           => n13, Y => TMP_3_2_port);
   MUX21_K_2_3 : MUX21_L_92 port map( A => TMP_2_3_port, B => TMP_2_7_port, S 
                           => n13, Y => TMP_3_3_port);
   MUX21_K_2_4 : MUX21_L_91 port map( A => TMP_2_4_port, B => TMP_2_8_port, S 
                           => n13, Y => TMP_3_4_port);
   MUX21_K_2_5 : MUX21_L_90 port map( A => TMP_2_5_port, B => TMP_2_9_port, S 
                           => n13, Y => TMP_3_5_port);
   MUX21_K_2_6 : MUX21_L_89 port map( A => TMP_2_6_port, B => TMP_2_10_port, S 
                           => n13, Y => TMP_3_6_port);
   MUX21_K_2_7 : MUX21_L_88 port map( A => TMP_2_7_port, B => TMP_2_11_port, S 
                           => n13, Y => TMP_3_7_port);
   MUX21_K_2_8 : MUX21_L_87 port map( A => TMP_2_8_port, B => TMP_2_12_port, S 
                           => n13, Y => TMP_3_8_port);
   MUX21_K_2_9 : MUX21_L_86 port map( A => TMP_2_9_port, B => TMP_2_13_port, S 
                           => n13, Y => TMP_3_9_port);
   MUX21_K_2_10 : MUX21_L_85 port map( A => TMP_2_10_port, B => TMP_2_14_port, 
                           S => n13, Y => TMP_3_10_port);
   MUX21_K_2_11 : MUX21_L_84 port map( A => TMP_2_11_port, B => TMP_2_15_port, 
                           S => n13, Y => TMP_3_11_port);
   MUX21_K_2_12 : MUX21_L_83 port map( A => TMP_2_12_port, B => TMP_2_16_port, 
                           S => n14, Y => TMP_3_12_port);
   MUX21_K_2_13 : MUX21_L_82 port map( A => TMP_2_13_port, B => TMP_2_17_port, 
                           S => n14, Y => TMP_3_13_port);
   MUX21_K_2_14 : MUX21_L_81 port map( A => TMP_2_14_port, B => TMP_2_18_port, 
                           S => n14, Y => TMP_3_14_port);
   MUX21_K_2_15 : MUX21_L_80 port map( A => TMP_2_15_port, B => TMP_2_19_port, 
                           S => n14, Y => TMP_3_15_port);
   MUX21_K_2_16 : MUX21_L_79 port map( A => TMP_2_16_port, B => TMP_2_20_port, 
                           S => n14, Y => TMP_3_16_port);
   MUX21_K_2_17 : MUX21_L_78 port map( A => TMP_2_17_port, B => TMP_2_21_port, 
                           S => n14, Y => TMP_3_17_port);
   MUX21_K_2_18 : MUX21_L_77 port map( A => TMP_2_18_port, B => TMP_2_22_port, 
                           S => n14, Y => TMP_3_18_port);
   MUX21_K_2_19 : MUX21_L_76 port map( A => TMP_2_19_port, B => TMP_2_23_port, 
                           S => n14, Y => TMP_3_19_port);
   MUX21_K_2_20 : MUX21_L_75 port map( A => TMP_2_20_port, B => TMP_2_24_port, 
                           S => n14, Y => TMP_3_20_port);
   MUX21_K_2_21 : MUX21_L_74 port map( A => TMP_2_21_port, B => TMP_2_25_port, 
                           S => n14, Y => TMP_3_21_port);
   MUX21_K_2_22 : MUX21_L_73 port map( A => TMP_2_22_port, B => TMP_2_26_port, 
                           S => n14, Y => TMP_3_22_port);
   MUX21_K_2_23 : MUX21_L_72 port map( A => TMP_2_23_port, B => TMP_2_27_port, 
                           S => n14, Y => TMP_3_23_port);
   MUX21_K_2_24 : MUX21_L_71 port map( A => TMP_2_24_port, B => TMP_2_28_port, 
                           S => n15, Y => TMP_3_24_port);
   MUX21_K_2_25 : MUX21_L_70 port map( A => TMP_2_25_port, B => TMP_2_29_port, 
                           S => n15, Y => TMP_3_25_port);
   MUX21_K_2_26 : MUX21_L_69 port map( A => TMP_2_26_port, B => TMP_2_30_port, 
                           S => n15, Y => TMP_3_26_port);
   MUX21_K_2_27 : MUX21_L_68 port map( A => TMP_2_27_port, B => TMP_2_31_port, 
                           S => n15, Y => TMP_3_27_port);
   MUX21_J_2_0 : MUX21_L_67 port map( A => TMP_2_28_port, B => n1, S => n15, Y 
                           => TMP_3_28_port);
   MUX21_J_2_1 : MUX21_L_66 port map( A => TMP_2_29_port, B => n1, S => n15, Y 
                           => TMP_3_29_port);
   MUX21_J_2_2 : MUX21_L_65 port map( A => TMP_2_30_port, B => n1, S => n15, Y 
                           => TMP_3_30_port);
   MUX21_J_2_3 : MUX21_L_64 port map( A => TMP_2_31_port, B => n1, S => n15, Y 
                           => TMP_3_31_port);
   MUX21_K_3_0 : MUX21_L_63 port map( A => TMP_3_0_port, B => TMP_3_8_port, S 
                           => n17, Y => TMP_4_0_port);
   MUX21_K_3_1 : MUX21_L_62 port map( A => TMP_3_1_port, B => TMP_3_9_port, S 
                           => n17, Y => TMP_4_1_port);
   MUX21_K_3_2 : MUX21_L_61 port map( A => TMP_3_2_port, B => TMP_3_10_port, S 
                           => n17, Y => TMP_4_2_port);
   MUX21_K_3_3 : MUX21_L_60 port map( A => TMP_3_3_port, B => TMP_3_11_port, S 
                           => n17, Y => TMP_4_3_port);
   MUX21_K_3_4 : MUX21_L_59 port map( A => TMP_3_4_port, B => TMP_3_12_port, S 
                           => n17, Y => TMP_4_4_port);
   MUX21_K_3_5 : MUX21_L_58 port map( A => TMP_3_5_port, B => TMP_3_13_port, S 
                           => n17, Y => TMP_4_5_port);
   MUX21_K_3_6 : MUX21_L_57 port map( A => TMP_3_6_port, B => TMP_3_14_port, S 
                           => n17, Y => TMP_4_6_port);
   MUX21_K_3_7 : MUX21_L_56 port map( A => TMP_3_7_port, B => TMP_3_15_port, S 
                           => n17, Y => TMP_4_7_port);
   MUX21_K_3_8 : MUX21_L_55 port map( A => TMP_3_8_port, B => TMP_3_16_port, S 
                           => n17, Y => TMP_4_8_port);
   MUX21_K_3_9 : MUX21_L_54 port map( A => TMP_3_9_port, B => TMP_3_17_port, S 
                           => n17, Y => TMP_4_9_port);
   MUX21_K_3_10 : MUX21_L_53 port map( A => TMP_3_10_port, B => TMP_3_18_port, 
                           S => n17, Y => TMP_4_10_port);
   MUX21_K_3_11 : MUX21_L_52 port map( A => TMP_3_11_port, B => TMP_3_19_port, 
                           S => n17, Y => TMP_4_11_port);
   MUX21_K_3_12 : MUX21_L_51 port map( A => TMP_3_12_port, B => TMP_3_20_port, 
                           S => n18, Y => TMP_4_12_port);
   MUX21_K_3_13 : MUX21_L_50 port map( A => TMP_3_13_port, B => TMP_3_21_port, 
                           S => n18, Y => TMP_4_13_port);
   MUX21_K_3_14 : MUX21_L_49 port map( A => TMP_3_14_port, B => TMP_3_22_port, 
                           S => n18, Y => TMP_4_14_port);
   MUX21_K_3_15 : MUX21_L_48 port map( A => TMP_3_15_port, B => TMP_3_23_port, 
                           S => n18, Y => TMP_4_15_port);
   MUX21_K_3_16 : MUX21_L_47 port map( A => TMP_3_16_port, B => TMP_3_24_port, 
                           S => n18, Y => TMP_4_16_port);
   MUX21_K_3_17 : MUX21_L_46 port map( A => TMP_3_17_port, B => TMP_3_25_port, 
                           S => n18, Y => TMP_4_17_port);
   MUX21_K_3_18 : MUX21_L_45 port map( A => TMP_3_18_port, B => TMP_3_26_port, 
                           S => n18, Y => TMP_4_18_port);
   MUX21_K_3_19 : MUX21_L_44 port map( A => TMP_3_19_port, B => TMP_3_27_port, 
                           S => n18, Y => TMP_4_19_port);
   MUX21_K_3_20 : MUX21_L_43 port map( A => TMP_3_20_port, B => TMP_3_28_port, 
                           S => n18, Y => TMP_4_20_port);
   MUX21_K_3_21 : MUX21_L_42 port map( A => TMP_3_21_port, B => TMP_3_29_port, 
                           S => n18, Y => TMP_4_21_port);
   MUX21_K_3_22 : MUX21_L_41 port map( A => TMP_3_22_port, B => TMP_3_30_port, 
                           S => n18, Y => TMP_4_22_port);
   MUX21_K_3_23 : MUX21_L_40 port map( A => TMP_3_23_port, B => TMP_3_31_port, 
                           S => n18, Y => TMP_4_23_port);
   MUX21_J_3_0 : MUX21_L_39 port map( A => TMP_3_24_port, B => n1, S => n19, Y 
                           => TMP_4_24_port);
   MUX21_J_3_1 : MUX21_L_38 port map( A => TMP_3_25_port, B => n1, S => n19, Y 
                           => TMP_4_25_port);
   MUX21_J_3_2 : MUX21_L_37 port map( A => TMP_3_26_port, B => n1, S => n19, Y 
                           => TMP_4_26_port);
   MUX21_J_3_3 : MUX21_L_36 port map( A => TMP_3_27_port, B => n1, S => n19, Y 
                           => TMP_4_27_port);
   MUX21_J_3_4 : MUX21_L_35 port map( A => TMP_3_28_port, B => n1, S => n19, Y 
                           => TMP_4_28_port);
   MUX21_J_3_5 : MUX21_L_34 port map( A => TMP_3_29_port, B => n2, S => n19, Y 
                           => TMP_4_29_port);
   MUX21_J_3_6 : MUX21_L_33 port map( A => TMP_3_30_port, B => n2, S => n19, Y 
                           => TMP_4_30_port);
   MUX21_J_3_7 : MUX21_L_32 port map( A => TMP_3_31_port, B => n2, S => n19, Y 
                           => TMP_4_31_port);
   MUX21_K_4_0 : MUX21_L_31 port map( A => TMP_4_0_port, B => TMP_4_16_port, S 
                           => n21, Y => Y(0));
   MUX21_K_4_1 : MUX21_L_30 port map( A => TMP_4_1_port, B => TMP_4_17_port, S 
                           => n21, Y => Y(1));
   MUX21_K_4_2 : MUX21_L_29 port map( A => TMP_4_2_port, B => TMP_4_18_port, S 
                           => n21, Y => Y(2));
   MUX21_K_4_3 : MUX21_L_28 port map( A => TMP_4_3_port, B => TMP_4_19_port, S 
                           => n21, Y => Y(3));
   MUX21_K_4_4 : MUX21_L_27 port map( A => TMP_4_4_port, B => TMP_4_20_port, S 
                           => n21, Y => Y(4));
   MUX21_K_4_5 : MUX21_L_26 port map( A => TMP_4_5_port, B => TMP_4_21_port, S 
                           => n21, Y => Y(5));
   MUX21_K_4_6 : MUX21_L_25 port map( A => TMP_4_6_port, B => TMP_4_22_port, S 
                           => n21, Y => Y(6));
   MUX21_K_4_7 : MUX21_L_24 port map( A => TMP_4_7_port, B => TMP_4_23_port, S 
                           => n21, Y => Y(7));
   MUX21_K_4_8 : MUX21_L_23 port map( A => TMP_4_8_port, B => TMP_4_24_port, S 
                           => n21, Y => Y(8));
   MUX21_K_4_9 : MUX21_L_22 port map( A => TMP_4_9_port, B => TMP_4_25_port, S 
                           => n21, Y => Y(9));
   MUX21_K_4_10 : MUX21_L_21 port map( A => TMP_4_10_port, B => TMP_4_26_port, 
                           S => n21, Y => Y(10));
   MUX21_K_4_11 : MUX21_L_20 port map( A => TMP_4_11_port, B => TMP_4_27_port, 
                           S => n21, Y => Y(11));
   MUX21_K_4_12 : MUX21_L_19 port map( A => TMP_4_12_port, B => TMP_4_28_port, 
                           S => n22, Y => Y(12));
   MUX21_K_4_13 : MUX21_L_18 port map( A => TMP_4_13_port, B => TMP_4_29_port, 
                           S => n22, Y => Y(13));
   MUX21_K_4_14 : MUX21_L_17 port map( A => TMP_4_14_port, B => TMP_4_30_port, 
                           S => n22, Y => Y(14));
   MUX21_K_4_15 : MUX21_L_16 port map( A => TMP_4_15_port, B => TMP_4_31_port, 
                           S => n22, Y => Y(15));
   MUX21_J_4_0 : MUX21_L_15 port map( A => TMP_4_16_port, B => n2, S => n22, Y 
                           => Y(16));
   MUX21_J_4_1 : MUX21_L_14 port map( A => TMP_4_17_port, B => n2, S => n22, Y 
                           => Y(17));
   MUX21_J_4_2 : MUX21_L_13 port map( A => TMP_4_18_port, B => n2, S => n22, Y 
                           => Y(18));
   MUX21_J_4_3 : MUX21_L_12 port map( A => TMP_4_19_port, B => n2, S => n22, Y 
                           => Y(19));
   MUX21_J_4_4 : MUX21_L_11 port map( A => TMP_4_20_port, B => n2, S => n22, Y 
                           => Y(20));
   MUX21_J_4_5 : MUX21_L_10 port map( A => TMP_4_21_port, B => n2, S => n22, Y 
                           => Y(21));
   MUX21_J_4_6 : MUX21_L_9 port map( A => TMP_4_22_port, B => n2, S => n22, Y 
                           => Y(22));
   MUX21_J_4_7 : MUX21_L_8 port map( A => TMP_4_23_port, B => n2, S => n22, Y 
                           => Y(23));
   MUX21_J_4_8 : MUX21_L_7 port map( A => TMP_4_24_port, B => n2, S => n23, Y 
                           => Y(24));
   MUX21_J_4_9 : MUX21_L_6 port map( A => TMP_4_25_port, B => n3, S => n23, Y 
                           => Y(25));
   MUX21_J_4_10 : MUX21_L_5 port map( A => TMP_4_26_port, B => n3, S => n23, Y 
                           => Y(26));
   MUX21_J_4_11 : MUX21_L_4 port map( A => TMP_4_27_port, B => n3, S => n23, Y 
                           => Y(27));
   MUX21_J_4_12 : MUX21_L_3 port map( A => TMP_4_28_port, B => n3, S => n23, Y 
                           => Y(28));
   MUX21_J_4_13 : MUX21_L_2 port map( A => TMP_4_29_port, B => n3, S => n23, Y 
                           => Y(29));
   MUX21_J_4_14 : MUX21_L_1 port map( A => TMP_4_30_port, B => n3, S => n23, Y 
                           => Y(30));
   MUX21_J_4_15 : MUX21_L_0 port map( A => TMP_4_31_port, B => n3, S => n23, Y 
                           => Y(31));
   U1 : BUF_X1 port map( A => n24, Z => n22);
   U2 : BUF_X1 port map( A => n20, Z => n17);
   U3 : BUF_X1 port map( A => n20, Z => n18);
   U4 : BUF_X1 port map( A => n16, Z => n13);
   U5 : BUF_X1 port map( A => n24, Z => n21);
   U6 : BUF_X1 port map( A => B(3), Z => n20);
   U7 : BUF_X1 port map( A => B(4), Z => n24);
   U8 : BUF_X1 port map( A => B(2), Z => n16);
   U9 : BUF_X1 port map( A => B(1), Z => n12);
   U10 : BUF_X1 port map( A => B(0), Z => n8);
   U11 : BUF_X1 port map( A => S, Z => n4);
   U12 : BUF_X1 port map( A => n8, Z => n5);
   U13 : BUF_X1 port map( A => n8, Z => n6);
   U14 : BUF_X1 port map( A => n12, Z => n9);
   U15 : BUF_X1 port map( A => n12, Z => n10);
   U16 : BUF_X1 port map( A => n16, Z => n14);
   U17 : BUF_X1 port map( A => n8, Z => n7);
   U18 : BUF_X1 port map( A => n12, Z => n11);
   U19 : BUF_X1 port map( A => n16, Z => n15);
   U20 : BUF_X1 port map( A => n20, Z => n19);
   U21 : BUF_X1 port map( A => n24, Z => n23);
   U22 : BUF_X1 port map( A => n4, Z => n1);
   U23 : BUF_X1 port map( A => n4, Z => n2);
   U24 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BARREL_SHIFTER_LEFT_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
         (31 downto 0));

end BARREL_SHIFTER_LEFT_N32;

architecture SYN_STRUCTURAL of BARREL_SHIFTER_LEFT_N32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_L_160
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_161
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_162
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_163
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_164
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_165
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_166
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_167
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_168
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_169
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_170
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_171
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_172
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_173
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_174
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_175
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_176
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_177
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_178
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_179
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_180
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_181
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_182
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_183
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_184
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_185
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_186
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_187
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_188
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_189
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_190
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_191
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_192
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_193
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_194
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_195
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_196
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_197
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_198
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_199
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_200
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_201
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_202
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_203
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_204
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_205
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_206
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_207
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_208
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_209
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_210
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_211
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_212
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_213
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_214
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_215
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_216
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_217
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_218
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_219
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_220
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_221
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_222
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_223
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_224
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_225
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_226
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_227
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_228
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_229
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_230
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_231
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_232
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_233
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_234
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_235
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_236
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_237
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_238
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_239
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_240
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_241
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_242
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_243
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_244
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_245
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_246
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_247
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_248
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_249
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_250
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_251
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_252
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_253
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_254
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_255
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_256
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_257
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_258
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_259
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_260
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_261
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_262
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_263
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_264
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_265
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_266
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_267
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_268
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_269
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_270
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_271
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_272
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_273
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_274
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_275
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_276
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_277
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_278
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_279
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_280
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_281
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_282
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_283
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_284
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_285
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_286
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_287
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_288
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_289
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_290
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_291
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_292
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_293
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_294
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_295
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_296
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_297
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_298
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_299
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_300
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_301
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_302
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_303
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_304
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_305
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_306
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_307
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_308
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_309
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_310
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_311
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_312
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_313
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_314
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_315
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_316
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_317
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_318
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_319
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, TMP_4_31_port, TMP_4_30_port, TMP_4_29_port, 
      TMP_4_28_port, TMP_4_27_port, TMP_4_26_port, TMP_4_25_port, TMP_4_24_port
      , TMP_4_23_port, TMP_4_22_port, TMP_4_21_port, TMP_4_20_port, 
      TMP_4_19_port, TMP_4_18_port, TMP_4_17_port, TMP_4_16_port, TMP_4_15_port
      , TMP_4_14_port, TMP_4_13_port, TMP_4_12_port, TMP_4_11_port, 
      TMP_4_10_port, TMP_4_9_port, TMP_4_8_port, TMP_4_7_port, TMP_4_6_port, 
      TMP_4_5_port, TMP_4_4_port, TMP_4_3_port, TMP_4_2_port, TMP_4_1_port, 
      TMP_4_0_port, TMP_3_31_port, TMP_3_30_port, TMP_3_29_port, TMP_3_28_port,
      TMP_3_27_port, TMP_3_26_port, TMP_3_25_port, TMP_3_24_port, TMP_3_23_port
      , TMP_3_22_port, TMP_3_21_port, TMP_3_20_port, TMP_3_19_port, 
      TMP_3_18_port, TMP_3_17_port, TMP_3_16_port, TMP_3_15_port, TMP_3_14_port
      , TMP_3_13_port, TMP_3_12_port, TMP_3_11_port, TMP_3_10_port, 
      TMP_3_9_port, TMP_3_8_port, TMP_3_7_port, TMP_3_6_port, TMP_3_5_port, 
      TMP_3_4_port, TMP_3_3_port, TMP_3_2_port, TMP_3_1_port, TMP_3_0_port, 
      TMP_2_31_port, TMP_2_30_port, TMP_2_29_port, TMP_2_28_port, TMP_2_27_port
      , TMP_2_26_port, TMP_2_25_port, TMP_2_24_port, TMP_2_23_port, 
      TMP_2_22_port, TMP_2_21_port, TMP_2_20_port, TMP_2_19_port, TMP_2_18_port
      , TMP_2_17_port, TMP_2_16_port, TMP_2_15_port, TMP_2_14_port, 
      TMP_2_13_port, TMP_2_12_port, TMP_2_11_port, TMP_2_10_port, TMP_2_9_port,
      TMP_2_8_port, TMP_2_7_port, TMP_2_6_port, TMP_2_5_port, TMP_2_4_port, 
      TMP_2_3_port, TMP_2_2_port, TMP_2_1_port, TMP_2_0_port, TMP_1_31_port, 
      TMP_1_30_port, TMP_1_29_port, TMP_1_28_port, TMP_1_27_port, TMP_1_26_port
      , TMP_1_25_port, TMP_1_24_port, TMP_1_23_port, TMP_1_22_port, 
      TMP_1_21_port, TMP_1_20_port, TMP_1_19_port, TMP_1_18_port, TMP_1_17_port
      , TMP_1_16_port, TMP_1_15_port, TMP_1_14_port, TMP_1_13_port, 
      TMP_1_12_port, TMP_1_11_port, TMP_1_10_port, TMP_1_9_port, TMP_1_8_port, 
      TMP_1_7_port, TMP_1_6_port, TMP_1_5_port, TMP_1_4_port, TMP_1_3_port, 
      TMP_1_2_port, TMP_1_1_port, TMP_1_0_port, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20 : std_logic;

begin
   
   X_Logic0_port <= '0';
   MUX21_J_0_0 : MUX21_L_319 port map( A => A(0), B => X_Logic0_port, S => n1, 
                           Y => TMP_1_0_port);
   MUX21_K_0_0 : MUX21_L_318 port map( A => A(1), B => A(0), S => n1, Y => 
                           TMP_1_1_port);
   MUX21_K_0_1 : MUX21_L_317 port map( A => A(2), B => A(1), S => n1, Y => 
                           TMP_1_2_port);
   MUX21_K_0_2 : MUX21_L_316 port map( A => A(3), B => A(2), S => n1, Y => 
                           TMP_1_3_port);
   MUX21_K_0_3 : MUX21_L_315 port map( A => A(4), B => A(3), S => n1, Y => 
                           TMP_1_4_port);
   MUX21_K_0_4 : MUX21_L_314 port map( A => A(5), B => A(4), S => n1, Y => 
                           TMP_1_5_port);
   MUX21_K_0_5 : MUX21_L_313 port map( A => A(6), B => A(5), S => n1, Y => 
                           TMP_1_6_port);
   MUX21_K_0_6 : MUX21_L_312 port map( A => A(7), B => A(6), S => n1, Y => 
                           TMP_1_7_port);
   MUX21_K_0_7 : MUX21_L_311 port map( A => A(8), B => A(7), S => n1, Y => 
                           TMP_1_8_port);
   MUX21_K_0_8 : MUX21_L_310 port map( A => A(9), B => A(8), S => n1, Y => 
                           TMP_1_9_port);
   MUX21_K_0_9 : MUX21_L_309 port map( A => A(10), B => A(9), S => n1, Y => 
                           TMP_1_10_port);
   MUX21_K_0_10 : MUX21_L_308 port map( A => A(11), B => A(10), S => n1, Y => 
                           TMP_1_11_port);
   MUX21_K_0_11 : MUX21_L_307 port map( A => A(12), B => A(11), S => n2, Y => 
                           TMP_1_12_port);
   MUX21_K_0_12 : MUX21_L_306 port map( A => A(13), B => A(12), S => n2, Y => 
                           TMP_1_13_port);
   MUX21_K_0_13 : MUX21_L_305 port map( A => A(14), B => A(13), S => n2, Y => 
                           TMP_1_14_port);
   MUX21_K_0_14 : MUX21_L_304 port map( A => A(15), B => A(14), S => n2, Y => 
                           TMP_1_15_port);
   MUX21_K_0_15 : MUX21_L_303 port map( A => A(16), B => A(15), S => n2, Y => 
                           TMP_1_16_port);
   MUX21_K_0_16 : MUX21_L_302 port map( A => A(17), B => A(16), S => n2, Y => 
                           TMP_1_17_port);
   MUX21_K_0_17 : MUX21_L_301 port map( A => A(18), B => A(17), S => n2, Y => 
                           TMP_1_18_port);
   MUX21_K_0_18 : MUX21_L_300 port map( A => A(19), B => A(18), S => n2, Y => 
                           TMP_1_19_port);
   MUX21_K_0_19 : MUX21_L_299 port map( A => A(20), B => A(19), S => n2, Y => 
                           TMP_1_20_port);
   MUX21_K_0_20 : MUX21_L_298 port map( A => A(21), B => A(20), S => n2, Y => 
                           TMP_1_21_port);
   MUX21_K_0_21 : MUX21_L_297 port map( A => A(22), B => A(21), S => n2, Y => 
                           TMP_1_22_port);
   MUX21_K_0_22 : MUX21_L_296 port map( A => A(23), B => A(22), S => n2, Y => 
                           TMP_1_23_port);
   MUX21_K_0_23 : MUX21_L_295 port map( A => A(24), B => A(23), S => n3, Y => 
                           TMP_1_24_port);
   MUX21_K_0_24 : MUX21_L_294 port map( A => A(25), B => A(24), S => n3, Y => 
                           TMP_1_25_port);
   MUX21_K_0_25 : MUX21_L_293 port map( A => A(26), B => A(25), S => n3, Y => 
                           TMP_1_26_port);
   MUX21_K_0_26 : MUX21_L_292 port map( A => A(27), B => A(26), S => n3, Y => 
                           TMP_1_27_port);
   MUX21_K_0_27 : MUX21_L_291 port map( A => A(28), B => A(27), S => n3, Y => 
                           TMP_1_28_port);
   MUX21_K_0_28 : MUX21_L_290 port map( A => A(29), B => A(28), S => n3, Y => 
                           TMP_1_29_port);
   MUX21_K_0_29 : MUX21_L_289 port map( A => A(30), B => A(29), S => n3, Y => 
                           TMP_1_30_port);
   MUX21_K_0_30 : MUX21_L_288 port map( A => A(31), B => A(30), S => n3, Y => 
                           TMP_1_31_port);
   MUX21_J_1_0 : MUX21_L_287 port map( A => TMP_1_0_port, B => X_Logic0_port, S
                           => n5, Y => TMP_2_0_port);
   MUX21_J_1_1 : MUX21_L_286 port map( A => TMP_1_1_port, B => X_Logic0_port, S
                           => n5, Y => TMP_2_1_port);
   MUX21_K_1_0 : MUX21_L_285 port map( A => TMP_1_2_port, B => TMP_1_0_port, S 
                           => n5, Y => TMP_2_2_port);
   MUX21_K_1_1 : MUX21_L_284 port map( A => TMP_1_3_port, B => TMP_1_1_port, S 
                           => n5, Y => TMP_2_3_port);
   MUX21_K_1_2 : MUX21_L_283 port map( A => TMP_1_4_port, B => TMP_1_2_port, S 
                           => n5, Y => TMP_2_4_port);
   MUX21_K_1_3 : MUX21_L_282 port map( A => TMP_1_5_port, B => TMP_1_3_port, S 
                           => n5, Y => TMP_2_5_port);
   MUX21_K_1_4 : MUX21_L_281 port map( A => TMP_1_6_port, B => TMP_1_4_port, S 
                           => n5, Y => TMP_2_6_port);
   MUX21_K_1_5 : MUX21_L_280 port map( A => TMP_1_7_port, B => TMP_1_5_port, S 
                           => n5, Y => TMP_2_7_port);
   MUX21_K_1_6 : MUX21_L_279 port map( A => TMP_1_8_port, B => TMP_1_6_port, S 
                           => n5, Y => TMP_2_8_port);
   MUX21_K_1_7 : MUX21_L_278 port map( A => TMP_1_9_port, B => TMP_1_7_port, S 
                           => n5, Y => TMP_2_9_port);
   MUX21_K_1_8 : MUX21_L_277 port map( A => TMP_1_10_port, B => TMP_1_8_port, S
                           => n5, Y => TMP_2_10_port);
   MUX21_K_1_9 : MUX21_L_276 port map( A => TMP_1_11_port, B => TMP_1_9_port, S
                           => n5, Y => TMP_2_11_port);
   MUX21_K_1_10 : MUX21_L_275 port map( A => TMP_1_12_port, B => TMP_1_10_port,
                           S => n6, Y => TMP_2_12_port);
   MUX21_K_1_11 : MUX21_L_274 port map( A => TMP_1_13_port, B => TMP_1_11_port,
                           S => n6, Y => TMP_2_13_port);
   MUX21_K_1_12 : MUX21_L_273 port map( A => TMP_1_14_port, B => TMP_1_12_port,
                           S => n6, Y => TMP_2_14_port);
   MUX21_K_1_13 : MUX21_L_272 port map( A => TMP_1_15_port, B => TMP_1_13_port,
                           S => n6, Y => TMP_2_15_port);
   MUX21_K_1_14 : MUX21_L_271 port map( A => TMP_1_16_port, B => TMP_1_14_port,
                           S => n6, Y => TMP_2_16_port);
   MUX21_K_1_15 : MUX21_L_270 port map( A => TMP_1_17_port, B => TMP_1_15_port,
                           S => n6, Y => TMP_2_17_port);
   MUX21_K_1_16 : MUX21_L_269 port map( A => TMP_1_18_port, B => TMP_1_16_port,
                           S => n6, Y => TMP_2_18_port);
   MUX21_K_1_17 : MUX21_L_268 port map( A => TMP_1_19_port, B => TMP_1_17_port,
                           S => n6, Y => TMP_2_19_port);
   MUX21_K_1_18 : MUX21_L_267 port map( A => TMP_1_20_port, B => TMP_1_18_port,
                           S => n6, Y => TMP_2_20_port);
   MUX21_K_1_19 : MUX21_L_266 port map( A => TMP_1_21_port, B => TMP_1_19_port,
                           S => n6, Y => TMP_2_21_port);
   MUX21_K_1_20 : MUX21_L_265 port map( A => TMP_1_22_port, B => TMP_1_20_port,
                           S => n6, Y => TMP_2_22_port);
   MUX21_K_1_21 : MUX21_L_264 port map( A => TMP_1_23_port, B => TMP_1_21_port,
                           S => n6, Y => TMP_2_23_port);
   MUX21_K_1_22 : MUX21_L_263 port map( A => TMP_1_24_port, B => TMP_1_22_port,
                           S => n7, Y => TMP_2_24_port);
   MUX21_K_1_23 : MUX21_L_262 port map( A => TMP_1_25_port, B => TMP_1_23_port,
                           S => n7, Y => TMP_2_25_port);
   MUX21_K_1_24 : MUX21_L_261 port map( A => TMP_1_26_port, B => TMP_1_24_port,
                           S => n7, Y => TMP_2_26_port);
   MUX21_K_1_25 : MUX21_L_260 port map( A => TMP_1_27_port, B => TMP_1_25_port,
                           S => n7, Y => TMP_2_27_port);
   MUX21_K_1_26 : MUX21_L_259 port map( A => TMP_1_28_port, B => TMP_1_26_port,
                           S => n7, Y => TMP_2_28_port);
   MUX21_K_1_27 : MUX21_L_258 port map( A => TMP_1_29_port, B => TMP_1_27_port,
                           S => n7, Y => TMP_2_29_port);
   MUX21_K_1_28 : MUX21_L_257 port map( A => TMP_1_30_port, B => TMP_1_28_port,
                           S => n7, Y => TMP_2_30_port);
   MUX21_K_1_29 : MUX21_L_256 port map( A => TMP_1_31_port, B => TMP_1_29_port,
                           S => n7, Y => TMP_2_31_port);
   MUX21_J_2_0 : MUX21_L_255 port map( A => TMP_2_0_port, B => X_Logic0_port, S
                           => n9, Y => TMP_3_0_port);
   MUX21_J_2_1 : MUX21_L_254 port map( A => TMP_2_1_port, B => X_Logic0_port, S
                           => n9, Y => TMP_3_1_port);
   MUX21_J_2_2 : MUX21_L_253 port map( A => TMP_2_2_port, B => X_Logic0_port, S
                           => n9, Y => TMP_3_2_port);
   MUX21_J_2_3 : MUX21_L_252 port map( A => TMP_2_3_port, B => X_Logic0_port, S
                           => n9, Y => TMP_3_3_port);
   MUX21_K_2_0 : MUX21_L_251 port map( A => TMP_2_4_port, B => TMP_2_0_port, S 
                           => n9, Y => TMP_3_4_port);
   MUX21_K_2_1 : MUX21_L_250 port map( A => TMP_2_5_port, B => TMP_2_1_port, S 
                           => n9, Y => TMP_3_5_port);
   MUX21_K_2_2 : MUX21_L_249 port map( A => TMP_2_6_port, B => TMP_2_2_port, S 
                           => n9, Y => TMP_3_6_port);
   MUX21_K_2_3 : MUX21_L_248 port map( A => TMP_2_7_port, B => TMP_2_3_port, S 
                           => n9, Y => TMP_3_7_port);
   MUX21_K_2_4 : MUX21_L_247 port map( A => TMP_2_8_port, B => TMP_2_4_port, S 
                           => n9, Y => TMP_3_8_port);
   MUX21_K_2_5 : MUX21_L_246 port map( A => TMP_2_9_port, B => TMP_2_5_port, S 
                           => n9, Y => TMP_3_9_port);
   MUX21_K_2_6 : MUX21_L_245 port map( A => TMP_2_10_port, B => TMP_2_6_port, S
                           => n9, Y => TMP_3_10_port);
   MUX21_K_2_7 : MUX21_L_244 port map( A => TMP_2_11_port, B => TMP_2_7_port, S
                           => n9, Y => TMP_3_11_port);
   MUX21_K_2_8 : MUX21_L_243 port map( A => TMP_2_12_port, B => TMP_2_8_port, S
                           => n10, Y => TMP_3_12_port);
   MUX21_K_2_9 : MUX21_L_242 port map( A => TMP_2_13_port, B => TMP_2_9_port, S
                           => n10, Y => TMP_3_13_port);
   MUX21_K_2_10 : MUX21_L_241 port map( A => TMP_2_14_port, B => TMP_2_10_port,
                           S => n10, Y => TMP_3_14_port);
   MUX21_K_2_11 : MUX21_L_240 port map( A => TMP_2_15_port, B => TMP_2_11_port,
                           S => n10, Y => TMP_3_15_port);
   MUX21_K_2_12 : MUX21_L_239 port map( A => TMP_2_16_port, B => TMP_2_12_port,
                           S => n10, Y => TMP_3_16_port);
   MUX21_K_2_13 : MUX21_L_238 port map( A => TMP_2_17_port, B => TMP_2_13_port,
                           S => n10, Y => TMP_3_17_port);
   MUX21_K_2_14 : MUX21_L_237 port map( A => TMP_2_18_port, B => TMP_2_14_port,
                           S => n10, Y => TMP_3_18_port);
   MUX21_K_2_15 : MUX21_L_236 port map( A => TMP_2_19_port, B => TMP_2_15_port,
                           S => n10, Y => TMP_3_19_port);
   MUX21_K_2_16 : MUX21_L_235 port map( A => TMP_2_20_port, B => TMP_2_16_port,
                           S => n10, Y => TMP_3_20_port);
   MUX21_K_2_17 : MUX21_L_234 port map( A => TMP_2_21_port, B => TMP_2_17_port,
                           S => n10, Y => TMP_3_21_port);
   MUX21_K_2_18 : MUX21_L_233 port map( A => TMP_2_22_port, B => TMP_2_18_port,
                           S => n10, Y => TMP_3_22_port);
   MUX21_K_2_19 : MUX21_L_232 port map( A => TMP_2_23_port, B => TMP_2_19_port,
                           S => n10, Y => TMP_3_23_port);
   MUX21_K_2_20 : MUX21_L_231 port map( A => TMP_2_24_port, B => TMP_2_20_port,
                           S => n11, Y => TMP_3_24_port);
   MUX21_K_2_21 : MUX21_L_230 port map( A => TMP_2_25_port, B => TMP_2_21_port,
                           S => n11, Y => TMP_3_25_port);
   MUX21_K_2_22 : MUX21_L_229 port map( A => TMP_2_26_port, B => TMP_2_22_port,
                           S => n11, Y => TMP_3_26_port);
   MUX21_K_2_23 : MUX21_L_228 port map( A => TMP_2_27_port, B => TMP_2_23_port,
                           S => n11, Y => TMP_3_27_port);
   MUX21_K_2_24 : MUX21_L_227 port map( A => TMP_2_28_port, B => TMP_2_24_port,
                           S => n11, Y => TMP_3_28_port);
   MUX21_K_2_25 : MUX21_L_226 port map( A => TMP_2_29_port, B => TMP_2_25_port,
                           S => n11, Y => TMP_3_29_port);
   MUX21_K_2_26 : MUX21_L_225 port map( A => TMP_2_30_port, B => TMP_2_26_port,
                           S => n11, Y => TMP_3_30_port);
   MUX21_K_2_27 : MUX21_L_224 port map( A => TMP_2_31_port, B => TMP_2_27_port,
                           S => n11, Y => TMP_3_31_port);
   MUX21_J_3_0 : MUX21_L_223 port map( A => TMP_3_0_port, B => X_Logic0_port, S
                           => n13, Y => TMP_4_0_port);
   MUX21_J_3_1 : MUX21_L_222 port map( A => TMP_3_1_port, B => X_Logic0_port, S
                           => n13, Y => TMP_4_1_port);
   MUX21_J_3_2 : MUX21_L_221 port map( A => TMP_3_2_port, B => X_Logic0_port, S
                           => n13, Y => TMP_4_2_port);
   MUX21_J_3_3 : MUX21_L_220 port map( A => TMP_3_3_port, B => X_Logic0_port, S
                           => n13, Y => TMP_4_3_port);
   MUX21_J_3_4 : MUX21_L_219 port map( A => TMP_3_4_port, B => X_Logic0_port, S
                           => n13, Y => TMP_4_4_port);
   MUX21_J_3_5 : MUX21_L_218 port map( A => TMP_3_5_port, B => X_Logic0_port, S
                           => n13, Y => TMP_4_5_port);
   MUX21_J_3_6 : MUX21_L_217 port map( A => TMP_3_6_port, B => X_Logic0_port, S
                           => n13, Y => TMP_4_6_port);
   MUX21_J_3_7 : MUX21_L_216 port map( A => TMP_3_7_port, B => X_Logic0_port, S
                           => n13, Y => TMP_4_7_port);
   MUX21_K_3_0 : MUX21_L_215 port map( A => TMP_3_8_port, B => TMP_3_0_port, S 
                           => n13, Y => TMP_4_8_port);
   MUX21_K_3_1 : MUX21_L_214 port map( A => TMP_3_9_port, B => TMP_3_1_port, S 
                           => n13, Y => TMP_4_9_port);
   MUX21_K_3_2 : MUX21_L_213 port map( A => TMP_3_10_port, B => TMP_3_2_port, S
                           => n13, Y => TMP_4_10_port);
   MUX21_K_3_3 : MUX21_L_212 port map( A => TMP_3_11_port, B => TMP_3_3_port, S
                           => n13, Y => TMP_4_11_port);
   MUX21_K_3_4 : MUX21_L_211 port map( A => TMP_3_12_port, B => TMP_3_4_port, S
                           => n14, Y => TMP_4_12_port);
   MUX21_K_3_5 : MUX21_L_210 port map( A => TMP_3_13_port, B => TMP_3_5_port, S
                           => n14, Y => TMP_4_13_port);
   MUX21_K_3_6 : MUX21_L_209 port map( A => TMP_3_14_port, B => TMP_3_6_port, S
                           => n14, Y => TMP_4_14_port);
   MUX21_K_3_7 : MUX21_L_208 port map( A => TMP_3_15_port, B => TMP_3_7_port, S
                           => n14, Y => TMP_4_15_port);
   MUX21_K_3_8 : MUX21_L_207 port map( A => TMP_3_16_port, B => TMP_3_8_port, S
                           => n14, Y => TMP_4_16_port);
   MUX21_K_3_9 : MUX21_L_206 port map( A => TMP_3_17_port, B => TMP_3_9_port, S
                           => n14, Y => TMP_4_17_port);
   MUX21_K_3_10 : MUX21_L_205 port map( A => TMP_3_18_port, B => TMP_3_10_port,
                           S => n14, Y => TMP_4_18_port);
   MUX21_K_3_11 : MUX21_L_204 port map( A => TMP_3_19_port, B => TMP_3_11_port,
                           S => n14, Y => TMP_4_19_port);
   MUX21_K_3_12 : MUX21_L_203 port map( A => TMP_3_20_port, B => TMP_3_12_port,
                           S => n14, Y => TMP_4_20_port);
   MUX21_K_3_13 : MUX21_L_202 port map( A => TMP_3_21_port, B => TMP_3_13_port,
                           S => n14, Y => TMP_4_21_port);
   MUX21_K_3_14 : MUX21_L_201 port map( A => TMP_3_22_port, B => TMP_3_14_port,
                           S => n14, Y => TMP_4_22_port);
   MUX21_K_3_15 : MUX21_L_200 port map( A => TMP_3_23_port, B => TMP_3_15_port,
                           S => n14, Y => TMP_4_23_port);
   MUX21_K_3_16 : MUX21_L_199 port map( A => TMP_3_24_port, B => TMP_3_16_port,
                           S => n15, Y => TMP_4_24_port);
   MUX21_K_3_17 : MUX21_L_198 port map( A => TMP_3_25_port, B => TMP_3_17_port,
                           S => n15, Y => TMP_4_25_port);
   MUX21_K_3_18 : MUX21_L_197 port map( A => TMP_3_26_port, B => TMP_3_18_port,
                           S => n15, Y => TMP_4_26_port);
   MUX21_K_3_19 : MUX21_L_196 port map( A => TMP_3_27_port, B => TMP_3_19_port,
                           S => n15, Y => TMP_4_27_port);
   MUX21_K_3_20 : MUX21_L_195 port map( A => TMP_3_28_port, B => TMP_3_20_port,
                           S => n15, Y => TMP_4_28_port);
   MUX21_K_3_21 : MUX21_L_194 port map( A => TMP_3_29_port, B => TMP_3_21_port,
                           S => n15, Y => TMP_4_29_port);
   MUX21_K_3_22 : MUX21_L_193 port map( A => TMP_3_30_port, B => TMP_3_22_port,
                           S => n15, Y => TMP_4_30_port);
   MUX21_K_3_23 : MUX21_L_192 port map( A => TMP_3_31_port, B => TMP_3_23_port,
                           S => n15, Y => TMP_4_31_port);
   MUX21_J_4_0 : MUX21_L_191 port map( A => TMP_4_0_port, B => X_Logic0_port, S
                           => n17, Y => Y(0));
   MUX21_J_4_1 : MUX21_L_190 port map( A => TMP_4_1_port, B => X_Logic0_port, S
                           => n17, Y => Y(1));
   MUX21_J_4_2 : MUX21_L_189 port map( A => TMP_4_2_port, B => X_Logic0_port, S
                           => n17, Y => Y(2));
   MUX21_J_4_3 : MUX21_L_188 port map( A => TMP_4_3_port, B => X_Logic0_port, S
                           => n17, Y => Y(3));
   MUX21_J_4_4 : MUX21_L_187 port map( A => TMP_4_4_port, B => X_Logic0_port, S
                           => n17, Y => Y(4));
   MUX21_J_4_5 : MUX21_L_186 port map( A => TMP_4_5_port, B => X_Logic0_port, S
                           => n17, Y => Y(5));
   MUX21_J_4_6 : MUX21_L_185 port map( A => TMP_4_6_port, B => X_Logic0_port, S
                           => n17, Y => Y(6));
   MUX21_J_4_7 : MUX21_L_184 port map( A => TMP_4_7_port, B => X_Logic0_port, S
                           => n17, Y => Y(7));
   MUX21_J_4_8 : MUX21_L_183 port map( A => TMP_4_8_port, B => X_Logic0_port, S
                           => n17, Y => Y(8));
   MUX21_J_4_9 : MUX21_L_182 port map( A => TMP_4_9_port, B => X_Logic0_port, S
                           => n17, Y => Y(9));
   MUX21_J_4_10 : MUX21_L_181 port map( A => TMP_4_10_port, B => X_Logic0_port,
                           S => n17, Y => Y(10));
   MUX21_J_4_11 : MUX21_L_180 port map( A => TMP_4_11_port, B => X_Logic0_port,
                           S => n17, Y => Y(11));
   MUX21_J_4_12 : MUX21_L_179 port map( A => TMP_4_12_port, B => X_Logic0_port,
                           S => n18, Y => Y(12));
   MUX21_J_4_13 : MUX21_L_178 port map( A => TMP_4_13_port, B => X_Logic0_port,
                           S => n18, Y => Y(13));
   MUX21_J_4_14 : MUX21_L_177 port map( A => TMP_4_14_port, B => X_Logic0_port,
                           S => n18, Y => Y(14));
   MUX21_J_4_15 : MUX21_L_176 port map( A => TMP_4_15_port, B => X_Logic0_port,
                           S => n18, Y => Y(15));
   MUX21_K_4_0 : MUX21_L_175 port map( A => TMP_4_16_port, B => TMP_4_0_port, S
                           => n18, Y => Y(16));
   MUX21_K_4_1 : MUX21_L_174 port map( A => TMP_4_17_port, B => TMP_4_1_port, S
                           => n18, Y => Y(17));
   MUX21_K_4_2 : MUX21_L_173 port map( A => TMP_4_18_port, B => TMP_4_2_port, S
                           => n18, Y => Y(18));
   MUX21_K_4_3 : MUX21_L_172 port map( A => TMP_4_19_port, B => TMP_4_3_port, S
                           => n18, Y => Y(19));
   MUX21_K_4_4 : MUX21_L_171 port map( A => TMP_4_20_port, B => TMP_4_4_port, S
                           => n18, Y => Y(20));
   MUX21_K_4_5 : MUX21_L_170 port map( A => TMP_4_21_port, B => TMP_4_5_port, S
                           => n18, Y => Y(21));
   MUX21_K_4_6 : MUX21_L_169 port map( A => TMP_4_22_port, B => TMP_4_6_port, S
                           => n18, Y => Y(22));
   MUX21_K_4_7 : MUX21_L_168 port map( A => TMP_4_23_port, B => TMP_4_7_port, S
                           => n18, Y => Y(23));
   MUX21_K_4_8 : MUX21_L_167 port map( A => TMP_4_24_port, B => TMP_4_8_port, S
                           => n19, Y => Y(24));
   MUX21_K_4_9 : MUX21_L_166 port map( A => TMP_4_25_port, B => TMP_4_9_port, S
                           => n19, Y => Y(25));
   MUX21_K_4_10 : MUX21_L_165 port map( A => TMP_4_26_port, B => TMP_4_10_port,
                           S => n19, Y => Y(26));
   MUX21_K_4_11 : MUX21_L_164 port map( A => TMP_4_27_port, B => TMP_4_11_port,
                           S => n19, Y => Y(27));
   MUX21_K_4_12 : MUX21_L_163 port map( A => TMP_4_28_port, B => TMP_4_12_port,
                           S => n19, Y => Y(28));
   MUX21_K_4_13 : MUX21_L_162 port map( A => TMP_4_29_port, B => TMP_4_13_port,
                           S => n19, Y => Y(29));
   MUX21_K_4_14 : MUX21_L_161 port map( A => TMP_4_30_port, B => TMP_4_14_port,
                           S => n19, Y => Y(30));
   MUX21_K_4_15 : MUX21_L_160 port map( A => TMP_4_31_port, B => TMP_4_15_port,
                           S => n19, Y => Y(31));
   U2 : BUF_X1 port map( A => n12, Z => n9);
   U3 : BUF_X1 port map( A => n12, Z => n10);
   U4 : BUF_X1 port map( A => n20, Z => n19);
   U5 : BUF_X1 port map( A => n16, Z => n15);
   U6 : BUF_X1 port map( A => n16, Z => n14);
   U7 : BUF_X1 port map( A => B(3), Z => n16);
   U8 : BUF_X1 port map( A => B(2), Z => n12);
   U9 : BUF_X1 port map( A => B(4), Z => n20);
   U10 : BUF_X1 port map( A => B(1), Z => n8);
   U11 : BUF_X1 port map( A => B(0), Z => n4);
   U12 : BUF_X1 port map( A => n4, Z => n1);
   U13 : BUF_X1 port map( A => n4, Z => n2);
   U14 : BUF_X1 port map( A => n8, Z => n5);
   U15 : BUF_X1 port map( A => n8, Z => n6);
   U16 : BUF_X1 port map( A => n16, Z => n13);
   U17 : BUF_X1 port map( A => n20, Z => n17);
   U18 : BUF_X1 port map( A => n20, Z => n18);
   U19 : BUF_X1 port map( A => n4, Z => n3);
   U20 : BUF_X1 port map( A => n8, Z => n7);
   U21 : BUF_X1 port map( A => n12, Z => n11);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BOOTH_MULTIPLIER_N32 is

   port( A, B : in std_logic_vector (15 downto 0);  P : out std_logic_vector 
         (31 downto 0));

end BOOTH_MULTIPLIER_N32;

architecture SYN_STRUCTURAL of BOOTH_MULTIPLIER_N32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component RCA_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component MUX81_N32_0
      port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component RCA_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component MUX81_N32_1
      port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component RCA_N32_2
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component MUX81_N32_2
      port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX81_N32_3
      port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component BOOTH_ENCODER_N16
      port( B : in std_logic_vector (15 downto 0);  Bo : out std_logic_vector 
            (23 downto 0));
   end component;
   
   signal X_Logic0_port, Bo_signal_11_port, Bo_signal_10_port, Bo_signal_9_port
      , Bo_signal_8_port, Bo_signal_7_port, Bo_signal_6_port, Bo_signal_5_port,
      Bo_signal_4_port, Bo_signal_3_port, Bo_signal_2_port, Bo_signal_1_port, 
      Bo_signal_0_port, aMatrix_15_31_port, aMatrix_15_22_port, 
      aMatrix_15_21_port, aMatrix_15_20_port, aMatrix_15_19_port, 
      aMatrix_15_18_port, aMatrix_15_17_port, aMatrix_15_16_port, 
      aMatrix_15_15_port, aMatrix_15_14_port, aMatrix_15_13_port, 
      aMatrix_15_12_port, aMatrix_15_11_port, aMatrix_15_10_port, 
      aMatrix_15_9_port, aMatrix_15_8_port, aMatrix_15_0_port, 
      aMatrix_13_31_port, aMatrix_13_21_port, aMatrix_13_20_port, 
      aMatrix_13_19_port, aMatrix_13_18_port, aMatrix_13_17_port, 
      aMatrix_13_16_port, aMatrix_13_15_port, aMatrix_13_14_port, 
      aMatrix_13_13_port, aMatrix_13_12_port, aMatrix_13_11_port, 
      aMatrix_13_10_port, aMatrix_13_9_port, aMatrix_13_8_port, 
      aMatrix_13_7_port, aMatrix_13_0_port, aMatrix_11_31_port, 
      aMatrix_11_20_port, aMatrix_11_19_port, aMatrix_11_18_port, 
      aMatrix_11_17_port, aMatrix_11_16_port, aMatrix_11_15_port, 
      aMatrix_11_14_port, aMatrix_11_13_port, aMatrix_11_12_port, 
      aMatrix_11_11_port, aMatrix_11_10_port, aMatrix_11_9_port, 
      aMatrix_11_8_port, aMatrix_11_7_port, aMatrix_11_6_port, 
      aMatrix_11_0_port, aMatrix_9_31_port, aMatrix_9_19_port, 
      aMatrix_9_18_port, aMatrix_9_17_port, aMatrix_9_16_port, 
      aMatrix_9_15_port, aMatrix_9_14_port, aMatrix_9_13_port, 
      aMatrix_9_12_port, aMatrix_9_11_port, aMatrix_9_10_port, aMatrix_9_9_port
      , aMatrix_9_8_port, aMatrix_9_7_port, aMatrix_9_6_port, aMatrix_9_5_port,
      aMatrix_9_0_port, aMatrix_7_31_port, aMatrix_7_18_port, aMatrix_7_17_port
      , aMatrix_7_16_port, aMatrix_7_15_port, aMatrix_7_14_port, 
      aMatrix_7_13_port, aMatrix_7_12_port, aMatrix_7_11_port, 
      aMatrix_7_10_port, aMatrix_7_9_port, aMatrix_7_8_port, aMatrix_7_7_port, 
      aMatrix_7_6_port, aMatrix_7_5_port, aMatrix_7_4_port, aMatrix_7_0_port, 
      aMatrix_5_31_port, aMatrix_5_17_port, aMatrix_5_16_port, 
      aMatrix_5_15_port, aMatrix_5_14_port, aMatrix_5_13_port, 
      aMatrix_5_12_port, aMatrix_5_11_port, aMatrix_5_10_port, aMatrix_5_9_port
      , aMatrix_5_8_port, aMatrix_5_7_port, aMatrix_5_6_port, aMatrix_5_5_port,
      aMatrix_5_4_port, aMatrix_5_3_port, aMatrix_5_0_port, aMatrix_3_31_port, 
      aMatrix_3_16_port, aMatrix_3_15_port, aMatrix_3_14_port, 
      aMatrix_3_13_port, aMatrix_3_12_port, aMatrix_3_11_port, 
      aMatrix_3_10_port, aMatrix_3_9_port, aMatrix_3_8_port, aMatrix_3_7_port, 
      aMatrix_3_6_port, aMatrix_3_5_port, aMatrix_3_4_port, aMatrix_3_3_port, 
      aMatrix_3_2_port, aMatrix_3_0_port, aMatrix_1_31_port, aMatrix_1_15_port,
      aMatrix_1_14_port, aMatrix_1_13_port, aMatrix_1_12_port, 
      aMatrix_1_11_port, aMatrix_1_10_port, aMatrix_1_9_port, aMatrix_1_8_port,
      aMatrix_1_7_port, aMatrix_1_6_port, aMatrix_1_5_port, aMatrix_1_4_port, 
      aMatrix_1_3_port, aMatrix_1_2_port, aMatrix_1_1_port, 
      aEncMatrix_3_31_port, aEncMatrix_3_30_port, aEncMatrix_3_29_port, 
      aEncMatrix_3_28_port, aEncMatrix_3_27_port, aEncMatrix_3_26_port, 
      aEncMatrix_3_25_port, aEncMatrix_3_24_port, aEncMatrix_3_23_port, 
      aEncMatrix_3_22_port, aEncMatrix_3_21_port, aEncMatrix_3_20_port, 
      aEncMatrix_3_19_port, aEncMatrix_3_18_port, aEncMatrix_3_17_port, 
      aEncMatrix_3_16_port, aEncMatrix_3_15_port, aEncMatrix_3_14_port, 
      aEncMatrix_3_13_port, aEncMatrix_3_12_port, aEncMatrix_3_11_port, 
      aEncMatrix_3_10_port, aEncMatrix_3_9_port, aEncMatrix_3_8_port, 
      aEncMatrix_3_7_port, aEncMatrix_3_6_port, aEncMatrix_3_5_port, 
      aEncMatrix_3_4_port, aEncMatrix_3_3_port, aEncMatrix_3_2_port, 
      aEncMatrix_3_1_port, aEncMatrix_3_0_port, aEncMatrix_2_31_port, 
      aEncMatrix_2_30_port, aEncMatrix_2_29_port, aEncMatrix_2_28_port, 
      aEncMatrix_2_27_port, aEncMatrix_2_26_port, aEncMatrix_2_25_port, 
      aEncMatrix_2_24_port, aEncMatrix_2_23_port, aEncMatrix_2_22_port, 
      aEncMatrix_2_21_port, aEncMatrix_2_20_port, aEncMatrix_2_19_port, 
      aEncMatrix_2_18_port, aEncMatrix_2_17_port, aEncMatrix_2_16_port, 
      aEncMatrix_2_15_port, aEncMatrix_2_14_port, aEncMatrix_2_13_port, 
      aEncMatrix_2_12_port, aEncMatrix_2_11_port, aEncMatrix_2_10_port, 
      aEncMatrix_2_9_port, aEncMatrix_2_8_port, aEncMatrix_2_7_port, 
      aEncMatrix_2_6_port, aEncMatrix_2_5_port, aEncMatrix_2_4_port, 
      aEncMatrix_2_3_port, aEncMatrix_2_2_port, aEncMatrix_2_1_port, 
      aEncMatrix_2_0_port, aEncMatrix_1_31_port, aEncMatrix_1_30_port, 
      aEncMatrix_1_29_port, aEncMatrix_1_28_port, aEncMatrix_1_27_port, 
      aEncMatrix_1_26_port, aEncMatrix_1_25_port, aEncMatrix_1_24_port, 
      aEncMatrix_1_23_port, aEncMatrix_1_22_port, aEncMatrix_1_21_port, 
      aEncMatrix_1_20_port, aEncMatrix_1_19_port, aEncMatrix_1_18_port, 
      aEncMatrix_1_17_port, aEncMatrix_1_16_port, aEncMatrix_1_15_port, 
      aEncMatrix_1_14_port, aEncMatrix_1_13_port, aEncMatrix_1_12_port, 
      aEncMatrix_1_11_port, aEncMatrix_1_10_port, aEncMatrix_1_9_port, 
      aEncMatrix_1_8_port, aEncMatrix_1_7_port, aEncMatrix_1_6_port, 
      aEncMatrix_1_5_port, aEncMatrix_1_4_port, aEncMatrix_1_3_port, 
      aEncMatrix_1_2_port, aEncMatrix_1_1_port, aEncMatrix_1_0_port, 
      aEncMatrix_0_31_port, aEncMatrix_0_30_port, aEncMatrix_0_29_port, 
      aEncMatrix_0_28_port, aEncMatrix_0_27_port, aEncMatrix_0_26_port, 
      aEncMatrix_0_25_port, aEncMatrix_0_24_port, aEncMatrix_0_23_port, 
      aEncMatrix_0_22_port, aEncMatrix_0_21_port, aEncMatrix_0_20_port, 
      aEncMatrix_0_19_port, aEncMatrix_0_18_port, aEncMatrix_0_17_port, 
      aEncMatrix_0_16_port, aEncMatrix_0_15_port, aEncMatrix_0_14_port, 
      aEncMatrix_0_13_port, aEncMatrix_0_12_port, aEncMatrix_0_11_port, 
      aEncMatrix_0_10_port, aEncMatrix_0_9_port, aEncMatrix_0_8_port, 
      aEncMatrix_0_7_port, aEncMatrix_0_6_port, aEncMatrix_0_5_port, 
      aEncMatrix_0_4_port, aEncMatrix_0_3_port, aEncMatrix_0_2_port, 
      aEncMatrix_0_1_port, aEncMatrix_0_0_port, pSumMatrix_1_31_port, 
      pSumMatrix_1_30_port, pSumMatrix_1_29_port, pSumMatrix_1_28_port, 
      pSumMatrix_1_27_port, pSumMatrix_1_26_port, pSumMatrix_1_25_port, 
      pSumMatrix_1_24_port, pSumMatrix_1_23_port, pSumMatrix_1_22_port, 
      pSumMatrix_1_21_port, pSumMatrix_1_20_port, pSumMatrix_1_19_port, 
      pSumMatrix_1_18_port, pSumMatrix_1_17_port, pSumMatrix_1_16_port, 
      pSumMatrix_1_15_port, pSumMatrix_1_14_port, pSumMatrix_1_13_port, 
      pSumMatrix_1_12_port, pSumMatrix_1_11_port, pSumMatrix_1_10_port, 
      pSumMatrix_1_9_port, pSumMatrix_1_8_port, pSumMatrix_1_7_port, 
      pSumMatrix_1_6_port, pSumMatrix_1_5_port, pSumMatrix_1_4_port, 
      pSumMatrix_1_3_port, pSumMatrix_1_2_port, pSumMatrix_1_1_port, 
      pSumMatrix_1_0_port, pSumMatrix_0_31_port, pSumMatrix_0_30_port, 
      pSumMatrix_0_29_port, pSumMatrix_0_28_port, pSumMatrix_0_27_port, 
      pSumMatrix_0_26_port, pSumMatrix_0_25_port, pSumMatrix_0_24_port, 
      pSumMatrix_0_23_port, pSumMatrix_0_22_port, pSumMatrix_0_21_port, 
      pSumMatrix_0_20_port, pSumMatrix_0_19_port, pSumMatrix_0_18_port, 
      pSumMatrix_0_17_port, pSumMatrix_0_16_port, pSumMatrix_0_15_port, 
      pSumMatrix_0_14_port, pSumMatrix_0_13_port, pSumMatrix_0_12_port, 
      pSumMatrix_0_11_port, pSumMatrix_0_10_port, pSumMatrix_0_9_port, 
      pSumMatrix_0_8_port, pSumMatrix_0_7_port, pSumMatrix_0_6_port, 
      pSumMatrix_0_5_port, pSumMatrix_0_4_port, pSumMatrix_0_3_port, 
      pSumMatrix_0_2_port, pSumMatrix_0_1_port, pSumMatrix_0_0_port, 
      add_92_G8_carry_9_port, add_92_G8_carry_10_port, add_92_G8_carry_11_port,
      add_92_G8_carry_12_port, add_92_G8_carry_13_port, add_92_G8_carry_14_port
      , add_92_G8_carry_15_port, add_92_G8_carry_16_port, 
      add_92_G8_carry_17_port, add_92_G8_carry_18_port, add_92_G8_carry_19_port
      , add_92_G8_carry_20_port, add_92_G8_carry_21_port, 
      add_92_G8_carry_22_port, add_92_G7_carry_8_port, add_92_G7_carry_9_port, 
      add_92_G7_carry_10_port, add_92_G7_carry_11_port, add_92_G7_carry_12_port
      , add_92_G7_carry_13_port, add_92_G7_carry_14_port, 
      add_92_G7_carry_15_port, add_92_G7_carry_16_port, add_92_G7_carry_17_port
      , add_92_G7_carry_18_port, add_92_G7_carry_19_port, 
      add_92_G7_carry_20_port, add_92_G7_carry_21_port, add_92_G6_carry_7_port,
      add_92_G6_carry_8_port, add_92_G6_carry_9_port, add_92_G6_carry_10_port, 
      add_92_G6_carry_11_port, add_92_G6_carry_12_port, add_92_G6_carry_13_port
      , add_92_G6_carry_14_port, add_92_G6_carry_15_port, 
      add_92_G6_carry_16_port, add_92_G6_carry_17_port, add_92_G6_carry_18_port
      , add_92_G6_carry_19_port, add_92_G6_carry_20_port, 
      add_92_G5_carry_6_port, add_92_G5_carry_7_port, add_92_G5_carry_8_port, 
      add_92_G5_carry_9_port, add_92_G5_carry_10_port, add_92_G5_carry_11_port,
      add_92_G5_carry_12_port, add_92_G5_carry_13_port, add_92_G5_carry_14_port
      , add_92_G5_carry_15_port, add_92_G5_carry_16_port, 
      add_92_G5_carry_17_port, add_92_G5_carry_18_port, add_92_G5_carry_19_port
      , add_92_G4_carry_5_port, add_92_G4_carry_6_port, add_92_G4_carry_7_port,
      add_92_G4_carry_8_port, add_92_G4_carry_9_port, add_92_G4_carry_10_port, 
      add_92_G4_carry_11_port, add_92_G4_carry_12_port, add_92_G4_carry_13_port
      , add_92_G4_carry_14_port, add_92_G4_carry_15_port, 
      add_92_G4_carry_16_port, add_92_G4_carry_17_port, add_92_G4_carry_18_port
      , add_92_G3_carry_4_port, add_92_G3_carry_5_port, add_92_G3_carry_6_port,
      add_92_G3_carry_7_port, add_92_G3_carry_8_port, add_92_G3_carry_9_port, 
      add_92_G3_carry_10_port, add_92_G3_carry_11_port, add_92_G3_carry_12_port
      , add_92_G3_carry_13_port, add_92_G3_carry_14_port, 
      add_92_G3_carry_15_port, add_92_G3_carry_16_port, add_92_G3_carry_17_port
      , add_92_G2_carry_3_port, add_92_G2_carry_4_port, add_92_G2_carry_5_port,
      add_92_G2_carry_6_port, add_92_G2_carry_7_port, add_92_G2_carry_8_port, 
      add_92_G2_carry_9_port, add_92_G2_carry_10_port, add_92_G2_carry_11_port,
      add_92_G2_carry_12_port, add_92_G2_carry_13_port, add_92_G2_carry_14_port
      , add_92_G2_carry_15_port, add_92_G2_carry_16_port, add_92_carry_2_port, 
      add_92_carry_3_port, add_92_carry_4_port, add_92_carry_5_port, 
      add_92_carry_6_port, add_92_carry_7_port, add_92_carry_8_port, 
      add_92_carry_9_port, add_92_carry_10_port, add_92_carry_11_port, 
      add_92_carry_12_port, add_92_carry_13_port, add_92_carry_14_port, 
      add_92_carry_15_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   B_INSTANCE : BOOTH_ENCODER_N16 port map( B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           Bo(23) => n_1258, Bo(22) => n_1259, Bo(21) => n_1260
                           , Bo(20) => n_1261, Bo(19) => n_1262, Bo(18) => 
                           n_1263, Bo(17) => n_1264, Bo(16) => n_1265, Bo(15) 
                           => n_1266, Bo(14) => n_1267, Bo(13) => n_1268, 
                           Bo(12) => n_1269, Bo(11) => Bo_signal_11_port, 
                           Bo(10) => Bo_signal_10_port, Bo(9) => 
                           Bo_signal_9_port, Bo(8) => Bo_signal_8_port, Bo(7) 
                           => Bo_signal_7_port, Bo(6) => Bo_signal_6_port, 
                           Bo(5) => Bo_signal_5_port, Bo(4) => Bo_signal_4_port
                           , Bo(3) => Bo_signal_3_port, Bo(2) => 
                           Bo_signal_2_port, Bo(1) => Bo_signal_1_port, Bo(0) 
                           => Bo_signal_0_port);
   FIRST_MUX : MUX81_N32_3 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => n21, B(30) => n21, B(29) => 
                           n21, B(28) => n21, B(27) => n21, B(26) => n21, B(25)
                           => n21, B(24) => n21, B(23) => n21, B(22) => n21, 
                           B(21) => n21, B(20) => n21, B(19) => n20, B(18) => 
                           n21, B(17) => A(15), B(16) => n19, B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => n2
                           , B(0) => A(0), C(31) => aMatrix_1_31_port, C(30) =>
                           aMatrix_1_31_port, C(29) => aMatrix_1_31_port, C(28)
                           => aMatrix_1_31_port, C(27) => aMatrix_1_31_port, 
                           C(26) => aMatrix_1_31_port, C(25) => 
                           aMatrix_1_31_port, C(24) => aMatrix_1_31_port, C(23)
                           => aMatrix_1_31_port, C(22) => aMatrix_1_31_port, 
                           C(21) => aMatrix_1_31_port, C(20) => 
                           aMatrix_1_31_port, C(19) => aMatrix_1_31_port, C(18)
                           => aMatrix_1_31_port, C(17) => aMatrix_1_31_port, 
                           C(16) => aMatrix_1_31_port, C(15) => 
                           aMatrix_1_15_port, C(14) => aMatrix_1_14_port, C(13)
                           => aMatrix_1_13_port, C(12) => aMatrix_1_12_port, 
                           C(11) => aMatrix_1_11_port, C(10) => 
                           aMatrix_1_10_port, C(9) => aMatrix_1_9_port, C(8) =>
                           aMatrix_1_8_port, C(7) => aMatrix_1_7_port, C(6) => 
                           aMatrix_1_6_port, C(5) => aMatrix_1_5_port, C(4) => 
                           aMatrix_1_4_port, C(3) => aMatrix_1_3_port, C(2) => 
                           aMatrix_1_2_port, C(1) => aMatrix_1_1_port, C(0) => 
                           A(0), D(31) => n19, D(30) => n20, D(29) => n21, 
                           D(28) => A(15), D(27) => n17, D(26) => n20, D(25) =>
                           n18, D(24) => n20, D(23) => n20, D(22) => n20, D(21)
                           => n20, D(20) => n20, D(19) => n20, D(18) => n20, 
                           D(17) => n20, D(16) => n20, D(15) => A(14), D(14) =>
                           A(13), D(13) => A(12), D(12) => A(11), D(11) => 
                           A(10), D(10) => A(9), D(9) => A(8), D(8) => A(7), 
                           D(7) => A(6), D(6) => A(5), D(5) => A(4), D(4) => 
                           A(3), D(3) => A(2), D(2) => n2, D(1) => A(0), D(0) 
                           => X_Logic0_port, E(31) => aMatrix_3_31_port, E(30) 
                           => aMatrix_3_31_port, E(29) => aMatrix_3_31_port, 
                           E(28) => aMatrix_3_31_port, E(27) => 
                           aMatrix_3_31_port, E(26) => aMatrix_3_31_port, E(25)
                           => aMatrix_3_31_port, E(24) => aMatrix_3_31_port, 
                           E(23) => aMatrix_3_31_port, E(22) => 
                           aMatrix_3_31_port, E(21) => aMatrix_3_31_port, E(20)
                           => aMatrix_3_31_port, E(19) => aMatrix_3_31_port, 
                           E(18) => aMatrix_3_31_port, E(17) => 
                           aMatrix_3_31_port, E(16) => aMatrix_3_16_port, E(15)
                           => aMatrix_3_15_port, E(14) => aMatrix_3_14_port, 
                           E(13) => aMatrix_3_13_port, E(12) => 
                           aMatrix_3_12_port, E(11) => aMatrix_3_11_port, E(10)
                           => aMatrix_3_10_port, E(9) => aMatrix_3_9_port, E(8)
                           => aMatrix_3_8_port, E(7) => aMatrix_3_7_port, E(6) 
                           => aMatrix_3_6_port, E(5) => aMatrix_3_5_port, E(4) 
                           => aMatrix_3_4_port, E(3) => aMatrix_3_3_port, E(2) 
                           => aMatrix_3_2_port, E(1) => A(0), E(0) => 
                           aMatrix_3_0_port, F(31) => X_Logic0_port, F(30) => 
                           X_Logic0_port, F(29) => X_Logic0_port, F(28) => 
                           X_Logic0_port, F(27) => X_Logic0_port, F(26) => 
                           X_Logic0_port, F(25) => X_Logic0_port, F(24) => 
                           X_Logic0_port, F(23) => X_Logic0_port, F(22) => 
                           X_Logic0_port, F(21) => X_Logic0_port, F(20) => 
                           X_Logic0_port, F(19) => X_Logic0_port, F(18) => 
                           X_Logic0_port, F(17) => X_Logic0_port, F(16) => 
                           X_Logic0_port, F(15) => X_Logic0_port, F(14) => 
                           X_Logic0_port, F(13) => X_Logic0_port, F(12) => 
                           X_Logic0_port, F(11) => X_Logic0_port, F(10) => 
                           X_Logic0_port, F(9) => X_Logic0_port, F(8) => 
                           X_Logic0_port, F(7) => X_Logic0_port, F(6) => 
                           X_Logic0_port, F(5) => X_Logic0_port, F(4) => 
                           X_Logic0_port, F(3) => X_Logic0_port, F(2) => 
                           X_Logic0_port, F(1) => X_Logic0_port, F(0) => 
                           X_Logic0_port, G(31) => X_Logic0_port, G(30) => 
                           X_Logic0_port, G(29) => X_Logic0_port, G(28) => 
                           X_Logic0_port, G(27) => X_Logic0_port, G(26) => 
                           X_Logic0_port, G(25) => X_Logic0_port, G(24) => 
                           X_Logic0_port, G(23) => X_Logic0_port, G(22) => 
                           X_Logic0_port, G(21) => X_Logic0_port, G(20) => 
                           X_Logic0_port, G(19) => X_Logic0_port, G(18) => 
                           X_Logic0_port, G(17) => X_Logic0_port, G(16) => 
                           X_Logic0_port, G(15) => X_Logic0_port, G(14) => 
                           X_Logic0_port, G(13) => X_Logic0_port, G(12) => 
                           X_Logic0_port, G(11) => X_Logic0_port, G(10) => 
                           X_Logic0_port, G(9) => X_Logic0_port, G(8) => 
                           X_Logic0_port, G(7) => X_Logic0_port, G(6) => 
                           X_Logic0_port, G(5) => X_Logic0_port, G(4) => 
                           X_Logic0_port, G(3) => X_Logic0_port, G(2) => 
                           X_Logic0_port, G(1) => X_Logic0_port, G(0) => 
                           X_Logic0_port, H(31) => X_Logic0_port, H(30) => 
                           X_Logic0_port, H(29) => X_Logic0_port, H(28) => 
                           X_Logic0_port, H(27) => X_Logic0_port, H(26) => 
                           X_Logic0_port, H(25) => X_Logic0_port, H(24) => 
                           X_Logic0_port, H(23) => X_Logic0_port, H(22) => 
                           X_Logic0_port, H(21) => X_Logic0_port, H(20) => 
                           X_Logic0_port, H(19) => X_Logic0_port, H(18) => 
                           X_Logic0_port, H(17) => X_Logic0_port, H(16) => 
                           X_Logic0_port, H(15) => X_Logic0_port, H(14) => 
                           X_Logic0_port, H(13) => X_Logic0_port, H(12) => 
                           X_Logic0_port, H(11) => X_Logic0_port, H(10) => 
                           X_Logic0_port, H(9) => X_Logic0_port, H(8) => 
                           X_Logic0_port, H(7) => X_Logic0_port, H(6) => 
                           X_Logic0_port, H(5) => X_Logic0_port, H(4) => 
                           X_Logic0_port, H(3) => X_Logic0_port, H(2) => 
                           X_Logic0_port, H(1) => X_Logic0_port, H(0) => 
                           X_Logic0_port, S(2) => Bo_signal_2_port, S(1) => 
                           Bo_signal_1_port, S(0) => Bo_signal_0_port, Y(31) =>
                           aEncMatrix_0_31_port, Y(30) => aEncMatrix_0_30_port,
                           Y(29) => aEncMatrix_0_29_port, Y(28) => 
                           aEncMatrix_0_28_port, Y(27) => aEncMatrix_0_27_port,
                           Y(26) => aEncMatrix_0_26_port, Y(25) => 
                           aEncMatrix_0_25_port, Y(24) => aEncMatrix_0_24_port,
                           Y(23) => aEncMatrix_0_23_port, Y(22) => 
                           aEncMatrix_0_22_port, Y(21) => aEncMatrix_0_21_port,
                           Y(20) => aEncMatrix_0_20_port, Y(19) => 
                           aEncMatrix_0_19_port, Y(18) => aEncMatrix_0_18_port,
                           Y(17) => aEncMatrix_0_17_port, Y(16) => 
                           aEncMatrix_0_16_port, Y(15) => aEncMatrix_0_15_port,
                           Y(14) => aEncMatrix_0_14_port, Y(13) => 
                           aEncMatrix_0_13_port, Y(12) => aEncMatrix_0_12_port,
                           Y(11) => aEncMatrix_0_11_port, Y(10) => 
                           aEncMatrix_0_10_port, Y(9) => aEncMatrix_0_9_port, 
                           Y(8) => aEncMatrix_0_8_port, Y(7) => 
                           aEncMatrix_0_7_port, Y(6) => aEncMatrix_0_6_port, 
                           Y(5) => aEncMatrix_0_5_port, Y(4) => 
                           aEncMatrix_0_4_port, Y(3) => aEncMatrix_0_3_port, 
                           Y(2) => aEncMatrix_0_2_port, Y(1) => 
                           aEncMatrix_0_1_port, Y(0) => aEncMatrix_0_0_port);
   MUXES_1 : MUX81_N32_2 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => n19, B(30) => n19, B(29) => 
                           n19, B(28) => n19, B(27) => n19, B(26) => n18, B(25)
                           => n18, B(24) => n18, B(23) => n18, B(22) => n18, 
                           B(21) => n18, B(20) => n18, B(19) => n18, B(18) => 
                           n18, B(17) => n18, B(16) => A(14), B(15) => A(13), 
                           B(14) => A(12), B(13) => A(11), B(12) => A(10), 
                           B(11) => A(9), B(10) => A(8), B(9) => A(7), B(8) => 
                           A(6), B(7) => A(5), B(6) => A(4), B(5) => A(3), B(4)
                           => A(2), B(3) => n2, B(2) => A(0), B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => 
                           aMatrix_5_31_port, C(30) => aMatrix_5_31_port, C(29)
                           => aMatrix_5_31_port, C(28) => aMatrix_5_31_port, 
                           C(27) => aMatrix_5_31_port, C(26) => 
                           aMatrix_5_31_port, C(25) => aMatrix_5_31_port, C(24)
                           => aMatrix_5_31_port, C(23) => aMatrix_5_31_port, 
                           C(22) => aMatrix_5_31_port, C(21) => 
                           aMatrix_5_31_port, C(20) => aMatrix_5_31_port, C(19)
                           => aMatrix_5_31_port, C(18) => aMatrix_5_31_port, 
                           C(17) => aMatrix_5_17_port, C(16) => 
                           aMatrix_5_16_port, C(15) => aMatrix_5_15_port, C(14)
                           => aMatrix_5_14_port, C(13) => aMatrix_5_13_port, 
                           C(12) => aMatrix_5_12_port, C(11) => 
                           aMatrix_5_11_port, C(10) => aMatrix_5_10_port, C(9) 
                           => aMatrix_5_9_port, C(8) => aMatrix_5_8_port, C(7) 
                           => aMatrix_5_7_port, C(6) => aMatrix_5_6_port, C(5) 
                           => aMatrix_5_5_port, C(4) => aMatrix_5_4_port, C(3) 
                           => aMatrix_5_3_port, C(2) => A(0), C(1) => n29, C(0)
                           => aMatrix_5_0_port, D(31) => n18, D(30) => n18, 
                           D(29) => n17, D(28) => n17, D(27) => n17, D(26) => 
                           n17, D(25) => n17, D(24) => n17, D(23) => n17, D(22)
                           => n17, D(21) => n17, D(20) => n17, D(19) => n17, 
                           D(18) => n17, D(17) => A(14), D(16) => A(13), D(15) 
                           => A(12), D(14) => A(11), D(13) => A(10), D(12) => 
                           A(9), D(11) => A(8), D(10) => A(7), D(9) => A(6), 
                           D(8) => A(5), D(7) => A(4), D(6) => A(3), D(5) => 
                           A(2), D(4) => n2, D(3) => A(0), D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => aMatrix_7_31_port, E(30) => 
                           aMatrix_7_31_port, E(29) => aMatrix_7_31_port, E(28)
                           => aMatrix_7_31_port, E(27) => aMatrix_7_31_port, 
                           E(26) => aMatrix_7_31_port, E(25) => 
                           aMatrix_7_31_port, E(24) => aMatrix_7_31_port, E(23)
                           => aMatrix_7_31_port, E(22) => aMatrix_7_31_port, 
                           E(21) => aMatrix_7_31_port, E(20) => 
                           aMatrix_7_31_port, E(19) => aMatrix_7_31_port, E(18)
                           => aMatrix_7_18_port, E(17) => aMatrix_7_17_port, 
                           E(16) => aMatrix_7_16_port, E(15) => 
                           aMatrix_7_15_port, E(14) => aMatrix_7_14_port, E(13)
                           => aMatrix_7_13_port, E(12) => aMatrix_7_12_port, 
                           E(11) => aMatrix_7_11_port, E(10) => 
                           aMatrix_7_10_port, E(9) => aMatrix_7_9_port, E(8) =>
                           aMatrix_7_8_port, E(7) => aMatrix_7_7_port, E(6) => 
                           aMatrix_7_6_port, E(5) => aMatrix_7_5_port, E(4) => 
                           aMatrix_7_4_port, E(3) => A(0), E(2) => n29, E(1) =>
                           n29, E(0) => aMatrix_7_0_port, F(31) => 
                           X_Logic0_port, F(30) => X_Logic0_port, F(29) => 
                           X_Logic0_port, F(28) => X_Logic0_port, F(27) => 
                           X_Logic0_port, F(26) => X_Logic0_port, F(25) => 
                           X_Logic0_port, F(24) => X_Logic0_port, F(23) => 
                           X_Logic0_port, F(22) => X_Logic0_port, F(21) => 
                           X_Logic0_port, F(20) => X_Logic0_port, F(19) => 
                           X_Logic0_port, F(18) => X_Logic0_port, F(17) => 
                           X_Logic0_port, F(16) => X_Logic0_port, F(15) => 
                           X_Logic0_port, F(14) => X_Logic0_port, F(13) => 
                           X_Logic0_port, F(12) => X_Logic0_port, F(11) => 
                           X_Logic0_port, F(10) => X_Logic0_port, F(9) => 
                           X_Logic0_port, F(8) => X_Logic0_port, F(7) => 
                           X_Logic0_port, F(6) => X_Logic0_port, F(5) => 
                           X_Logic0_port, F(4) => X_Logic0_port, F(3) => 
                           X_Logic0_port, F(2) => X_Logic0_port, F(1) => 
                           X_Logic0_port, F(0) => X_Logic0_port, G(31) => 
                           X_Logic0_port, G(30) => X_Logic0_port, G(29) => 
                           X_Logic0_port, G(28) => X_Logic0_port, G(27) => 
                           X_Logic0_port, G(26) => X_Logic0_port, G(25) => 
                           X_Logic0_port, G(24) => X_Logic0_port, G(23) => 
                           X_Logic0_port, G(22) => X_Logic0_port, G(21) => 
                           X_Logic0_port, G(20) => X_Logic0_port, G(19) => 
                           X_Logic0_port, G(18) => X_Logic0_port, G(17) => 
                           X_Logic0_port, G(16) => X_Logic0_port, G(15) => 
                           X_Logic0_port, G(14) => X_Logic0_port, G(13) => 
                           X_Logic0_port, G(12) => X_Logic0_port, G(11) => 
                           X_Logic0_port, G(10) => X_Logic0_port, G(9) => 
                           X_Logic0_port, G(8) => X_Logic0_port, G(7) => 
                           X_Logic0_port, G(6) => X_Logic0_port, G(5) => 
                           X_Logic0_port, G(4) => X_Logic0_port, G(3) => 
                           X_Logic0_port, G(2) => X_Logic0_port, G(1) => 
                           X_Logic0_port, G(0) => X_Logic0_port, H(31) => 
                           X_Logic0_port, H(30) => X_Logic0_port, H(29) => 
                           X_Logic0_port, H(28) => X_Logic0_port, H(27) => 
                           X_Logic0_port, H(26) => X_Logic0_port, H(25) => 
                           X_Logic0_port, H(24) => X_Logic0_port, H(23) => 
                           X_Logic0_port, H(22) => X_Logic0_port, H(21) => 
                           X_Logic0_port, H(20) => X_Logic0_port, H(19) => 
                           X_Logic0_port, H(18) => X_Logic0_port, H(17) => 
                           X_Logic0_port, H(16) => X_Logic0_port, H(15) => 
                           X_Logic0_port, H(14) => X_Logic0_port, H(13) => 
                           X_Logic0_port, H(12) => X_Logic0_port, H(11) => 
                           X_Logic0_port, H(10) => X_Logic0_port, H(9) => 
                           X_Logic0_port, H(8) => X_Logic0_port, H(7) => 
                           X_Logic0_port, H(6) => X_Logic0_port, H(5) => 
                           X_Logic0_port, H(4) => X_Logic0_port, H(3) => 
                           X_Logic0_port, H(2) => X_Logic0_port, H(1) => 
                           X_Logic0_port, H(0) => X_Logic0_port, S(2) => 
                           Bo_signal_5_port, S(1) => Bo_signal_4_port, S(0) => 
                           Bo_signal_3_port, Y(31) => aEncMatrix_1_31_port, 
                           Y(30) => aEncMatrix_1_30_port, Y(29) => 
                           aEncMatrix_1_29_port, Y(28) => aEncMatrix_1_28_port,
                           Y(27) => aEncMatrix_1_27_port, Y(26) => 
                           aEncMatrix_1_26_port, Y(25) => aEncMatrix_1_25_port,
                           Y(24) => aEncMatrix_1_24_port, Y(23) => 
                           aEncMatrix_1_23_port, Y(22) => aEncMatrix_1_22_port,
                           Y(21) => aEncMatrix_1_21_port, Y(20) => 
                           aEncMatrix_1_20_port, Y(19) => aEncMatrix_1_19_port,
                           Y(18) => aEncMatrix_1_18_port, Y(17) => 
                           aEncMatrix_1_17_port, Y(16) => aEncMatrix_1_16_port,
                           Y(15) => aEncMatrix_1_15_port, Y(14) => 
                           aEncMatrix_1_14_port, Y(13) => aEncMatrix_1_13_port,
                           Y(12) => aEncMatrix_1_12_port, Y(11) => 
                           aEncMatrix_1_11_port, Y(10) => aEncMatrix_1_10_port,
                           Y(9) => aEncMatrix_1_9_port, Y(8) => 
                           aEncMatrix_1_8_port, Y(7) => aEncMatrix_1_7_port, 
                           Y(6) => aEncMatrix_1_6_port, Y(5) => 
                           aEncMatrix_1_5_port, Y(4) => aEncMatrix_1_4_port, 
                           Y(3) => aEncMatrix_1_3_port, Y(2) => 
                           aEncMatrix_1_2_port, Y(1) => aEncMatrix_1_1_port, 
                           Y(0) => aEncMatrix_1_0_port);
   FIRST_RCA_1 : RCA_N32_2 port map( A(31) => aEncMatrix_1_31_port, A(30) => 
                           aEncMatrix_1_30_port, A(29) => aEncMatrix_1_29_port,
                           A(28) => aEncMatrix_1_28_port, A(27) => 
                           aEncMatrix_1_27_port, A(26) => aEncMatrix_1_26_port,
                           A(25) => aEncMatrix_1_25_port, A(24) => 
                           aEncMatrix_1_24_port, A(23) => aEncMatrix_1_23_port,
                           A(22) => aEncMatrix_1_22_port, A(21) => 
                           aEncMatrix_1_21_port, A(20) => aEncMatrix_1_20_port,
                           A(19) => aEncMatrix_1_19_port, A(18) => 
                           aEncMatrix_1_18_port, A(17) => aEncMatrix_1_17_port,
                           A(16) => aEncMatrix_1_16_port, A(15) => 
                           aEncMatrix_1_15_port, A(14) => aEncMatrix_1_14_port,
                           A(13) => aEncMatrix_1_13_port, A(12) => 
                           aEncMatrix_1_12_port, A(11) => aEncMatrix_1_11_port,
                           A(10) => aEncMatrix_1_10_port, A(9) => 
                           aEncMatrix_1_9_port, A(8) => aEncMatrix_1_8_port, 
                           A(7) => aEncMatrix_1_7_port, A(6) => 
                           aEncMatrix_1_6_port, A(5) => aEncMatrix_1_5_port, 
                           A(4) => aEncMatrix_1_4_port, A(3) => 
                           aEncMatrix_1_3_port, A(2) => aEncMatrix_1_2_port, 
                           A(1) => aEncMatrix_1_1_port, A(0) => 
                           aEncMatrix_1_0_port, B(31) => aEncMatrix_0_31_port, 
                           B(30) => aEncMatrix_0_30_port, B(29) => 
                           aEncMatrix_0_29_port, B(28) => aEncMatrix_0_28_port,
                           B(27) => aEncMatrix_0_27_port, B(26) => 
                           aEncMatrix_0_26_port, B(25) => aEncMatrix_0_25_port,
                           B(24) => aEncMatrix_0_24_port, B(23) => 
                           aEncMatrix_0_23_port, B(22) => aEncMatrix_0_22_port,
                           B(21) => aEncMatrix_0_21_port, B(20) => 
                           aEncMatrix_0_20_port, B(19) => aEncMatrix_0_19_port,
                           B(18) => aEncMatrix_0_18_port, B(17) => 
                           aEncMatrix_0_17_port, B(16) => aEncMatrix_0_16_port,
                           B(15) => aEncMatrix_0_15_port, B(14) => 
                           aEncMatrix_0_14_port, B(13) => aEncMatrix_0_13_port,
                           B(12) => aEncMatrix_0_12_port, B(11) => 
                           aEncMatrix_0_11_port, B(10) => aEncMatrix_0_10_port,
                           B(9) => aEncMatrix_0_9_port, B(8) => 
                           aEncMatrix_0_8_port, B(7) => aEncMatrix_0_7_port, 
                           B(6) => aEncMatrix_0_6_port, B(5) => 
                           aEncMatrix_0_5_port, B(4) => aEncMatrix_0_4_port, 
                           B(3) => aEncMatrix_0_3_port, B(2) => 
                           aEncMatrix_0_2_port, B(1) => aEncMatrix_0_1_port, 
                           B(0) => aEncMatrix_0_0_port, Ci => X_Logic0_port, 
                           S(31) => pSumMatrix_0_31_port, S(30) => 
                           pSumMatrix_0_30_port, S(29) => pSumMatrix_0_29_port,
                           S(28) => pSumMatrix_0_28_port, S(27) => 
                           pSumMatrix_0_27_port, S(26) => pSumMatrix_0_26_port,
                           S(25) => pSumMatrix_0_25_port, S(24) => 
                           pSumMatrix_0_24_port, S(23) => pSumMatrix_0_23_port,
                           S(22) => pSumMatrix_0_22_port, S(21) => 
                           pSumMatrix_0_21_port, S(20) => pSumMatrix_0_20_port,
                           S(19) => pSumMatrix_0_19_port, S(18) => 
                           pSumMatrix_0_18_port, S(17) => pSumMatrix_0_17_port,
                           S(16) => pSumMatrix_0_16_port, S(15) => 
                           pSumMatrix_0_15_port, S(14) => pSumMatrix_0_14_port,
                           S(13) => pSumMatrix_0_13_port, S(12) => 
                           pSumMatrix_0_12_port, S(11) => pSumMatrix_0_11_port,
                           S(10) => pSumMatrix_0_10_port, S(9) => 
                           pSumMatrix_0_9_port, S(8) => pSumMatrix_0_8_port, 
                           S(7) => pSumMatrix_0_7_port, S(6) => 
                           pSumMatrix_0_6_port, S(5) => pSumMatrix_0_5_port, 
                           S(4) => pSumMatrix_0_4_port, S(3) => 
                           pSumMatrix_0_3_port, S(2) => pSumMatrix_0_2_port, 
                           S(1) => pSumMatrix_0_1_port, S(0) => 
                           pSumMatrix_0_0_port, Co => n_1270);
   MUXES_2 : MUX81_N32_1 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => n21, B(30) => n20, B(29) => 
                           n18, B(28) => A(15), B(27) => n17, B(26) => n19, 
                           B(25) => n21, B(24) => n20, B(23) => A(15), B(22) =>
                           n17, B(21) => n19, B(20) => n18, B(19) => n21, B(18)
                           => A(14), B(17) => A(13), B(16) => A(12), B(15) => 
                           A(11), B(14) => A(10), B(13) => A(9), B(12) => A(8),
                           B(11) => A(7), B(10) => A(6), B(9) => A(5), B(8) => 
                           A(4), B(7) => A(3), B(6) => A(2), B(5) => n2, B(4) 
                           => A(0), B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, C(31) => aMatrix_9_31_port, C(30) => 
                           aMatrix_9_31_port, C(29) => aMatrix_9_31_port, C(28)
                           => aMatrix_9_31_port, C(27) => aMatrix_9_31_port, 
                           C(26) => aMatrix_9_31_port, C(25) => 
                           aMatrix_9_31_port, C(24) => aMatrix_9_31_port, C(23)
                           => aMatrix_9_31_port, C(22) => aMatrix_9_31_port, 
                           C(21) => aMatrix_9_31_port, C(20) => 
                           aMatrix_9_31_port, C(19) => aMatrix_9_19_port, C(18)
                           => aMatrix_9_18_port, C(17) => aMatrix_9_17_port, 
                           C(16) => aMatrix_9_16_port, C(15) => 
                           aMatrix_9_15_port, C(14) => aMatrix_9_14_port, C(13)
                           => aMatrix_9_13_port, C(12) => aMatrix_9_12_port, 
                           C(11) => aMatrix_9_11_port, C(10) => 
                           aMatrix_9_10_port, C(9) => aMatrix_9_9_port, C(8) =>
                           aMatrix_9_8_port, C(7) => aMatrix_9_7_port, C(6) => 
                           aMatrix_9_6_port, C(5) => aMatrix_9_5_port, C(4) => 
                           A(0), C(3) => n29, C(2) => n29, C(1) => n29, C(0) =>
                           aMatrix_9_0_port, D(31) => n20, D(30) => n18, D(29) 
                           => A(15), D(28) => n17, D(27) => n19, D(26) => n19, 
                           D(25) => n19, D(24) => n19, D(23) => n19, D(22) => 
                           n19, D(21) => n19, D(20) => n19, D(19) => A(14), 
                           D(18) => A(13), D(17) => A(12), D(16) => A(11), 
                           D(15) => A(10), D(14) => A(9), D(13) => A(8), D(12) 
                           => A(7), D(11) => A(6), D(10) => A(5), D(9) => A(4),
                           D(8) => A(3), D(7) => A(2), D(6) => n2, D(5) => A(0)
                           , D(4) => X_Logic0_port, D(3) => X_Logic0_port, D(2)
                           => X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => aMatrix_11_31_port, E(30) =>
                           aMatrix_11_31_port, E(29) => aMatrix_11_31_port, 
                           E(28) => aMatrix_11_31_port, E(27) => 
                           aMatrix_11_31_port, E(26) => aMatrix_11_31_port, 
                           E(25) => aMatrix_11_31_port, E(24) => 
                           aMatrix_11_31_port, E(23) => aMatrix_11_31_port, 
                           E(22) => aMatrix_11_31_port, E(21) => 
                           aMatrix_11_31_port, E(20) => aMatrix_11_20_port, 
                           E(19) => aMatrix_11_19_port, E(18) => 
                           aMatrix_11_18_port, E(17) => aMatrix_11_17_port, 
                           E(16) => aMatrix_11_16_port, E(15) => 
                           aMatrix_11_15_port, E(14) => aMatrix_11_14_port, 
                           E(13) => aMatrix_11_13_port, E(12) => 
                           aMatrix_11_12_port, E(11) => aMatrix_11_11_port, 
                           E(10) => aMatrix_11_10_port, E(9) => 
                           aMatrix_11_9_port, E(8) => aMatrix_11_8_port, E(7) 
                           => aMatrix_11_7_port, E(6) => aMatrix_11_6_port, 
                           E(5) => A(0), E(4) => n29, E(3) => n29, E(2) => n29,
                           E(1) => n29, E(0) => aMatrix_11_0_port, F(31) => 
                           X_Logic0_port, F(30) => X_Logic0_port, F(29) => 
                           X_Logic0_port, F(28) => X_Logic0_port, F(27) => 
                           X_Logic0_port, F(26) => X_Logic0_port, F(25) => 
                           X_Logic0_port, F(24) => X_Logic0_port, F(23) => 
                           X_Logic0_port, F(22) => X_Logic0_port, F(21) => 
                           X_Logic0_port, F(20) => X_Logic0_port, F(19) => 
                           X_Logic0_port, F(18) => X_Logic0_port, F(17) => 
                           X_Logic0_port, F(16) => X_Logic0_port, F(15) => 
                           X_Logic0_port, F(14) => X_Logic0_port, F(13) => 
                           X_Logic0_port, F(12) => X_Logic0_port, F(11) => 
                           X_Logic0_port, F(10) => X_Logic0_port, F(9) => 
                           X_Logic0_port, F(8) => X_Logic0_port, F(7) => 
                           X_Logic0_port, F(6) => X_Logic0_port, F(5) => 
                           X_Logic0_port, F(4) => X_Logic0_port, F(3) => 
                           X_Logic0_port, F(2) => X_Logic0_port, F(1) => 
                           X_Logic0_port, F(0) => X_Logic0_port, G(31) => 
                           X_Logic0_port, G(30) => X_Logic0_port, G(29) => 
                           X_Logic0_port, G(28) => X_Logic0_port, G(27) => 
                           X_Logic0_port, G(26) => X_Logic0_port, G(25) => 
                           X_Logic0_port, G(24) => X_Logic0_port, G(23) => 
                           X_Logic0_port, G(22) => X_Logic0_port, G(21) => 
                           X_Logic0_port, G(20) => X_Logic0_port, G(19) => 
                           X_Logic0_port, G(18) => X_Logic0_port, G(17) => 
                           X_Logic0_port, G(16) => X_Logic0_port, G(15) => 
                           X_Logic0_port, G(14) => X_Logic0_port, G(13) => 
                           X_Logic0_port, G(12) => X_Logic0_port, G(11) => 
                           X_Logic0_port, G(10) => X_Logic0_port, G(9) => 
                           X_Logic0_port, G(8) => X_Logic0_port, G(7) => 
                           X_Logic0_port, G(6) => X_Logic0_port, G(5) => 
                           X_Logic0_port, G(4) => X_Logic0_port, G(3) => 
                           X_Logic0_port, G(2) => X_Logic0_port, G(1) => 
                           X_Logic0_port, G(0) => X_Logic0_port, H(31) => 
                           X_Logic0_port, H(30) => X_Logic0_port, H(29) => 
                           X_Logic0_port, H(28) => X_Logic0_port, H(27) => 
                           X_Logic0_port, H(26) => X_Logic0_port, H(25) => 
                           X_Logic0_port, H(24) => X_Logic0_port, H(23) => 
                           X_Logic0_port, H(22) => X_Logic0_port, H(21) => 
                           X_Logic0_port, H(20) => X_Logic0_port, H(19) => 
                           X_Logic0_port, H(18) => X_Logic0_port, H(17) => 
                           X_Logic0_port, H(16) => X_Logic0_port, H(15) => 
                           X_Logic0_port, H(14) => X_Logic0_port, H(13) => 
                           X_Logic0_port, H(12) => X_Logic0_port, H(11) => 
                           X_Logic0_port, H(10) => X_Logic0_port, H(9) => 
                           X_Logic0_port, H(8) => X_Logic0_port, H(7) => 
                           X_Logic0_port, H(6) => X_Logic0_port, H(5) => 
                           X_Logic0_port, H(4) => X_Logic0_port, H(3) => 
                           X_Logic0_port, H(2) => X_Logic0_port, H(1) => 
                           X_Logic0_port, H(0) => X_Logic0_port, S(2) => 
                           Bo_signal_8_port, S(1) => Bo_signal_7_port, S(0) => 
                           Bo_signal_6_port, Y(31) => aEncMatrix_2_31_port, 
                           Y(30) => aEncMatrix_2_30_port, Y(29) => 
                           aEncMatrix_2_29_port, Y(28) => aEncMatrix_2_28_port,
                           Y(27) => aEncMatrix_2_27_port, Y(26) => 
                           aEncMatrix_2_26_port, Y(25) => aEncMatrix_2_25_port,
                           Y(24) => aEncMatrix_2_24_port, Y(23) => 
                           aEncMatrix_2_23_port, Y(22) => aEncMatrix_2_22_port,
                           Y(21) => aEncMatrix_2_21_port, Y(20) => 
                           aEncMatrix_2_20_port, Y(19) => aEncMatrix_2_19_port,
                           Y(18) => aEncMatrix_2_18_port, Y(17) => 
                           aEncMatrix_2_17_port, Y(16) => aEncMatrix_2_16_port,
                           Y(15) => aEncMatrix_2_15_port, Y(14) => 
                           aEncMatrix_2_14_port, Y(13) => aEncMatrix_2_13_port,
                           Y(12) => aEncMatrix_2_12_port, Y(11) => 
                           aEncMatrix_2_11_port, Y(10) => aEncMatrix_2_10_port,
                           Y(9) => aEncMatrix_2_9_port, Y(8) => 
                           aEncMatrix_2_8_port, Y(7) => aEncMatrix_2_7_port, 
                           Y(6) => aEncMatrix_2_6_port, Y(5) => 
                           aEncMatrix_2_5_port, Y(4) => aEncMatrix_2_4_port, 
                           Y(3) => aEncMatrix_2_3_port, Y(2) => 
                           aEncMatrix_2_2_port, Y(1) => aEncMatrix_2_1_port, 
                           Y(0) => aEncMatrix_2_0_port);
   RCAS_2 : RCA_N32_1 port map( A(31) => aEncMatrix_2_31_port, A(30) => 
                           aEncMatrix_2_30_port, A(29) => aEncMatrix_2_29_port,
                           A(28) => aEncMatrix_2_28_port, A(27) => 
                           aEncMatrix_2_27_port, A(26) => aEncMatrix_2_26_port,
                           A(25) => aEncMatrix_2_25_port, A(24) => 
                           aEncMatrix_2_24_port, A(23) => aEncMatrix_2_23_port,
                           A(22) => aEncMatrix_2_22_port, A(21) => 
                           aEncMatrix_2_21_port, A(20) => aEncMatrix_2_20_port,
                           A(19) => aEncMatrix_2_19_port, A(18) => 
                           aEncMatrix_2_18_port, A(17) => aEncMatrix_2_17_port,
                           A(16) => aEncMatrix_2_16_port, A(15) => 
                           aEncMatrix_2_15_port, A(14) => aEncMatrix_2_14_port,
                           A(13) => aEncMatrix_2_13_port, A(12) => 
                           aEncMatrix_2_12_port, A(11) => aEncMatrix_2_11_port,
                           A(10) => aEncMatrix_2_10_port, A(9) => 
                           aEncMatrix_2_9_port, A(8) => aEncMatrix_2_8_port, 
                           A(7) => aEncMatrix_2_7_port, A(6) => 
                           aEncMatrix_2_6_port, A(5) => aEncMatrix_2_5_port, 
                           A(4) => aEncMatrix_2_4_port, A(3) => 
                           aEncMatrix_2_3_port, A(2) => aEncMatrix_2_2_port, 
                           A(1) => aEncMatrix_2_1_port, A(0) => 
                           aEncMatrix_2_0_port, B(31) => pSumMatrix_0_31_port, 
                           B(30) => pSumMatrix_0_30_port, B(29) => 
                           pSumMatrix_0_29_port, B(28) => pSumMatrix_0_28_port,
                           B(27) => pSumMatrix_0_27_port, B(26) => 
                           pSumMatrix_0_26_port, B(25) => pSumMatrix_0_25_port,
                           B(24) => pSumMatrix_0_24_port, B(23) => 
                           pSumMatrix_0_23_port, B(22) => pSumMatrix_0_22_port,
                           B(21) => pSumMatrix_0_21_port, B(20) => 
                           pSumMatrix_0_20_port, B(19) => pSumMatrix_0_19_port,
                           B(18) => pSumMatrix_0_18_port, B(17) => 
                           pSumMatrix_0_17_port, B(16) => pSumMatrix_0_16_port,
                           B(15) => pSumMatrix_0_15_port, B(14) => 
                           pSumMatrix_0_14_port, B(13) => pSumMatrix_0_13_port,
                           B(12) => pSumMatrix_0_12_port, B(11) => 
                           pSumMatrix_0_11_port, B(10) => pSumMatrix_0_10_port,
                           B(9) => pSumMatrix_0_9_port, B(8) => 
                           pSumMatrix_0_8_port, B(7) => pSumMatrix_0_7_port, 
                           B(6) => pSumMatrix_0_6_port, B(5) => 
                           pSumMatrix_0_5_port, B(4) => pSumMatrix_0_4_port, 
                           B(3) => pSumMatrix_0_3_port, B(2) => 
                           pSumMatrix_0_2_port, B(1) => pSumMatrix_0_1_port, 
                           B(0) => pSumMatrix_0_0_port, Ci => X_Logic0_port, 
                           S(31) => pSumMatrix_1_31_port, S(30) => 
                           pSumMatrix_1_30_port, S(29) => pSumMatrix_1_29_port,
                           S(28) => pSumMatrix_1_28_port, S(27) => 
                           pSumMatrix_1_27_port, S(26) => pSumMatrix_1_26_port,
                           S(25) => pSumMatrix_1_25_port, S(24) => 
                           pSumMatrix_1_24_port, S(23) => pSumMatrix_1_23_port,
                           S(22) => pSumMatrix_1_22_port, S(21) => 
                           pSumMatrix_1_21_port, S(20) => pSumMatrix_1_20_port,
                           S(19) => pSumMatrix_1_19_port, S(18) => 
                           pSumMatrix_1_18_port, S(17) => pSumMatrix_1_17_port,
                           S(16) => pSumMatrix_1_16_port, S(15) => 
                           pSumMatrix_1_15_port, S(14) => pSumMatrix_1_14_port,
                           S(13) => pSumMatrix_1_13_port, S(12) => 
                           pSumMatrix_1_12_port, S(11) => pSumMatrix_1_11_port,
                           S(10) => pSumMatrix_1_10_port, S(9) => 
                           pSumMatrix_1_9_port, S(8) => pSumMatrix_1_8_port, 
                           S(7) => pSumMatrix_1_7_port, S(6) => 
                           pSumMatrix_1_6_port, S(5) => pSumMatrix_1_5_port, 
                           S(4) => pSumMatrix_1_4_port, S(3) => 
                           pSumMatrix_1_3_port, S(2) => pSumMatrix_1_2_port, 
                           S(1) => pSumMatrix_1_1_port, S(0) => 
                           pSumMatrix_1_0_port, Co => n_1271);
   MUXES_3 : MUX81_N32_0 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => n20, B(30) => n20, B(29) => 
                           n20, B(28) => n21, B(27) => n20, B(26) => A(15), 
                           B(25) => n17, B(24) => n19, B(23) => n18, B(22) => 
                           n19, B(21) => n17, B(20) => A(14), B(19) => A(13), 
                           B(18) => A(12), B(17) => A(11), B(16) => A(10), 
                           B(15) => A(9), B(14) => A(8), B(13) => A(7), B(12) 
                           => A(6), B(11) => A(5), B(10) => A(4), B(9) => A(3),
                           B(8) => A(2), B(7) => n2, B(6) => A(0), B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => 
                           aMatrix_13_31_port, C(30) => aMatrix_13_31_port, 
                           C(29) => aMatrix_13_31_port, C(28) => 
                           aMatrix_13_31_port, C(27) => aMatrix_13_31_port, 
                           C(26) => aMatrix_13_31_port, C(25) => 
                           aMatrix_13_31_port, C(24) => aMatrix_13_31_port, 
                           C(23) => aMatrix_13_31_port, C(22) => 
                           aMatrix_13_31_port, C(21) => aMatrix_13_21_port, 
                           C(20) => aMatrix_13_20_port, C(19) => 
                           aMatrix_13_19_port, C(18) => aMatrix_13_18_port, 
                           C(17) => aMatrix_13_17_port, C(16) => 
                           aMatrix_13_16_port, C(15) => aMatrix_13_15_port, 
                           C(14) => aMatrix_13_14_port, C(13) => 
                           aMatrix_13_13_port, C(12) => aMatrix_13_12_port, 
                           C(11) => aMatrix_13_11_port, C(10) => 
                           aMatrix_13_10_port, C(9) => aMatrix_13_9_port, C(8) 
                           => aMatrix_13_8_port, C(7) => aMatrix_13_7_port, 
                           C(6) => A(0), C(5) => n29, C(4) => n29, C(3) => n29,
                           C(2) => n29, C(1) => n29, C(0) => aMatrix_13_0_port,
                           D(31) => n21, D(30) => n20, D(29) => A(15), D(28) =>
                           n17, D(27) => n21, D(26) => n20, D(25) => n18, D(24)
                           => A(15), D(23) => n17, D(22) => n19, D(21) => A(14)
                           , D(20) => A(13), D(19) => A(12), D(18) => A(11), 
                           D(17) => A(10), D(16) => A(9), D(15) => A(8), D(14) 
                           => A(7), D(13) => A(6), D(12) => A(5), D(11) => A(4)
                           , D(10) => A(3), D(9) => A(2), D(8) => n2, D(7) => 
                           A(0), D(6) => X_Logic0_port, D(5) => X_Logic0_port, 
                           D(4) => X_Logic0_port, D(3) => X_Logic0_port, D(2) 
                           => X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(31) => aMatrix_15_31_port, E(30) =>
                           aMatrix_15_31_port, E(29) => aMatrix_15_31_port, 
                           E(28) => aMatrix_15_31_port, E(27) => 
                           aMatrix_15_31_port, E(26) => aMatrix_15_31_port, 
                           E(25) => aMatrix_15_31_port, E(24) => 
                           aMatrix_15_31_port, E(23) => aMatrix_15_31_port, 
                           E(22) => aMatrix_15_22_port, E(21) => 
                           aMatrix_15_21_port, E(20) => aMatrix_15_20_port, 
                           E(19) => aMatrix_15_19_port, E(18) => 
                           aMatrix_15_18_port, E(17) => aMatrix_15_17_port, 
                           E(16) => aMatrix_15_16_port, E(15) => 
                           aMatrix_15_15_port, E(14) => aMatrix_15_14_port, 
                           E(13) => aMatrix_15_13_port, E(12) => 
                           aMatrix_15_12_port, E(11) => aMatrix_15_11_port, 
                           E(10) => aMatrix_15_10_port, E(9) => 
                           aMatrix_15_9_port, E(8) => aMatrix_15_8_port, E(7) 
                           => A(0), E(6) => n29, E(5) => n29, E(4) => n29, E(3)
                           => n29, E(2) => n29, E(1) => n29, E(0) => 
                           aMatrix_15_0_port, F(31) => X_Logic0_port, F(30) => 
                           X_Logic0_port, F(29) => X_Logic0_port, F(28) => 
                           X_Logic0_port, F(27) => X_Logic0_port, F(26) => 
                           X_Logic0_port, F(25) => X_Logic0_port, F(24) => 
                           X_Logic0_port, F(23) => X_Logic0_port, F(22) => 
                           X_Logic0_port, F(21) => X_Logic0_port, F(20) => 
                           X_Logic0_port, F(19) => X_Logic0_port, F(18) => 
                           X_Logic0_port, F(17) => X_Logic0_port, F(16) => 
                           X_Logic0_port, F(15) => X_Logic0_port, F(14) => 
                           X_Logic0_port, F(13) => X_Logic0_port, F(12) => 
                           X_Logic0_port, F(11) => X_Logic0_port, F(10) => 
                           X_Logic0_port, F(9) => X_Logic0_port, F(8) => 
                           X_Logic0_port, F(7) => X_Logic0_port, F(6) => 
                           X_Logic0_port, F(5) => X_Logic0_port, F(4) => 
                           X_Logic0_port, F(3) => X_Logic0_port, F(2) => 
                           X_Logic0_port, F(1) => X_Logic0_port, F(0) => 
                           X_Logic0_port, G(31) => X_Logic0_port, G(30) => 
                           X_Logic0_port, G(29) => X_Logic0_port, G(28) => 
                           X_Logic0_port, G(27) => X_Logic0_port, G(26) => 
                           X_Logic0_port, G(25) => X_Logic0_port, G(24) => 
                           X_Logic0_port, G(23) => X_Logic0_port, G(22) => 
                           X_Logic0_port, G(21) => X_Logic0_port, G(20) => 
                           X_Logic0_port, G(19) => X_Logic0_port, G(18) => 
                           X_Logic0_port, G(17) => X_Logic0_port, G(16) => 
                           X_Logic0_port, G(15) => X_Logic0_port, G(14) => 
                           X_Logic0_port, G(13) => X_Logic0_port, G(12) => 
                           X_Logic0_port, G(11) => X_Logic0_port, G(10) => 
                           X_Logic0_port, G(9) => X_Logic0_port, G(8) => 
                           X_Logic0_port, G(7) => X_Logic0_port, G(6) => 
                           X_Logic0_port, G(5) => X_Logic0_port, G(4) => 
                           X_Logic0_port, G(3) => X_Logic0_port, G(2) => 
                           X_Logic0_port, G(1) => X_Logic0_port, G(0) => 
                           X_Logic0_port, H(31) => X_Logic0_port, H(30) => 
                           X_Logic0_port, H(29) => X_Logic0_port, H(28) => 
                           X_Logic0_port, H(27) => X_Logic0_port, H(26) => 
                           X_Logic0_port, H(25) => X_Logic0_port, H(24) => 
                           X_Logic0_port, H(23) => X_Logic0_port, H(22) => 
                           X_Logic0_port, H(21) => X_Logic0_port, H(20) => 
                           X_Logic0_port, H(19) => X_Logic0_port, H(18) => 
                           X_Logic0_port, H(17) => X_Logic0_port, H(16) => 
                           X_Logic0_port, H(15) => X_Logic0_port, H(14) => 
                           X_Logic0_port, H(13) => X_Logic0_port, H(12) => 
                           X_Logic0_port, H(11) => X_Logic0_port, H(10) => 
                           X_Logic0_port, H(9) => X_Logic0_port, H(8) => 
                           X_Logic0_port, H(7) => X_Logic0_port, H(6) => 
                           X_Logic0_port, H(5) => X_Logic0_port, H(4) => 
                           X_Logic0_port, H(3) => X_Logic0_port, H(2) => 
                           X_Logic0_port, H(1) => X_Logic0_port, H(0) => 
                           X_Logic0_port, S(2) => Bo_signal_11_port, S(1) => 
                           Bo_signal_10_port, S(0) => Bo_signal_9_port, Y(31) 
                           => aEncMatrix_3_31_port, Y(30) => 
                           aEncMatrix_3_30_port, Y(29) => aEncMatrix_3_29_port,
                           Y(28) => aEncMatrix_3_28_port, Y(27) => 
                           aEncMatrix_3_27_port, Y(26) => aEncMatrix_3_26_port,
                           Y(25) => aEncMatrix_3_25_port, Y(24) => 
                           aEncMatrix_3_24_port, Y(23) => aEncMatrix_3_23_port,
                           Y(22) => aEncMatrix_3_22_port, Y(21) => 
                           aEncMatrix_3_21_port, Y(20) => aEncMatrix_3_20_port,
                           Y(19) => aEncMatrix_3_19_port, Y(18) => 
                           aEncMatrix_3_18_port, Y(17) => aEncMatrix_3_17_port,
                           Y(16) => aEncMatrix_3_16_port, Y(15) => 
                           aEncMatrix_3_15_port, Y(14) => aEncMatrix_3_14_port,
                           Y(13) => aEncMatrix_3_13_port, Y(12) => 
                           aEncMatrix_3_12_port, Y(11) => aEncMatrix_3_11_port,
                           Y(10) => aEncMatrix_3_10_port, Y(9) => 
                           aEncMatrix_3_9_port, Y(8) => aEncMatrix_3_8_port, 
                           Y(7) => aEncMatrix_3_7_port, Y(6) => 
                           aEncMatrix_3_6_port, Y(5) => aEncMatrix_3_5_port, 
                           Y(4) => aEncMatrix_3_4_port, Y(3) => 
                           aEncMatrix_3_3_port, Y(2) => aEncMatrix_3_2_port, 
                           Y(1) => aEncMatrix_3_1_port, Y(0) => 
                           aEncMatrix_3_0_port);
   RCAS_3 : RCA_N32_0 port map( A(31) => aEncMatrix_3_31_port, A(30) => 
                           aEncMatrix_3_30_port, A(29) => aEncMatrix_3_29_port,
                           A(28) => aEncMatrix_3_28_port, A(27) => 
                           aEncMatrix_3_27_port, A(26) => aEncMatrix_3_26_port,
                           A(25) => aEncMatrix_3_25_port, A(24) => 
                           aEncMatrix_3_24_port, A(23) => aEncMatrix_3_23_port,
                           A(22) => aEncMatrix_3_22_port, A(21) => 
                           aEncMatrix_3_21_port, A(20) => aEncMatrix_3_20_port,
                           A(19) => aEncMatrix_3_19_port, A(18) => 
                           aEncMatrix_3_18_port, A(17) => aEncMatrix_3_17_port,
                           A(16) => aEncMatrix_3_16_port, A(15) => 
                           aEncMatrix_3_15_port, A(14) => aEncMatrix_3_14_port,
                           A(13) => aEncMatrix_3_13_port, A(12) => 
                           aEncMatrix_3_12_port, A(11) => aEncMatrix_3_11_port,
                           A(10) => aEncMatrix_3_10_port, A(9) => 
                           aEncMatrix_3_9_port, A(8) => aEncMatrix_3_8_port, 
                           A(7) => aEncMatrix_3_7_port, A(6) => 
                           aEncMatrix_3_6_port, A(5) => aEncMatrix_3_5_port, 
                           A(4) => aEncMatrix_3_4_port, A(3) => 
                           aEncMatrix_3_3_port, A(2) => aEncMatrix_3_2_port, 
                           A(1) => aEncMatrix_3_1_port, A(0) => 
                           aEncMatrix_3_0_port, B(31) => pSumMatrix_1_31_port, 
                           B(30) => pSumMatrix_1_30_port, B(29) => 
                           pSumMatrix_1_29_port, B(28) => pSumMatrix_1_28_port,
                           B(27) => pSumMatrix_1_27_port, B(26) => 
                           pSumMatrix_1_26_port, B(25) => pSumMatrix_1_25_port,
                           B(24) => pSumMatrix_1_24_port, B(23) => 
                           pSumMatrix_1_23_port, B(22) => pSumMatrix_1_22_port,
                           B(21) => pSumMatrix_1_21_port, B(20) => 
                           pSumMatrix_1_20_port, B(19) => pSumMatrix_1_19_port,
                           B(18) => pSumMatrix_1_18_port, B(17) => 
                           pSumMatrix_1_17_port, B(16) => pSumMatrix_1_16_port,
                           B(15) => pSumMatrix_1_15_port, B(14) => 
                           pSumMatrix_1_14_port, B(13) => pSumMatrix_1_13_port,
                           B(12) => pSumMatrix_1_12_port, B(11) => 
                           pSumMatrix_1_11_port, B(10) => pSumMatrix_1_10_port,
                           B(9) => pSumMatrix_1_9_port, B(8) => 
                           pSumMatrix_1_8_port, B(7) => pSumMatrix_1_7_port, 
                           B(6) => pSumMatrix_1_6_port, B(5) => 
                           pSumMatrix_1_5_port, B(4) => pSumMatrix_1_4_port, 
                           B(3) => pSumMatrix_1_3_port, B(2) => 
                           pSumMatrix_1_2_port, B(1) => pSumMatrix_1_1_port, 
                           B(0) => pSumMatrix_1_0_port, Ci => X_Logic0_port, 
                           S(31) => P(31), S(30) => P(30), S(29) => P(29), 
                           S(28) => P(28), S(27) => P(27), S(26) => P(26), 
                           S(25) => P(25), S(24) => P(24), S(23) => P(23), 
                           S(22) => P(22), S(21) => P(21), S(20) => P(20), 
                           S(19) => P(19), S(18) => P(18), S(17) => P(17), 
                           S(16) => P(16), S(15) => P(15), S(14) => P(14), 
                           S(13) => P(13), S(12) => P(12), S(11) => P(11), 
                           S(10) => P(10), S(9) => P(9), S(8) => P(8), S(7) => 
                           P(7), S(6) => P(6), S(5) => P(5), S(4) => P(4), S(3)
                           => P(3), S(2) => P(2), S(1) => P(1), S(0) => P(0), 
                           Co => n_1272);
   add_92_G8_U1_1_8 : HA_X1 port map( A => n3, B => n1, CO => 
                           add_92_G8_carry_9_port, S => aMatrix_15_8_port);
   add_92_G8_U1_1_9 : HA_X1 port map( A => n4, B => add_92_G8_carry_9_port, CO 
                           => add_92_G8_carry_10_port, S => aMatrix_15_9_port);
   add_92_G8_U1_1_10 : HA_X1 port map( A => n5, B => add_92_G8_carry_10_port, 
                           CO => add_92_G8_carry_11_port, S => 
                           aMatrix_15_10_port);
   add_92_G8_U1_1_11 : HA_X1 port map( A => n6, B => add_92_G8_carry_11_port, 
                           CO => add_92_G8_carry_12_port, S => 
                           aMatrix_15_11_port);
   add_92_G8_U1_1_12 : HA_X1 port map( A => n7, B => add_92_G8_carry_12_port, 
                           CO => add_92_G8_carry_13_port, S => 
                           aMatrix_15_12_port);
   add_92_G8_U1_1_13 : HA_X1 port map( A => n8, B => add_92_G8_carry_13_port, 
                           CO => add_92_G8_carry_14_port, S => 
                           aMatrix_15_13_port);
   add_92_G8_U1_1_14 : HA_X1 port map( A => n9, B => add_92_G8_carry_14_port, 
                           CO => add_92_G8_carry_15_port, S => 
                           aMatrix_15_14_port);
   add_92_G8_U1_1_15 : HA_X1 port map( A => n10, B => add_92_G8_carry_15_port, 
                           CO => add_92_G8_carry_16_port, S => 
                           aMatrix_15_15_port);
   add_92_G8_U1_1_16 : HA_X1 port map( A => n11, B => add_92_G8_carry_16_port, 
                           CO => add_92_G8_carry_17_port, S => 
                           aMatrix_15_16_port);
   add_92_G8_U1_1_17 : HA_X1 port map( A => n12, B => add_92_G8_carry_17_port, 
                           CO => add_92_G8_carry_18_port, S => 
                           aMatrix_15_17_port);
   add_92_G8_U1_1_18 : HA_X1 port map( A => n13, B => add_92_G8_carry_18_port, 
                           CO => add_92_G8_carry_19_port, S => 
                           aMatrix_15_18_port);
   add_92_G8_U1_1_19 : HA_X1 port map( A => n14, B => add_92_G8_carry_19_port, 
                           CO => add_92_G8_carry_20_port, S => 
                           aMatrix_15_19_port);
   add_92_G8_U1_1_20 : HA_X1 port map( A => n15, B => add_92_G8_carry_20_port, 
                           CO => add_92_G8_carry_21_port, S => 
                           aMatrix_15_20_port);
   add_92_G8_U1_1_21 : HA_X1 port map( A => n16, B => add_92_G8_carry_21_port, 
                           CO => add_92_G8_carry_22_port, S => 
                           aMatrix_15_21_port);
   add_92_G7_U1_1_7 : HA_X1 port map( A => n3, B => n1, CO => 
                           add_92_G7_carry_8_port, S => aMatrix_13_7_port);
   add_92_G7_U1_1_8 : HA_X1 port map( A => n4, B => add_92_G7_carry_8_port, CO 
                           => add_92_G7_carry_9_port, S => aMatrix_13_8_port);
   add_92_G7_U1_1_9 : HA_X1 port map( A => n5, B => add_92_G7_carry_9_port, CO 
                           => add_92_G7_carry_10_port, S => aMatrix_13_9_port);
   add_92_G7_U1_1_10 : HA_X1 port map( A => n6, B => add_92_G7_carry_10_port, 
                           CO => add_92_G7_carry_11_port, S => 
                           aMatrix_13_10_port);
   add_92_G7_U1_1_11 : HA_X1 port map( A => n7, B => add_92_G7_carry_11_port, 
                           CO => add_92_G7_carry_12_port, S => 
                           aMatrix_13_11_port);
   add_92_G7_U1_1_12 : HA_X1 port map( A => n8, B => add_92_G7_carry_12_port, 
                           CO => add_92_G7_carry_13_port, S => 
                           aMatrix_13_12_port);
   add_92_G7_U1_1_13 : HA_X1 port map( A => n9, B => add_92_G7_carry_13_port, 
                           CO => add_92_G7_carry_14_port, S => 
                           aMatrix_13_13_port);
   add_92_G7_U1_1_14 : HA_X1 port map( A => n10, B => add_92_G7_carry_14_port, 
                           CO => add_92_G7_carry_15_port, S => 
                           aMatrix_13_14_port);
   add_92_G7_U1_1_15 : HA_X1 port map( A => n11, B => add_92_G7_carry_15_port, 
                           CO => add_92_G7_carry_16_port, S => 
                           aMatrix_13_15_port);
   add_92_G7_U1_1_16 : HA_X1 port map( A => n12, B => add_92_G7_carry_16_port, 
                           CO => add_92_G7_carry_17_port, S => 
                           aMatrix_13_16_port);
   add_92_G7_U1_1_17 : HA_X1 port map( A => n13, B => add_92_G7_carry_17_port, 
                           CO => add_92_G7_carry_18_port, S => 
                           aMatrix_13_17_port);
   add_92_G7_U1_1_18 : HA_X1 port map( A => n14, B => add_92_G7_carry_18_port, 
                           CO => add_92_G7_carry_19_port, S => 
                           aMatrix_13_18_port);
   add_92_G7_U1_1_19 : HA_X1 port map( A => n15, B => add_92_G7_carry_19_port, 
                           CO => add_92_G7_carry_20_port, S => 
                           aMatrix_13_19_port);
   add_92_G7_U1_1_20 : HA_X1 port map( A => n16, B => add_92_G7_carry_20_port, 
                           CO => add_92_G7_carry_21_port, S => 
                           aMatrix_13_20_port);
   add_92_G6_U1_1_6 : HA_X1 port map( A => n3, B => n1, CO => 
                           add_92_G6_carry_7_port, S => aMatrix_11_6_port);
   add_92_G6_U1_1_7 : HA_X1 port map( A => n4, B => add_92_G6_carry_7_port, CO 
                           => add_92_G6_carry_8_port, S => aMatrix_11_7_port);
   add_92_G6_U1_1_8 : HA_X1 port map( A => n5, B => add_92_G6_carry_8_port, CO 
                           => add_92_G6_carry_9_port, S => aMatrix_11_8_port);
   add_92_G6_U1_1_9 : HA_X1 port map( A => n6, B => add_92_G6_carry_9_port, CO 
                           => add_92_G6_carry_10_port, S => aMatrix_11_9_port);
   add_92_G6_U1_1_10 : HA_X1 port map( A => n7, B => add_92_G6_carry_10_port, 
                           CO => add_92_G6_carry_11_port, S => 
                           aMatrix_11_10_port);
   add_92_G6_U1_1_11 : HA_X1 port map( A => n8, B => add_92_G6_carry_11_port, 
                           CO => add_92_G6_carry_12_port, S => 
                           aMatrix_11_11_port);
   add_92_G6_U1_1_12 : HA_X1 port map( A => n9, B => add_92_G6_carry_12_port, 
                           CO => add_92_G6_carry_13_port, S => 
                           aMatrix_11_12_port);
   add_92_G6_U1_1_13 : HA_X1 port map( A => n10, B => add_92_G6_carry_13_port, 
                           CO => add_92_G6_carry_14_port, S => 
                           aMatrix_11_13_port);
   add_92_G6_U1_1_14 : HA_X1 port map( A => n11, B => add_92_G6_carry_14_port, 
                           CO => add_92_G6_carry_15_port, S => 
                           aMatrix_11_14_port);
   add_92_G6_U1_1_15 : HA_X1 port map( A => n12, B => add_92_G6_carry_15_port, 
                           CO => add_92_G6_carry_16_port, S => 
                           aMatrix_11_15_port);
   add_92_G6_U1_1_16 : HA_X1 port map( A => n13, B => add_92_G6_carry_16_port, 
                           CO => add_92_G6_carry_17_port, S => 
                           aMatrix_11_16_port);
   add_92_G6_U1_1_17 : HA_X1 port map( A => n14, B => add_92_G6_carry_17_port, 
                           CO => add_92_G6_carry_18_port, S => 
                           aMatrix_11_17_port);
   add_92_G6_U1_1_18 : HA_X1 port map( A => n15, B => add_92_G6_carry_18_port, 
                           CO => add_92_G6_carry_19_port, S => 
                           aMatrix_11_18_port);
   add_92_G6_U1_1_19 : HA_X1 port map( A => n16, B => add_92_G6_carry_19_port, 
                           CO => add_92_G6_carry_20_port, S => 
                           aMatrix_11_19_port);
   add_92_G5_U1_1_5 : HA_X1 port map( A => n3, B => n1, CO => 
                           add_92_G5_carry_6_port, S => aMatrix_9_5_port);
   add_92_G5_U1_1_6 : HA_X1 port map( A => n4, B => add_92_G5_carry_6_port, CO 
                           => add_92_G5_carry_7_port, S => aMatrix_9_6_port);
   add_92_G5_U1_1_7 : HA_X1 port map( A => n5, B => add_92_G5_carry_7_port, CO 
                           => add_92_G5_carry_8_port, S => aMatrix_9_7_port);
   add_92_G5_U1_1_8 : HA_X1 port map( A => n6, B => add_92_G5_carry_8_port, CO 
                           => add_92_G5_carry_9_port, S => aMatrix_9_8_port);
   add_92_G5_U1_1_9 : HA_X1 port map( A => n7, B => add_92_G5_carry_9_port, CO 
                           => add_92_G5_carry_10_port, S => aMatrix_9_9_port);
   add_92_G5_U1_1_10 : HA_X1 port map( A => n8, B => add_92_G5_carry_10_port, 
                           CO => add_92_G5_carry_11_port, S => 
                           aMatrix_9_10_port);
   add_92_G5_U1_1_11 : HA_X1 port map( A => n9, B => add_92_G5_carry_11_port, 
                           CO => add_92_G5_carry_12_port, S => 
                           aMatrix_9_11_port);
   add_92_G5_U1_1_12 : HA_X1 port map( A => n10, B => add_92_G5_carry_12_port, 
                           CO => add_92_G5_carry_13_port, S => 
                           aMatrix_9_12_port);
   add_92_G5_U1_1_13 : HA_X1 port map( A => n11, B => add_92_G5_carry_13_port, 
                           CO => add_92_G5_carry_14_port, S => 
                           aMatrix_9_13_port);
   add_92_G5_U1_1_14 : HA_X1 port map( A => n12, B => add_92_G5_carry_14_port, 
                           CO => add_92_G5_carry_15_port, S => 
                           aMatrix_9_14_port);
   add_92_G5_U1_1_15 : HA_X1 port map( A => n13, B => add_92_G5_carry_15_port, 
                           CO => add_92_G5_carry_16_port, S => 
                           aMatrix_9_15_port);
   add_92_G5_U1_1_16 : HA_X1 port map( A => n14, B => add_92_G5_carry_16_port, 
                           CO => add_92_G5_carry_17_port, S => 
                           aMatrix_9_16_port);
   add_92_G5_U1_1_17 : HA_X1 port map( A => n15, B => add_92_G5_carry_17_port, 
                           CO => add_92_G5_carry_18_port, S => 
                           aMatrix_9_17_port);
   add_92_G5_U1_1_18 : HA_X1 port map( A => n16, B => add_92_G5_carry_18_port, 
                           CO => add_92_G5_carry_19_port, S => 
                           aMatrix_9_18_port);
   add_92_G4_U1_1_4 : HA_X1 port map( A => n3, B => n1, CO => 
                           add_92_G4_carry_5_port, S => aMatrix_7_4_port);
   add_92_G4_U1_1_5 : HA_X1 port map( A => n4, B => add_92_G4_carry_5_port, CO 
                           => add_92_G4_carry_6_port, S => aMatrix_7_5_port);
   add_92_G4_U1_1_6 : HA_X1 port map( A => n5, B => add_92_G4_carry_6_port, CO 
                           => add_92_G4_carry_7_port, S => aMatrix_7_6_port);
   add_92_G4_U1_1_7 : HA_X1 port map( A => n6, B => add_92_G4_carry_7_port, CO 
                           => add_92_G4_carry_8_port, S => aMatrix_7_7_port);
   add_92_G4_U1_1_8 : HA_X1 port map( A => n7, B => add_92_G4_carry_8_port, CO 
                           => add_92_G4_carry_9_port, S => aMatrix_7_8_port);
   add_92_G4_U1_1_9 : HA_X1 port map( A => n8, B => add_92_G4_carry_9_port, CO 
                           => add_92_G4_carry_10_port, S => aMatrix_7_9_port);
   add_92_G4_U1_1_10 : HA_X1 port map( A => n9, B => add_92_G4_carry_10_port, 
                           CO => add_92_G4_carry_11_port, S => 
                           aMatrix_7_10_port);
   add_92_G4_U1_1_11 : HA_X1 port map( A => n10, B => add_92_G4_carry_11_port, 
                           CO => add_92_G4_carry_12_port, S => 
                           aMatrix_7_11_port);
   add_92_G4_U1_1_12 : HA_X1 port map( A => n11, B => add_92_G4_carry_12_port, 
                           CO => add_92_G4_carry_13_port, S => 
                           aMatrix_7_12_port);
   add_92_G4_U1_1_13 : HA_X1 port map( A => n12, B => add_92_G4_carry_13_port, 
                           CO => add_92_G4_carry_14_port, S => 
                           aMatrix_7_13_port);
   add_92_G4_U1_1_14 : HA_X1 port map( A => n13, B => add_92_G4_carry_14_port, 
                           CO => add_92_G4_carry_15_port, S => 
                           aMatrix_7_14_port);
   add_92_G4_U1_1_15 : HA_X1 port map( A => n14, B => add_92_G4_carry_15_port, 
                           CO => add_92_G4_carry_16_port, S => 
                           aMatrix_7_15_port);
   add_92_G4_U1_1_16 : HA_X1 port map( A => n15, B => add_92_G4_carry_16_port, 
                           CO => add_92_G4_carry_17_port, S => 
                           aMatrix_7_16_port);
   add_92_G4_U1_1_17 : HA_X1 port map( A => n16, B => add_92_G4_carry_17_port, 
                           CO => add_92_G4_carry_18_port, S => 
                           aMatrix_7_17_port);
   add_92_G3_U1_1_3 : HA_X1 port map( A => n3, B => n1, CO => 
                           add_92_G3_carry_4_port, S => aMatrix_5_3_port);
   add_92_G3_U1_1_4 : HA_X1 port map( A => n4, B => add_92_G3_carry_4_port, CO 
                           => add_92_G3_carry_5_port, S => aMatrix_5_4_port);
   add_92_G3_U1_1_5 : HA_X1 port map( A => n5, B => add_92_G3_carry_5_port, CO 
                           => add_92_G3_carry_6_port, S => aMatrix_5_5_port);
   add_92_G3_U1_1_6 : HA_X1 port map( A => n6, B => add_92_G3_carry_6_port, CO 
                           => add_92_G3_carry_7_port, S => aMatrix_5_6_port);
   add_92_G3_U1_1_7 : HA_X1 port map( A => n7, B => add_92_G3_carry_7_port, CO 
                           => add_92_G3_carry_8_port, S => aMatrix_5_7_port);
   add_92_G3_U1_1_8 : HA_X1 port map( A => n8, B => add_92_G3_carry_8_port, CO 
                           => add_92_G3_carry_9_port, S => aMatrix_5_8_port);
   add_92_G3_U1_1_9 : HA_X1 port map( A => n9, B => add_92_G3_carry_9_port, CO 
                           => add_92_G3_carry_10_port, S => aMatrix_5_9_port);
   add_92_G3_U1_1_10 : HA_X1 port map( A => n10, B => add_92_G3_carry_10_port, 
                           CO => add_92_G3_carry_11_port, S => 
                           aMatrix_5_10_port);
   add_92_G3_U1_1_11 : HA_X1 port map( A => n11, B => add_92_G3_carry_11_port, 
                           CO => add_92_G3_carry_12_port, S => 
                           aMatrix_5_11_port);
   add_92_G3_U1_1_12 : HA_X1 port map( A => n12, B => add_92_G3_carry_12_port, 
                           CO => add_92_G3_carry_13_port, S => 
                           aMatrix_5_12_port);
   add_92_G3_U1_1_13 : HA_X1 port map( A => n13, B => add_92_G3_carry_13_port, 
                           CO => add_92_G3_carry_14_port, S => 
                           aMatrix_5_13_port);
   add_92_G3_U1_1_14 : HA_X1 port map( A => n14, B => add_92_G3_carry_14_port, 
                           CO => add_92_G3_carry_15_port, S => 
                           aMatrix_5_14_port);
   add_92_G3_U1_1_15 : HA_X1 port map( A => n15, B => add_92_G3_carry_15_port, 
                           CO => add_92_G3_carry_16_port, S => 
                           aMatrix_5_15_port);
   add_92_G3_U1_1_16 : HA_X1 port map( A => n16, B => add_92_G3_carry_16_port, 
                           CO => add_92_G3_carry_17_port, S => 
                           aMatrix_5_16_port);
   add_92_G2_U1_1_2 : HA_X1 port map( A => n3, B => n1, CO => 
                           add_92_G2_carry_3_port, S => aMatrix_3_2_port);
   add_92_G2_U1_1_3 : HA_X1 port map( A => n4, B => add_92_G2_carry_3_port, CO 
                           => add_92_G2_carry_4_port, S => aMatrix_3_3_port);
   add_92_G2_U1_1_4 : HA_X1 port map( A => n5, B => add_92_G2_carry_4_port, CO 
                           => add_92_G2_carry_5_port, S => aMatrix_3_4_port);
   add_92_G2_U1_1_5 : HA_X1 port map( A => n6, B => add_92_G2_carry_5_port, CO 
                           => add_92_G2_carry_6_port, S => aMatrix_3_5_port);
   add_92_G2_U1_1_6 : HA_X1 port map( A => n7, B => add_92_G2_carry_6_port, CO 
                           => add_92_G2_carry_7_port, S => aMatrix_3_6_port);
   add_92_G2_U1_1_7 : HA_X1 port map( A => n8, B => add_92_G2_carry_7_port, CO 
                           => add_92_G2_carry_8_port, S => aMatrix_3_7_port);
   add_92_G2_U1_1_8 : HA_X1 port map( A => n9, B => add_92_G2_carry_8_port, CO 
                           => add_92_G2_carry_9_port, S => aMatrix_3_8_port);
   add_92_G2_U1_1_9 : HA_X1 port map( A => n10, B => add_92_G2_carry_9_port, CO
                           => add_92_G2_carry_10_port, S => aMatrix_3_9_port);
   add_92_G2_U1_1_10 : HA_X1 port map( A => n11, B => add_92_G2_carry_10_port, 
                           CO => add_92_G2_carry_11_port, S => 
                           aMatrix_3_10_port);
   add_92_G2_U1_1_11 : HA_X1 port map( A => n12, B => add_92_G2_carry_11_port, 
                           CO => add_92_G2_carry_12_port, S => 
                           aMatrix_3_11_port);
   add_92_G2_U1_1_12 : HA_X1 port map( A => n13, B => add_92_G2_carry_12_port, 
                           CO => add_92_G2_carry_13_port, S => 
                           aMatrix_3_12_port);
   add_92_G2_U1_1_13 : HA_X1 port map( A => n14, B => add_92_G2_carry_13_port, 
                           CO => add_92_G2_carry_14_port, S => 
                           aMatrix_3_13_port);
   add_92_G2_U1_1_14 : HA_X1 port map( A => n15, B => add_92_G2_carry_14_port, 
                           CO => add_92_G2_carry_15_port, S => 
                           aMatrix_3_14_port);
   add_92_G2_U1_1_15 : HA_X1 port map( A => n16, B => add_92_G2_carry_15_port, 
                           CO => add_92_G2_carry_16_port, S => 
                           aMatrix_3_15_port);
   add_92_U1_1_1 : HA_X1 port map( A => n3, B => n1, CO => add_92_carry_2_port,
                           S => aMatrix_1_1_port);
   add_92_U1_1_2 : HA_X1 port map( A => n4, B => add_92_carry_2_port, CO => 
                           add_92_carry_3_port, S => aMatrix_1_2_port);
   add_92_U1_1_3 : HA_X1 port map( A => n5, B => add_92_carry_3_port, CO => 
                           add_92_carry_4_port, S => aMatrix_1_3_port);
   add_92_U1_1_4 : HA_X1 port map( A => n6, B => add_92_carry_4_port, CO => 
                           add_92_carry_5_port, S => aMatrix_1_4_port);
   add_92_U1_1_5 : HA_X1 port map( A => n7, B => add_92_carry_5_port, CO => 
                           add_92_carry_6_port, S => aMatrix_1_5_port);
   add_92_U1_1_6 : HA_X1 port map( A => n8, B => add_92_carry_6_port, CO => 
                           add_92_carry_7_port, S => aMatrix_1_6_port);
   add_92_U1_1_7 : HA_X1 port map( A => n9, B => add_92_carry_7_port, CO => 
                           add_92_carry_8_port, S => aMatrix_1_7_port);
   add_92_U1_1_8 : HA_X1 port map( A => n10, B => add_92_carry_8_port, CO => 
                           add_92_carry_9_port, S => aMatrix_1_8_port);
   add_92_U1_1_9 : HA_X1 port map( A => n11, B => add_92_carry_9_port, CO => 
                           add_92_carry_10_port, S => aMatrix_1_9_port);
   add_92_U1_1_10 : HA_X1 port map( A => n12, B => add_92_carry_10_port, CO => 
                           add_92_carry_11_port, S => aMatrix_1_10_port);
   add_92_U1_1_11 : HA_X1 port map( A => n13, B => add_92_carry_11_port, CO => 
                           add_92_carry_12_port, S => aMatrix_1_11_port);
   add_92_U1_1_12 : HA_X1 port map( A => n14, B => add_92_carry_12_port, CO => 
                           add_92_carry_13_port, S => aMatrix_1_12_port);
   add_92_U1_1_13 : HA_X1 port map( A => n15, B => add_92_carry_13_port, CO => 
                           add_92_carry_14_port, S => aMatrix_1_13_port);
   add_92_U1_1_14 : HA_X1 port map( A => n16, B => add_92_carry_14_port, CO => 
                           add_92_carry_15_port, S => aMatrix_1_14_port);
   U3 : NOR2_X2 port map( A1 => add_92_G4_carry_18_port, A2 => A(15), ZN => 
                           aMatrix_7_31_port);
   U4 : NOR2_X2 port map( A1 => add_92_G3_carry_17_port, A2 => A(15), ZN => 
                           aMatrix_5_31_port);
   U5 : NOR2_X2 port map( A1 => add_92_G2_carry_16_port, A2 => n17, ZN => 
                           aMatrix_3_31_port);
   U6 : BUF_X1 port map( A => n26, Z => n25);
   U7 : BUF_X1 port map( A => n26, Z => n24);
   U8 : BUF_X1 port map( A => n26, Z => n23);
   U9 : BUF_X1 port map( A => n28, Z => n26);
   U10 : BUF_X1 port map( A => n27, Z => n22);
   U11 : INV_X1 port map( A => n24, ZN => n18);
   U12 : INV_X1 port map( A => n23, ZN => n20);
   U13 : INV_X1 port map( A => n24, ZN => n19);
   U14 : INV_X1 port map( A => n25, ZN => n17);
   U15 : NOR2_X1 port map( A1 => add_92_G8_carry_22_port, A2 => n19, ZN => 
                           aMatrix_15_31_port);
   U16 : NOR2_X2 port map( A1 => add_92_carry_15_port, A2 => n18, ZN => 
                           aMatrix_1_31_port);
   U17 : NOR2_X2 port map( A1 => add_92_G5_carry_19_port, A2 => n18, ZN => 
                           aMatrix_9_31_port);
   U18 : NOR2_X1 port map( A1 => add_92_G6_carry_20_port, A2 => n19, ZN => 
                           aMatrix_11_31_port);
   U19 : NOR2_X1 port map( A1 => add_92_G7_carry_21_port, A2 => n21, ZN => 
                           aMatrix_13_31_port);
   U20 : INV_X1 port map( A => n22, ZN => n21);
   U21 : BUF_X1 port map( A => n28, Z => n27);
   U22 : INV_X1 port map( A => n3, ZN => n2);
   U23 : INV_X1 port map( A => A(0), ZN => n1);
   U24 : INV_X1 port map( A => A(1), ZN => n3);
   U25 : INV_X1 port map( A => A(2), ZN => n4);
   U26 : INV_X1 port map( A => A(3), ZN => n5);
   U27 : INV_X1 port map( A => A(4), ZN => n6);
   U28 : INV_X1 port map( A => A(5), ZN => n7);
   U29 : INV_X1 port map( A => A(6), ZN => n8);
   U30 : INV_X1 port map( A => A(7), ZN => n9);
   U31 : INV_X1 port map( A => A(8), ZN => n10);
   U32 : INV_X1 port map( A => A(9), ZN => n11);
   U33 : INV_X1 port map( A => A(10), ZN => n12);
   U34 : INV_X1 port map( A => A(11), ZN => n13);
   U35 : INV_X1 port map( A => A(12), ZN => n14);
   U36 : INV_X1 port map( A => A(13), ZN => n15);
   U37 : INV_X1 port map( A => A(14), ZN => n16);
   U38 : INV_X1 port map( A => A(15), ZN => n28);
   U39 : XOR2_X1 port map( A => add_92_carry_15_port, B => n25, Z => 
                           aMatrix_1_15_port);
   U40 : XOR2_X1 port map( A => add_92_G2_carry_16_port, B => n25, Z => 
                           aMatrix_3_16_port);
   U41 : XOR2_X1 port map( A => add_92_G3_carry_17_port, B => n25, Z => 
                           aMatrix_5_17_port);
   U42 : XOR2_X1 port map( A => add_92_G4_carry_18_port, B => n25, Z => 
                           aMatrix_7_18_port);
   U43 : XOR2_X1 port map( A => add_92_G5_carry_19_port, B => n25, Z => 
                           aMatrix_9_19_port);
   U44 : XOR2_X1 port map( A => add_92_G6_carry_20_port, B => n25, Z => 
                           aMatrix_11_20_port);
   U45 : XOR2_X1 port map( A => add_92_G7_carry_21_port, B => n25, Z => 
                           aMatrix_13_21_port);
   U46 : XOR2_X1 port map( A => add_92_G8_carry_22_port, B => n25, Z => 
                           aMatrix_15_22_port);
   n29 <= '0';
   aMatrix_3_0_port <= '0';
   aMatrix_5_0_port <= '0';
   aMatrix_7_0_port <= '0';
   aMatrix_9_0_port <= '0';
   aMatrix_11_0_port <= '0';
   aMatrix_13_0_port <= '0';
   aMatrix_15_0_port <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity P4_ADDER_N32_NB8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end P4_ADDER_N32_NB8;

architecture SYN_STRUCTURAL of P4_ADDER_N32_NB8 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GENERATOR_N32_NB8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_N32_NB8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Co :
            out std_logic_vector (7 downto 0));
   end component;
   
   signal CarriesOut_6_port, CarriesOut_5_port, CarriesOut_4_port, 
      CarriesOut_3_port, CarriesOut_2_port, CarriesOut_1_port, 
      CarriesOut_0_port, n1, n2 : std_logic;

begin
   
   CARRY_GENERATOR_INSTANCE : CARRY_GENERATOR_N32_NB8 port map( A(31) => A(31),
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => n2, B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => n1, Ci => Ci, Co(7) => 
                           Co, Co(6) => CarriesOut_6_port, Co(5) => 
                           CarriesOut_5_port, Co(4) => CarriesOut_4_port, Co(3)
                           => CarriesOut_3_port, Co(2) => CarriesOut_2_port, 
                           Co(1) => CarriesOut_1_port, Co(0) => 
                           CarriesOut_0_port);
   SUM_GENERATOR_INSTANCE : SUM_GENERATOR_N32_NB8 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => n2, B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => n1, Ci(7) => 
                           CarriesOut_6_port, Ci(6) => CarriesOut_5_port, Ci(5)
                           => CarriesOut_4_port, Ci(4) => CarriesOut_3_port, 
                           Ci(3) => CarriesOut_2_port, Ci(2) => 
                           CarriesOut_1_port, Ci(1) => CarriesOut_0_port, Ci(0)
                           => Ci, S(31) => S(31), S(30) => S(30), S(29) => 
                           S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   U1 : BUF_X1 port map( A => B(0), Z => n1);
   U2 : BUF_X1 port map( A => A(0), Z => n2);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_31 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_31;

architecture SYN_BEHAVIORAL of FFD_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n3, n4, n1, n2, n_1273 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n4, CK => CLK, Q => Q_port, QN => n_1273);
   U3 : NOR2_X1 port map( A1 => n3, A2 => n1, ZN => n4);
   U4 : INV_X1 port map( A => RST, ZN => n1);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n3)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_224 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_224;

architecture SYN_BEHAVIORAL of LD_224 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U4 : INV_X1 port map( A => EN, ZN => n1);
   U5 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FU_N5 is

   port( RS1, RS2, RD_MEM, RD_WB : in std_logic_vector (4 downto 0);  RF_WE_MEM
         , RF_WE_WB : in std_logic;  FORWARD_A, FORWARD_B : out 
         std_logic_vector (1 downto 0));

end FU_N5;

architecture SYN_BEHAVIORAL of FU_N5 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27 : std_logic;

begin
   
   U2 : INV_X1 port map( A => n1, ZN => FORWARD_A(0));
   U3 : INV_X1 port map( A => n2, ZN => FORWARD_B(0));
   U4 : NOR4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => 
                           FORWARD_B(1));
   U5 : XOR2_X1 port map( A => RS2(1), B => RD_WB(1), Z => n6);
   U6 : XOR2_X1 port map( A => RS2(4), B => RD_WB(4), Z => n5);
   U7 : XOR2_X1 port map( A => RS2(2), B => RD_WB(2), Z => n4);
   U8 : NAND4_X1 port map( A1 => n7, A2 => n8, A3 => RF_WE_WB, A4 => n2, ZN => 
                           n3);
   U9 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n2)
                           ;
   U10 : NOR3_X1 port map( A1 => n13, A2 => n14, A3 => n15, ZN => n12);
   U11 : XOR2_X1 port map( A => RS2(1), B => RD_MEM(1), Z => n15);
   U12 : XOR2_X1 port map( A => RS2(0), B => RD_MEM(0), Z => n13);
   U13 : XNOR2_X1 port map( A => RD_MEM(3), B => RS2(3), ZN => n11);
   U14 : XNOR2_X1 port map( A => RD_MEM(4), B => RS2(4), ZN => n10);
   U15 : XNOR2_X1 port map( A => RD_MEM(2), B => RS2(2), ZN => n9);
   U16 : XNOR2_X1 port map( A => RD_WB(3), B => RS2(3), ZN => n8);
   U17 : XNOR2_X1 port map( A => RD_WB(0), B => RS2(0), ZN => n7);
   U18 : NOR4_X1 port map( A1 => n16, A2 => n17, A3 => n18, A4 => n19, ZN => 
                           FORWARD_A(1));
   U19 : XOR2_X1 port map( A => RS1(1), B => RD_WB(1), Z => n19);
   U20 : XOR2_X1 port map( A => RS1(4), B => RD_WB(4), Z => n18);
   U21 : XOR2_X1 port map( A => RS1(2), B => RD_WB(2), Z => n17);
   U22 : NAND4_X1 port map( A1 => n20, A2 => n21, A3 => RF_WE_WB, A4 => n1, ZN 
                           => n16);
   U23 : NAND4_X1 port map( A1 => n22, A2 => n23, A3 => n24, A4 => n25, ZN => 
                           n1);
   U24 : NOR3_X1 port map( A1 => n26, A2 => n14, A3 => n27, ZN => n25);
   U25 : XOR2_X1 port map( A => RS1(1), B => RD_MEM(1), Z => n27);
   U26 : INV_X1 port map( A => RF_WE_MEM, ZN => n14);
   U27 : XOR2_X1 port map( A => RS1(0), B => RD_MEM(0), Z => n26);
   U28 : XNOR2_X1 port map( A => RD_MEM(3), B => RS1(3), ZN => n24);
   U29 : XNOR2_X1 port map( A => RD_MEM(4), B => RS1(4), ZN => n23);
   U30 : XNOR2_X1 port map( A => RD_MEM(2), B => RS1(2), ZN => n22);
   U31 : XNOR2_X1 port map( A => RD_WB(3), B => RS1(3), ZN => n21);
   U32 : XNOR2_X1 port map( A => RD_WB(0), B => RS1(0), ZN => n20);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ZERO_DETECTOR_N32_1 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic);

end ZERO_DETECTOR_N32_1;

architecture SYN_STRUCTURAL of ZERO_DETECTOR_N32_1 is

   component AND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, M_4_1_port, M_4_0_port, M_3_3_port, M_3_2_port, 
      M_3_1_port, M_3_0_port, M_2_7_port, M_2_6_port, M_2_5_port, M_2_4_port, 
      M_2_3_port, M_2_2_port, M_2_1_port, M_2_0_port, M_1_15_port, M_1_14_port,
      M_1_13_port, M_1_12_port, M_1_11_port, M_1_10_port, M_1_9_port, 
      M_1_8_port, M_1_7_port, M_1_6_port, M_1_5_port, M_1_4_port, M_1_3_port, 
      M_1_2_port, M_1_1_port, M_1_0_port, M_0_31_port, M_0_30_port, M_0_29_port
      , M_0_28_port, M_0_27_port, M_0_26_port, M_0_25_port, M_0_24_port, 
      M_0_23_port, M_0_22_port, M_0_21_port, M_0_20_port, M_0_19_port, 
      M_0_18_port, M_0_17_port, M_0_16_port, M_0_15_port, M_0_14_port, 
      M_0_13_port, M_0_12_port, M_0_11_port, M_0_10_port, M_0_9_port, 
      M_0_8_port, M_0_7_port, M_0_6_port, M_0_5_port, M_0_4_port, M_0_3_port, 
      M_0_2_port, M_0_1_port, M_0_0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   XOR0_i_0_0 : XNOR2_63 port map( A => A(0), B => X_Logic0_port, Y => 
                           M_0_0_port);
   XOR0_i_0_1 : XNOR2_62 port map( A => A(1), B => X_Logic0_port, Y => 
                           M_0_1_port);
   XOR0_i_0_2 : XNOR2_61 port map( A => A(2), B => X_Logic0_port, Y => 
                           M_0_2_port);
   XOR0_i_0_3 : XNOR2_60 port map( A => A(3), B => X_Logic0_port, Y => 
                           M_0_3_port);
   XOR0_i_0_4 : XNOR2_59 port map( A => A(4), B => X_Logic0_port, Y => 
                           M_0_4_port);
   XOR0_i_0_5 : XNOR2_58 port map( A => A(5), B => X_Logic0_port, Y => 
                           M_0_5_port);
   XOR0_i_0_6 : XNOR2_57 port map( A => A(6), B => X_Logic0_port, Y => 
                           M_0_6_port);
   XOR0_i_0_7 : XNOR2_56 port map( A => A(7), B => X_Logic0_port, Y => 
                           M_0_7_port);
   XOR0_i_0_8 : XNOR2_55 port map( A => A(8), B => X_Logic0_port, Y => 
                           M_0_8_port);
   XOR0_i_0_9 : XNOR2_54 port map( A => A(9), B => X_Logic0_port, Y => 
                           M_0_9_port);
   XOR0_i_0_10 : XNOR2_53 port map( A => A(10), B => X_Logic0_port, Y => 
                           M_0_10_port);
   XOR0_i_0_11 : XNOR2_52 port map( A => A(11), B => X_Logic0_port, Y => 
                           M_0_11_port);
   XOR0_i_0_12 : XNOR2_51 port map( A => A(12), B => X_Logic0_port, Y => 
                           M_0_12_port);
   XOR0_i_0_13 : XNOR2_50 port map( A => A(13), B => X_Logic0_port, Y => 
                           M_0_13_port);
   XOR0_i_0_14 : XNOR2_49 port map( A => A(14), B => X_Logic0_port, Y => 
                           M_0_14_port);
   XOR0_i_0_15 : XNOR2_48 port map( A => A(15), B => X_Logic0_port, Y => 
                           M_0_15_port);
   XOR0_i_0_16 : XNOR2_47 port map( A => A(16), B => X_Logic0_port, Y => 
                           M_0_16_port);
   XOR0_i_0_17 : XNOR2_46 port map( A => A(17), B => X_Logic0_port, Y => 
                           M_0_17_port);
   XOR0_i_0_18 : XNOR2_45 port map( A => A(18), B => X_Logic0_port, Y => 
                           M_0_18_port);
   XOR0_i_0_19 : XNOR2_44 port map( A => A(19), B => X_Logic0_port, Y => 
                           M_0_19_port);
   XOR0_i_0_20 : XNOR2_43 port map( A => A(20), B => X_Logic0_port, Y => 
                           M_0_20_port);
   XOR0_i_0_21 : XNOR2_42 port map( A => A(21), B => X_Logic0_port, Y => 
                           M_0_21_port);
   XOR0_i_0_22 : XNOR2_41 port map( A => A(22), B => X_Logic0_port, Y => 
                           M_0_22_port);
   XOR0_i_0_23 : XNOR2_40 port map( A => A(23), B => X_Logic0_port, Y => 
                           M_0_23_port);
   XOR0_i_0_24 : XNOR2_39 port map( A => A(24), B => X_Logic0_port, Y => 
                           M_0_24_port);
   XOR0_i_0_25 : XNOR2_38 port map( A => A(25), B => X_Logic0_port, Y => 
                           M_0_25_port);
   XOR0_i_0_26 : XNOR2_37 port map( A => A(26), B => X_Logic0_port, Y => 
                           M_0_26_port);
   XOR0_i_0_27 : XNOR2_36 port map( A => A(27), B => X_Logic0_port, Y => 
                           M_0_27_port);
   XOR0_i_0_28 : XNOR2_35 port map( A => A(28), B => X_Logic0_port, Y => 
                           M_0_28_port);
   XOR0_i_0_29 : XNOR2_34 port map( A => A(29), B => X_Logic0_port, Y => 
                           M_0_29_port);
   XOR0_i_0_30 : XNOR2_33 port map( A => A(30), B => X_Logic0_port, Y => 
                           M_0_30_port);
   XOR0_i_0_31 : XNOR2_32 port map( A => A(31), B => X_Logic0_port, Y => 
                           M_0_31_port);
   AND_i_1_0 : AND2_61 port map( A => M_0_0_port, B => M_0_1_port, Y => 
                           M_1_0_port);
   AND_i_1_1 : AND2_60 port map( A => M_0_2_port, B => M_0_3_port, Y => 
                           M_1_1_port);
   AND_i_1_2 : AND2_59 port map( A => M_0_4_port, B => M_0_5_port, Y => 
                           M_1_2_port);
   AND_i_1_3 : AND2_58 port map( A => M_0_6_port, B => M_0_7_port, Y => 
                           M_1_3_port);
   AND_i_1_4 : AND2_57 port map( A => M_0_8_port, B => M_0_9_port, Y => 
                           M_1_4_port);
   AND_i_1_5 : AND2_56 port map( A => M_0_10_port, B => M_0_11_port, Y => 
                           M_1_5_port);
   AND_i_1_6 : AND2_55 port map( A => M_0_12_port, B => M_0_13_port, Y => 
                           M_1_6_port);
   AND_i_1_7 : AND2_54 port map( A => M_0_14_port, B => M_0_15_port, Y => 
                           M_1_7_port);
   AND_i_1_8 : AND2_53 port map( A => M_0_16_port, B => M_0_17_port, Y => 
                           M_1_8_port);
   AND_i_1_9 : AND2_52 port map( A => M_0_18_port, B => M_0_19_port, Y => 
                           M_1_9_port);
   AND_i_1_10 : AND2_51 port map( A => M_0_20_port, B => M_0_21_port, Y => 
                           M_1_10_port);
   AND_i_1_11 : AND2_50 port map( A => M_0_22_port, B => M_0_23_port, Y => 
                           M_1_11_port);
   AND_i_1_12 : AND2_49 port map( A => M_0_24_port, B => M_0_25_port, Y => 
                           M_1_12_port);
   AND_i_1_13 : AND2_48 port map( A => M_0_26_port, B => M_0_27_port, Y => 
                           M_1_13_port);
   AND_i_1_14 : AND2_47 port map( A => M_0_28_port, B => M_0_29_port, Y => 
                           M_1_14_port);
   AND_i_1_15 : AND2_46 port map( A => M_0_30_port, B => M_0_31_port, Y => 
                           M_1_15_port);
   AND_i_2_0 : AND2_45 port map( A => M_1_0_port, B => M_1_1_port, Y => 
                           M_2_0_port);
   AND_i_2_1 : AND2_44 port map( A => M_1_2_port, B => M_1_3_port, Y => 
                           M_2_1_port);
   AND_i_2_2 : AND2_43 port map( A => M_1_4_port, B => M_1_5_port, Y => 
                           M_2_2_port);
   AND_i_2_3 : AND2_42 port map( A => M_1_6_port, B => M_1_7_port, Y => 
                           M_2_3_port);
   AND_i_2_4 : AND2_41 port map( A => M_1_8_port, B => M_1_9_port, Y => 
                           M_2_4_port);
   AND_i_2_5 : AND2_40 port map( A => M_1_10_port, B => M_1_11_port, Y => 
                           M_2_5_port);
   AND_i_2_6 : AND2_39 port map( A => M_1_12_port, B => M_1_13_port, Y => 
                           M_2_6_port);
   AND_i_2_7 : AND2_38 port map( A => M_1_14_port, B => M_1_15_port, Y => 
                           M_2_7_port);
   AND_i_3_0 : AND2_37 port map( A => M_2_0_port, B => M_2_1_port, Y => 
                           M_3_0_port);
   AND_i_3_1 : AND2_36 port map( A => M_2_2_port, B => M_2_3_port, Y => 
                           M_3_1_port);
   AND_i_3_2 : AND2_35 port map( A => M_2_4_port, B => M_2_5_port, Y => 
                           M_3_2_port);
   AND_i_3_3 : AND2_34 port map( A => M_2_6_port, B => M_2_7_port, Y => 
                           M_3_3_port);
   AND_i_4_0 : AND2_33 port map( A => M_3_0_port, B => M_3_1_port, Y => 
                           M_4_0_port);
   AND_i_4_1 : AND2_32 port map( A => M_3_2_port, B => M_3_3_port, Y => 
                           M_4_1_port);
   AND_i_5_0 : AND2_31 port map( A => M_4_0_port, B => M_4_1_port, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_320 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_320;

architecture SYN_BEHAVIORAL of MUX21_L_320 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n3);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_NB8 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
         std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);  Z
         : out std_logic);

end ALU_N32_NB8;

architecture SYN_BEHAVIORAL of ALU_N32_NB8 is

   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component ZERO_DETECTOR_N32_0
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic);
   end component;
   
   component COMPARATOR_N32
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic_vector 
            (3 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component LOGIC_N32
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic_vector 
            (1 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component BARREL_SHIFTER_RIGHT_N32
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component BARREL_SHIFTER_LEFT_N32
      port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector
            (31 downto 0));
   end component;
   
   component BOOTH_MULTIPLIER_N32
      port( A, B : in std_logic_vector (15 downto 0);  P : out std_logic_vector
            (31 downto 0));
   end component;
   
   component P4_ADDER_N32_NB8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal Y_31_port, Y_30_port, Y_29_port, Y_28_port, Y_27_port, Y_26_port, 
      Y_25_port, Y_24_port, Y_23_port, Y_22_port, Y_21_port, Y_20_port, 
      Y_19_port, Y_18_port, Y_17_port, Y_16_port, Y_15_port, Y_14_port, 
      Y_13_port, Y_12_port, Y_11_port, Y_10_port, Y_9_port, Y_8_port, Y_7_port,
      Y_6_port, Y_5_port, Y_4_port, Y_3_port, Y_2_port, Y_1_port, Y_0_port, N96
      , OP_A_31_port, OP_A_30_port, OP_A_29_port, OP_A_28_port, OP_A_27_port, 
      OP_A_26_port, OP_A_25_port, OP_A_24_port, OP_A_23_port, OP_A_22_port, 
      OP_A_21_port, OP_A_20_port, OP_A_19_port, OP_A_18_port, OP_A_17_port, 
      OP_A_16_port, OP_A_15_port, OP_A_14_port, OP_A_13_port, OP_A_12_port, 
      OP_A_11_port, OP_A_10_port, OP_A_9_port, OP_A_8_port, OP_A_7_port, 
      OP_A_6_port, OP_A_5_port, OP_A_4_port, OP_A_3_port, OP_A_2_port, 
      OP_A_1_port, OP_A_0_port, OP_B_31_port, OP_B_30_port, OP_B_29_port, 
      OP_B_28_port, OP_B_27_port, OP_B_26_port, OP_B_25_port, OP_B_24_port, 
      OP_B_23_port, OP_B_22_port, OP_B_21_port, OP_B_20_port, OP_B_19_port, 
      OP_B_18_port, OP_B_17_port, OP_B_16_port, OP_B_15_port, OP_B_14_port, 
      OP_B_13_port, OP_B_12_port, OP_B_11_port, OP_B_10_port, OP_B_9_port, 
      OP_B_8_port, OP_B_7_port, OP_B_6_port, OP_B_5_port, OP_B_4_port, 
      OP_B_3_port, OP_B_2_port, OP_B_1_port, OP_B_0_port, Y_SHIFTL_31_port, 
      Y_SHIFTL_30_port, Y_SHIFTL_29_port, Y_SHIFTL_28_port, Y_SHIFTL_27_port, 
      Y_SHIFTL_26_port, Y_SHIFTL_25_port, Y_SHIFTL_24_port, Y_SHIFTL_23_port, 
      Y_SHIFTL_22_port, Y_SHIFTL_21_port, Y_SHIFTL_20_port, Y_SHIFTL_19_port, 
      Y_SHIFTL_18_port, Y_SHIFTL_17_port, Y_SHIFTL_16_port, Y_SHIFTL_15_port, 
      Y_SHIFTL_14_port, Y_SHIFTL_13_port, Y_SHIFTL_12_port, Y_SHIFTL_11_port, 
      Y_SHIFTL_10_port, Y_SHIFTL_9_port, Y_SHIFTL_8_port, Y_SHIFTL_7_port, 
      Y_SHIFTL_6_port, Y_SHIFTL_5_port, Y_SHIFTL_4_port, Y_SHIFTL_3_port, 
      Y_SHIFTL_2_port, Y_SHIFTL_1_port, Y_SHIFTL_0_port, Y_MUL_31_port, 
      Y_MUL_30_port, Y_MUL_29_port, Y_MUL_28_port, Y_MUL_27_port, Y_MUL_26_port
      , Y_MUL_25_port, Y_MUL_24_port, Y_MUL_23_port, Y_MUL_22_port, 
      Y_MUL_21_port, Y_MUL_20_port, Y_MUL_19_port, Y_MUL_18_port, Y_MUL_17_port
      , Y_MUL_16_port, Y_MUL_15_port, Y_MUL_14_port, Y_MUL_13_port, 
      Y_MUL_12_port, Y_MUL_11_port, Y_MUL_10_port, Y_MUL_9_port, Y_MUL_8_port, 
      Y_MUL_7_port, Y_MUL_6_port, Y_MUL_5_port, Y_MUL_4_port, Y_MUL_3_port, 
      Y_MUL_2_port, Y_MUL_1_port, Y_MUL_0_port, OP_Ci, Y_SUM_31_port, 
      Y_SUM_30_port, Y_SUM_29_port, Y_SUM_28_port, Y_SUM_27_port, Y_SUM_26_port
      , Y_SUM_25_port, Y_SUM_24_port, Y_SUM_23_port, Y_SUM_22_port, 
      Y_SUM_21_port, Y_SUM_20_port, Y_SUM_19_port, Y_SUM_18_port, Y_SUM_17_port
      , Y_SUM_16_port, Y_SUM_15_port, Y_SUM_14_port, Y_SUM_13_port, 
      Y_SUM_12_port, Y_SUM_11_port, Y_SUM_10_port, Y_SUM_9_port, Y_SUM_8_port, 
      Y_SUM_7_port, Y_SUM_6_port, Y_SUM_5_port, Y_SUM_4_port, Y_SUM_3_port, 
      Y_SUM_2_port, Y_SUM_1_port, Y_SUM_0_port, OP_LOGIC_1_port, 
      OP_LOGIC_0_port, Y_LOGIC_31_port, Y_LOGIC_30_port, Y_LOGIC_29_port, 
      Y_LOGIC_28_port, Y_LOGIC_27_port, Y_LOGIC_26_port, Y_LOGIC_25_port, 
      Y_LOGIC_24_port, Y_LOGIC_23_port, Y_LOGIC_22_port, Y_LOGIC_21_port, 
      Y_LOGIC_20_port, Y_LOGIC_19_port, Y_LOGIC_18_port, Y_LOGIC_17_port, 
      Y_LOGIC_16_port, Y_LOGIC_15_port, Y_LOGIC_14_port, Y_LOGIC_13_port, 
      Y_LOGIC_12_port, Y_LOGIC_11_port, Y_LOGIC_10_port, Y_LOGIC_9_port, 
      Y_LOGIC_8_port, Y_LOGIC_7_port, Y_LOGIC_6_port, Y_LOGIC_5_port, 
      Y_LOGIC_4_port, Y_LOGIC_3_port, Y_LOGIC_2_port, Y_LOGIC_1_port, 
      Y_LOGIC_0_port, OP_SHIFT, Y_SHIFTR_31_port, Y_SHIFTR_30_port, 
      Y_SHIFTR_29_port, Y_SHIFTR_28_port, Y_SHIFTR_27_port, Y_SHIFTR_26_port, 
      Y_SHIFTR_25_port, Y_SHIFTR_24_port, Y_SHIFTR_23_port, Y_SHIFTR_22_port, 
      Y_SHIFTR_21_port, Y_SHIFTR_20_port, Y_SHIFTR_19_port, Y_SHIFTR_18_port, 
      Y_SHIFTR_17_port, Y_SHIFTR_16_port, Y_SHIFTR_15_port, Y_SHIFTR_14_port, 
      Y_SHIFTR_13_port, Y_SHIFTR_12_port, Y_SHIFTR_11_port, Y_SHIFTR_10_port, 
      Y_SHIFTR_9_port, Y_SHIFTR_8_port, Y_SHIFTR_7_port, Y_SHIFTR_6_port, 
      Y_SHIFTR_5_port, Y_SHIFTR_4_port, Y_SHIFTR_3_port, Y_SHIFTR_2_port, 
      Y_SHIFTR_1_port, Y_SHIFTR_0_port, OP_COMPARE_3_port, OP_COMPARE_2_port, 
      OP_COMPARE_1_port, OP_COMPARE_0_port, Y_COMPARE_0_port, N246, N247, N248,
      N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, 
      N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, 
      N273, N274, N275, N276, N277, N278, N280, N281, N285, N286, N287, N288, 
      N289, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96_port, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246_port, n247_port, n248_port, n249_port, n250_port, n251_port, 
      n252_port, n253_port, n254_port, n255_port, n256_port, n257_port, 
      n258_port, n259_port, n260_port, n261_port, n262_port, n263_port, 
      n264_port, n265_port, n266_port, n267_port, n268_port, n269_port, 
      n270_port, n271_port, n272_port, n273_port, n274_port, n275_port, 
      n276_port, n277_port, n278_port, n279, n280_port, n281_port, n282, n283, 
      n284, n285_port, n286_port, n287_port, n288_port, n289_port, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n_1274, n_1275, n_1276, n_1277,
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305 : std_logic;

begin
   Y <= ( Y_31_port, Y_30_port, Y_29_port, Y_28_port, Y_27_port, Y_26_port, 
      Y_25_port, Y_24_port, Y_23_port, Y_22_port, Y_21_port, Y_20_port, 
      Y_19_port, Y_18_port, Y_17_port, Y_16_port, Y_15_port, Y_14_port, 
      Y_13_port, Y_12_port, Y_11_port, Y_10_port, Y_9_port, Y_8_port, Y_7_port,
      Y_6_port, Y_5_port, Y_4_port, Y_3_port, Y_2_port, Y_1_port, Y_0_port );
   
   OP_COMPARE_reg_3_inst : DLH_X1 port map( G => N285, D => N289, Q => 
                           OP_COMPARE_3_port);
   OP_COMPARE_reg_2_inst : DLH_X1 port map( G => N285, D => N288, Q => 
                           OP_COMPARE_2_port);
   OP_COMPARE_reg_1_inst : DLH_X1 port map( G => N285, D => N287, Q => 
                           OP_COMPARE_1_port);
   OP_COMPARE_reg_0_inst : DLH_X1 port map( G => N285, D => N286, Q => 
                           OP_COMPARE_0_port);
   OP_A_reg_31_inst : DLH_X1 port map( G => n35, D => OP1(31), Q => 
                           OP_A_31_port);
   OP_A_reg_30_inst : DLH_X1 port map( G => n35, D => OP1(30), Q => 
                           OP_A_30_port);
   OP_A_reg_29_inst : DLH_X1 port map( G => n35, D => OP1(29), Q => 
                           OP_A_29_port);
   OP_A_reg_28_inst : DLH_X1 port map( G => n35, D => OP1(28), Q => 
                           OP_A_28_port);
   OP_A_reg_27_inst : DLH_X1 port map( G => n35, D => OP1(27), Q => 
                           OP_A_27_port);
   OP_A_reg_26_inst : DLH_X1 port map( G => n35, D => OP1(26), Q => 
                           OP_A_26_port);
   OP_A_reg_25_inst : DLH_X1 port map( G => n35, D => OP1(25), Q => 
                           OP_A_25_port);
   OP_A_reg_24_inst : DLH_X1 port map( G => n35, D => OP1(24), Q => 
                           OP_A_24_port);
   OP_A_reg_23_inst : DLH_X1 port map( G => n35, D => OP1(23), Q => 
                           OP_A_23_port);
   OP_A_reg_22_inst : DLH_X1 port map( G => n35, D => OP1(22), Q => 
                           OP_A_22_port);
   OP_A_reg_21_inst : DLH_X1 port map( G => n36, D => OP1(21), Q => 
                           OP_A_21_port);
   OP_A_reg_20_inst : DLH_X1 port map( G => n36, D => OP1(20), Q => 
                           OP_A_20_port);
   OP_A_reg_19_inst : DLH_X1 port map( G => n36, D => OP1(19), Q => 
                           OP_A_19_port);
   OP_A_reg_18_inst : DLH_X1 port map( G => n36, D => OP1(18), Q => 
                           OP_A_18_port);
   OP_A_reg_17_inst : DLH_X1 port map( G => n36, D => OP1(17), Q => 
                           OP_A_17_port);
   OP_A_reg_16_inst : DLH_X1 port map( G => n36, D => OP1(16), Q => 
                           OP_A_16_port);
   OP_A_reg_15_inst : DLH_X1 port map( G => n36, D => OP1(15), Q => 
                           OP_A_15_port);
   OP_A_reg_14_inst : DLH_X1 port map( G => n36, D => OP1(14), Q => 
                           OP_A_14_port);
   OP_A_reg_13_inst : DLH_X1 port map( G => n36, D => OP1(13), Q => 
                           OP_A_13_port);
   OP_A_reg_12_inst : DLH_X1 port map( G => n36, D => OP1(12), Q => 
                           OP_A_12_port);
   OP_A_reg_11_inst : DLH_X1 port map( G => n37, D => OP1(11), Q => 
                           OP_A_11_port);
   OP_A_reg_10_inst : DLH_X1 port map( G => n37, D => OP1(10), Q => 
                           OP_A_10_port);
   OP_A_reg_9_inst : DLH_X1 port map( G => n37, D => OP1(9), Q => OP_A_9_port);
   OP_A_reg_8_inst : DLH_X1 port map( G => n37, D => OP1(8), Q => OP_A_8_port);
   OP_A_reg_7_inst : DLH_X1 port map( G => n37, D => OP1(7), Q => OP_A_7_port);
   OP_A_reg_6_inst : DLH_X1 port map( G => n37, D => OP1(6), Q => OP_A_6_port);
   OP_A_reg_5_inst : DLH_X1 port map( G => n37, D => OP1(5), Q => OP_A_5_port);
   OP_A_reg_4_inst : DLH_X1 port map( G => n37, D => OP1(4), Q => OP_A_4_port);
   OP_A_reg_3_inst : DLH_X1 port map( G => n37, D => OP1(3), Q => OP_A_3_port);
   OP_A_reg_2_inst : DLH_X1 port map( G => n37, D => OP1(2), Q => OP_A_2_port);
   OP_A_reg_1_inst : DLH_X1 port map( G => n38, D => OP1(1), Q => OP_A_1_port);
   OP_A_reg_0_inst : DLH_X1 port map( G => n38, D => OP1(0), Q => OP_A_0_port);
   OP_B_reg_31_inst : DLH_X1 port map( G => n38, D => N278, Q => OP_B_31_port);
   OP_B_reg_30_inst : DLH_X1 port map( G => n38, D => N277, Q => OP_B_30_port);
   OP_B_reg_29_inst : DLH_X1 port map( G => n38, D => N276, Q => OP_B_29_port);
   OP_B_reg_28_inst : DLH_X1 port map( G => n38, D => N275, Q => OP_B_28_port);
   OP_B_reg_27_inst : DLH_X1 port map( G => n38, D => N274, Q => OP_B_27_port);
   OP_B_reg_26_inst : DLH_X1 port map( G => n38, D => N273, Q => OP_B_26_port);
   OP_B_reg_25_inst : DLH_X1 port map( G => n38, D => N272, Q => OP_B_25_port);
   OP_B_reg_24_inst : DLH_X1 port map( G => n38, D => N271, Q => OP_B_24_port);
   OP_B_reg_23_inst : DLH_X1 port map( G => n39, D => N270, Q => OP_B_23_port);
   OP_B_reg_22_inst : DLH_X1 port map( G => n39, D => N269, Q => OP_B_22_port);
   OP_B_reg_21_inst : DLH_X1 port map( G => n39, D => N268, Q => OP_B_21_port);
   OP_B_reg_20_inst : DLH_X1 port map( G => n39, D => N267, Q => OP_B_20_port);
   OP_B_reg_19_inst : DLH_X1 port map( G => n39, D => N266, Q => OP_B_19_port);
   OP_B_reg_18_inst : DLH_X1 port map( G => n39, D => N265, Q => OP_B_18_port);
   OP_B_reg_17_inst : DLH_X1 port map( G => n39, D => N264, Q => OP_B_17_port);
   OP_B_reg_16_inst : DLH_X1 port map( G => n39, D => N263, Q => OP_B_16_port);
   OP_B_reg_15_inst : DLH_X1 port map( G => n39, D => N262, Q => OP_B_15_port);
   OP_B_reg_14_inst : DLH_X1 port map( G => n39, D => N261, Q => OP_B_14_port);
   OP_B_reg_13_inst : DLH_X1 port map( G => n40, D => N260, Q => OP_B_13_port);
   OP_B_reg_12_inst : DLH_X1 port map( G => n40, D => N259, Q => OP_B_12_port);
   OP_B_reg_11_inst : DLH_X1 port map( G => n40, D => N258, Q => OP_B_11_port);
   OP_B_reg_10_inst : DLH_X1 port map( G => n40, D => N257, Q => OP_B_10_port);
   OP_B_reg_9_inst : DLH_X1 port map( G => n40, D => N256, Q => OP_B_9_port);
   OP_B_reg_8_inst : DLH_X1 port map( G => n40, D => N255, Q => OP_B_8_port);
   OP_B_reg_7_inst : DLH_X1 port map( G => n40, D => N254, Q => OP_B_7_port);
   OP_B_reg_6_inst : DLH_X1 port map( G => n40, D => N253, Q => OP_B_6_port);
   OP_B_reg_5_inst : DLH_X1 port map( G => n40, D => N252, Q => OP_B_5_port);
   OP_B_reg_4_inst : DLH_X1 port map( G => n40, D => N251, Q => OP_B_4_port);
   OP_B_reg_3_inst : DLH_X1 port map( G => n41, D => N250, Q => OP_B_3_port);
   OP_B_reg_2_inst : DLH_X1 port map( G => n41, D => N249, Q => OP_B_2_port);
   OP_B_reg_1_inst : DLH_X1 port map( G => n41, D => N248, Q => OP_B_1_port);
   OP_B_reg_0_inst : DLH_X1 port map( G => n41, D => N247, Q => OP_B_0_port);
   OP_Ci_reg : DLH_X1 port map( G => n33, D => N280, Q => OP_Ci);
   OP_LOGIC_reg_1_inst : DLH_X1 port map( G => n30, D => n282, Q => 
                           OP_LOGIC_1_port);
   OP_LOGIC_reg_0_inst : DLH_X1 port map( G => n30, D => n283, Q => 
                           OP_LOGIC_0_port);
   OP_SHIFT_reg : DLL_X1 port map( D => N96, GN => n225, Q => OP_SHIFT);
   U301 : NAND3_X1 port map( A1 => n214, A2 => n287_port, A3 => n215, ZN => 
                           n212);
   U302 : NAND3_X1 port map( A1 => n200, A2 => n201, A3 => n222, ZN => N281);
   U303 : NAND3_X1 port map( A1 => OPC(2), A2 => n289_port, A3 => n216, ZN => 
                           n231);
   U304 : NAND3_X1 port map( A1 => OPC(6), A2 => n297, A3 => OPC(4), ZN => n187
                           );
   U305 : XOR2_X1 port map( A => OPC(2), B => OPC(3), Z => n233);
   U306 : NAND3_X1 port map( A1 => n297, A2 => n294, A3 => n298, ZN => n189);
   U307 : NAND3_X1 port map( A1 => n290, A2 => n281_port, A3 => n224, ZN => 
                           n214);
   U308 : NAND3_X1 port map( A1 => n298, A2 => n294, A3 => OPC(5), ZN => n226);
   U309 : NAND3_X1 port map( A1 => OPC(3), A2 => n224, A3 => OPC(0), ZN => n190
                           );
   SUM : P4_ADDER_N32_NB8 port map( A(31) => OP_A_31_port, A(30) => 
                           OP_A_30_port, A(29) => OP_A_29_port, A(28) => 
                           OP_A_28_port, A(27) => OP_A_27_port, A(26) => 
                           OP_A_26_port, A(25) => OP_A_25_port, A(24) => 
                           OP_A_24_port, A(23) => OP_A_23_port, A(22) => 
                           OP_A_22_port, A(21) => OP_A_21_port, A(20) => 
                           OP_A_20_port, A(19) => OP_A_19_port, A(18) => 
                           OP_A_18_port, A(17) => OP_A_17_port, A(16) => 
                           OP_A_16_port, A(15) => n245, A(14) => n244, A(13) =>
                           n243, A(12) => n242, A(11) => n241, A(10) => n240, 
                           A(9) => n239, A(8) => n238, A(7) => n237, A(6) => 
                           n236, A(5) => n235, A(4) => n234, A(3) => n54, A(2) 
                           => n53, A(1) => n52, A(0) => n51, B(31) => 
                           OP_B_31_port, B(30) => OP_B_30_port, B(29) => 
                           OP_B_29_port, B(28) => OP_B_28_port, B(27) => 
                           OP_B_27_port, B(26) => OP_B_26_port, B(25) => 
                           OP_B_25_port, B(24) => OP_B_24_port, B(23) => 
                           OP_B_23_port, B(22) => OP_B_22_port, B(21) => 
                           OP_B_21_port, B(20) => OP_B_20_port, B(19) => 
                           OP_B_19_port, B(18) => OP_B_18_port, B(17) => 
                           OP_B_17_port, B(16) => OP_B_16_port, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n50, B(3) => n49, B(2) => n48, 
                           B(1) => n47, B(0) => n46, Ci => OP_Ci, S(31) => 
                           Y_SUM_31_port, S(30) => Y_SUM_30_port, S(29) => 
                           Y_SUM_29_port, S(28) => Y_SUM_28_port, S(27) => 
                           Y_SUM_27_port, S(26) => Y_SUM_26_port, S(25) => 
                           Y_SUM_25_port, S(24) => Y_SUM_24_port, S(23) => 
                           Y_SUM_23_port, S(22) => Y_SUM_22_port, S(21) => 
                           Y_SUM_21_port, S(20) => Y_SUM_20_port, S(19) => 
                           Y_SUM_19_port, S(18) => Y_SUM_18_port, S(17) => 
                           Y_SUM_17_port, S(16) => Y_SUM_16_port, S(15) => 
                           Y_SUM_15_port, S(14) => Y_SUM_14_port, S(13) => 
                           Y_SUM_13_port, S(12) => Y_SUM_12_port, S(11) => 
                           Y_SUM_11_port, S(10) => Y_SUM_10_port, S(9) => 
                           Y_SUM_9_port, S(8) => Y_SUM_8_port, S(7) => 
                           Y_SUM_7_port, S(6) => Y_SUM_6_port, S(5) => 
                           Y_SUM_5_port, S(4) => Y_SUM_4_port, S(3) => 
                           Y_SUM_3_port, S(2) => Y_SUM_2_port, S(1) => 
                           Y_SUM_1_port, S(0) => Y_SUM_0_port, Co => n_1274);
   MUL : BOOTH_MULTIPLIER_N32 port map( A(15) => n245, A(14) => n244, A(13) => 
                           n243, A(12) => n242, A(11) => n241, A(10) => n240, 
                           A(9) => n239, A(8) => n238, A(7) => n237, A(6) => 
                           n236, A(5) => n235, A(4) => n234, A(3) => n54, A(2) 
                           => n53, A(1) => n52, A(0) => n51, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n50, B(3) => n49, B(2) => n48, 
                           B(1) => n47, B(0) => n46, P(31) => Y_MUL_31_port, 
                           P(30) => Y_MUL_30_port, P(29) => Y_MUL_29_port, 
                           P(28) => Y_MUL_28_port, P(27) => Y_MUL_27_port, 
                           P(26) => Y_MUL_26_port, P(25) => Y_MUL_25_port, 
                           P(24) => Y_MUL_24_port, P(23) => Y_MUL_23_port, 
                           P(22) => Y_MUL_22_port, P(21) => Y_MUL_21_port, 
                           P(20) => Y_MUL_20_port, P(19) => Y_MUL_19_port, 
                           P(18) => Y_MUL_18_port, P(17) => Y_MUL_17_port, 
                           P(16) => Y_MUL_16_port, P(15) => Y_MUL_15_port, 
                           P(14) => Y_MUL_14_port, P(13) => Y_MUL_13_port, 
                           P(12) => Y_MUL_12_port, P(11) => Y_MUL_11_port, 
                           P(10) => Y_MUL_10_port, P(9) => Y_MUL_9_port, P(8) 
                           => Y_MUL_8_port, P(7) => Y_MUL_7_port, P(6) => 
                           Y_MUL_6_port, P(5) => Y_MUL_5_port, P(4) => 
                           Y_MUL_4_port, P(3) => Y_MUL_3_port, P(2) => 
                           Y_MUL_2_port, P(1) => Y_MUL_1_port, P(0) => 
                           Y_MUL_0_port);
   BSL : BARREL_SHIFTER_LEFT_N32 port map( A(31) => OP_A_31_port, A(30) => 
                           OP_A_30_port, A(29) => OP_A_29_port, A(28) => 
                           OP_A_28_port, A(27) => OP_A_27_port, A(26) => 
                           OP_A_26_port, A(25) => OP_A_25_port, A(24) => 
                           OP_A_24_port, A(23) => OP_A_23_port, A(22) => 
                           OP_A_22_port, A(21) => OP_A_21_port, A(20) => 
                           OP_A_20_port, A(19) => OP_A_19_port, A(18) => 
                           OP_A_18_port, A(17) => OP_A_17_port, A(16) => 
                           OP_A_16_port, A(15) => n245, A(14) => n244, A(13) =>
                           n243, A(12) => n242, A(11) => n241, A(10) => n240, 
                           A(9) => n239, A(8) => n238, A(7) => n237, A(6) => 
                           n236, A(5) => n235, A(4) => n234, A(3) => n54, A(2) 
                           => n53, A(1) => n52, A(0) => n51, B(31) => 
                           OP_B_31_port, B(30) => OP_B_30_port, B(29) => 
                           OP_B_29_port, B(28) => OP_B_28_port, B(27) => 
                           OP_B_27_port, B(26) => OP_B_26_port, B(25) => 
                           OP_B_25_port, B(24) => OP_B_24_port, B(23) => 
                           OP_B_23_port, B(22) => OP_B_22_port, B(21) => 
                           OP_B_21_port, B(20) => OP_B_20_port, B(19) => 
                           OP_B_19_port, B(18) => OP_B_18_port, B(17) => 
                           OP_B_17_port, B(16) => OP_B_16_port, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n50, B(3) => n49, B(2) => n48, 
                           B(1) => n47, B(0) => n46, Y(31) => Y_SHIFTL_31_port,
                           Y(30) => Y_SHIFTL_30_port, Y(29) => Y_SHIFTL_29_port
                           , Y(28) => Y_SHIFTL_28_port, Y(27) => 
                           Y_SHIFTL_27_port, Y(26) => Y_SHIFTL_26_port, Y(25) 
                           => Y_SHIFTL_25_port, Y(24) => Y_SHIFTL_24_port, 
                           Y(23) => Y_SHIFTL_23_port, Y(22) => Y_SHIFTL_22_port
                           , Y(21) => Y_SHIFTL_21_port, Y(20) => 
                           Y_SHIFTL_20_port, Y(19) => Y_SHIFTL_19_port, Y(18) 
                           => Y_SHIFTL_18_port, Y(17) => Y_SHIFTL_17_port, 
                           Y(16) => Y_SHIFTL_16_port, Y(15) => Y_SHIFTL_15_port
                           , Y(14) => Y_SHIFTL_14_port, Y(13) => 
                           Y_SHIFTL_13_port, Y(12) => Y_SHIFTL_12_port, Y(11) 
                           => Y_SHIFTL_11_port, Y(10) => Y_SHIFTL_10_port, Y(9)
                           => Y_SHIFTL_9_port, Y(8) => Y_SHIFTL_8_port, Y(7) =>
                           Y_SHIFTL_7_port, Y(6) => Y_SHIFTL_6_port, Y(5) => 
                           Y_SHIFTL_5_port, Y(4) => Y_SHIFTL_4_port, Y(3) => 
                           Y_SHIFTL_3_port, Y(2) => Y_SHIFTL_2_port, Y(1) => 
                           Y_SHIFTL_1_port, Y(0) => Y_SHIFTL_0_port);
   BSR : BARREL_SHIFTER_RIGHT_N32 port map( A(31) => OP_A_31_port, A(30) => 
                           OP_A_30_port, A(29) => OP_A_29_port, A(28) => 
                           OP_A_28_port, A(27) => OP_A_27_port, A(26) => 
                           OP_A_26_port, A(25) => OP_A_25_port, A(24) => 
                           OP_A_24_port, A(23) => OP_A_23_port, A(22) => 
                           OP_A_22_port, A(21) => OP_A_21_port, A(20) => 
                           OP_A_20_port, A(19) => OP_A_19_port, A(18) => 
                           OP_A_18_port, A(17) => OP_A_17_port, A(16) => 
                           OP_A_16_port, A(15) => n245, A(14) => n244, A(13) =>
                           n243, A(12) => n242, A(11) => n241, A(10) => n240, 
                           A(9) => n239, A(8) => n238, A(7) => n237, A(6) => 
                           n236, A(5) => n235, A(4) => n234, A(3) => n54, A(2) 
                           => n53, A(1) => n52, A(0) => n51, B(31) => 
                           OP_B_31_port, B(30) => OP_B_30_port, B(29) => 
                           OP_B_29_port, B(28) => OP_B_28_port, B(27) => 
                           OP_B_27_port, B(26) => OP_B_26_port, B(25) => 
                           OP_B_25_port, B(24) => OP_B_24_port, B(23) => 
                           OP_B_23_port, B(22) => OP_B_22_port, B(21) => 
                           OP_B_21_port, B(20) => OP_B_20_port, B(19) => 
                           OP_B_19_port, B(18) => OP_B_18_port, B(17) => 
                           OP_B_17_port, B(16) => OP_B_16_port, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n50, B(3) => n49, B(2) => n48, 
                           B(1) => n47, B(0) => n46, S => OP_SHIFT, Y(31) => 
                           Y_SHIFTR_31_port, Y(30) => Y_SHIFTR_30_port, Y(29) 
                           => Y_SHIFTR_29_port, Y(28) => Y_SHIFTR_28_port, 
                           Y(27) => Y_SHIFTR_27_port, Y(26) => Y_SHIFTR_26_port
                           , Y(25) => Y_SHIFTR_25_port, Y(24) => 
                           Y_SHIFTR_24_port, Y(23) => Y_SHIFTR_23_port, Y(22) 
                           => Y_SHIFTR_22_port, Y(21) => Y_SHIFTR_21_port, 
                           Y(20) => Y_SHIFTR_20_port, Y(19) => Y_SHIFTR_19_port
                           , Y(18) => Y_SHIFTR_18_port, Y(17) => 
                           Y_SHIFTR_17_port, Y(16) => Y_SHIFTR_16_port, Y(15) 
                           => Y_SHIFTR_15_port, Y(14) => Y_SHIFTR_14_port, 
                           Y(13) => Y_SHIFTR_13_port, Y(12) => Y_SHIFTR_12_port
                           , Y(11) => Y_SHIFTR_11_port, Y(10) => 
                           Y_SHIFTR_10_port, Y(9) => Y_SHIFTR_9_port, Y(8) => 
                           Y_SHIFTR_8_port, Y(7) => Y_SHIFTR_7_port, Y(6) => 
                           Y_SHIFTR_6_port, Y(5) => Y_SHIFTR_5_port, Y(4) => 
                           Y_SHIFTR_4_port, Y(3) => Y_SHIFTR_3_port, Y(2) => 
                           Y_SHIFTR_2_port, Y(1) => Y_SHIFTR_1_port, Y(0) => 
                           Y_SHIFTR_0_port);
   LOG : LOGIC_N32 port map( A(31) => OP_A_31_port, A(30) => OP_A_30_port, 
                           A(29) => OP_A_29_port, A(28) => OP_A_28_port, A(27) 
                           => OP_A_27_port, A(26) => OP_A_26_port, A(25) => 
                           OP_A_25_port, A(24) => OP_A_24_port, A(23) => 
                           OP_A_23_port, A(22) => OP_A_22_port, A(21) => 
                           OP_A_21_port, A(20) => OP_A_20_port, A(19) => 
                           OP_A_19_port, A(18) => OP_A_18_port, A(17) => 
                           OP_A_17_port, A(16) => OP_A_16_port, A(15) => n245, 
                           A(14) => n244, A(13) => n243, A(12) => n242, A(11) 
                           => n241, A(10) => n240, A(9) => n239, A(8) => n238, 
                           A(7) => n237, A(6) => n236, A(5) => n235, A(4) => 
                           n234, A(3) => n54, A(2) => n53, A(1) => n52, A(0) =>
                           n51, B(31) => OP_B_31_port, B(30) => OP_B_30_port, 
                           B(29) => OP_B_29_port, B(28) => OP_B_28_port, B(27) 
                           => OP_B_27_port, B(26) => OP_B_26_port, B(25) => 
                           OP_B_25_port, B(24) => OP_B_24_port, B(23) => 
                           OP_B_23_port, B(22) => OP_B_22_port, B(21) => 
                           OP_B_21_port, B(20) => OP_B_20_port, B(19) => 
                           OP_B_19_port, B(18) => OP_B_18_port, B(17) => 
                           OP_B_17_port, B(16) => OP_B_16_port, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n50, B(3) => n49, B(2) => n48, 
                           B(1) => n47, B(0) => n46, S(1) => OP_LOGIC_1_port, 
                           S(0) => OP_LOGIC_0_port, Y(31) => Y_LOGIC_31_port, 
                           Y(30) => Y_LOGIC_30_port, Y(29) => Y_LOGIC_29_port, 
                           Y(28) => Y_LOGIC_28_port, Y(27) => Y_LOGIC_27_port, 
                           Y(26) => Y_LOGIC_26_port, Y(25) => Y_LOGIC_25_port, 
                           Y(24) => Y_LOGIC_24_port, Y(23) => Y_LOGIC_23_port, 
                           Y(22) => Y_LOGIC_22_port, Y(21) => Y_LOGIC_21_port, 
                           Y(20) => Y_LOGIC_20_port, Y(19) => Y_LOGIC_19_port, 
                           Y(18) => Y_LOGIC_18_port, Y(17) => Y_LOGIC_17_port, 
                           Y(16) => Y_LOGIC_16_port, Y(15) => Y_LOGIC_15_port, 
                           Y(14) => Y_LOGIC_14_port, Y(13) => Y_LOGIC_13_port, 
                           Y(12) => Y_LOGIC_12_port, Y(11) => Y_LOGIC_11_port, 
                           Y(10) => Y_LOGIC_10_port, Y(9) => Y_LOGIC_9_port, 
                           Y(8) => Y_LOGIC_8_port, Y(7) => Y_LOGIC_7_port, Y(6)
                           => Y_LOGIC_6_port, Y(5) => Y_LOGIC_5_port, Y(4) => 
                           Y_LOGIC_4_port, Y(3) => Y_LOGIC_3_port, Y(2) => 
                           Y_LOGIC_2_port, Y(1) => Y_LOGIC_1_port, Y(0) => 
                           Y_LOGIC_0_port);
   CMP : COMPARATOR_N32 port map( A(31) => OP_A_31_port, A(30) => OP_A_30_port,
                           A(29) => OP_A_29_port, A(28) => OP_A_28_port, A(27) 
                           => OP_A_27_port, A(26) => OP_A_26_port, A(25) => 
                           OP_A_25_port, A(24) => OP_A_24_port, A(23) => 
                           OP_A_23_port, A(22) => OP_A_22_port, A(21) => 
                           OP_A_21_port, A(20) => OP_A_20_port, A(19) => 
                           OP_A_19_port, A(18) => OP_A_18_port, A(17) => 
                           OP_A_17_port, A(16) => OP_A_16_port, A(15) => n245, 
                           A(14) => n244, A(13) => n243, A(12) => n242, A(11) 
                           => n241, A(10) => n240, A(9) => n239, A(8) => n238, 
                           A(7) => n237, A(6) => n236, A(5) => n235, A(4) => 
                           n234, A(3) => n54, A(2) => n53, A(1) => n52, A(0) =>
                           n51, B(31) => OP_B_31_port, B(30) => OP_B_30_port, 
                           B(29) => OP_B_29_port, B(28) => OP_B_28_port, B(27) 
                           => OP_B_27_port, B(26) => OP_B_26_port, B(25) => 
                           OP_B_25_port, B(24) => OP_B_24_port, B(23) => 
                           OP_B_23_port, B(22) => OP_B_22_port, B(21) => 
                           OP_B_21_port, B(20) => OP_B_20_port, B(19) => 
                           OP_B_19_port, B(18) => OP_B_18_port, B(17) => 
                           OP_B_17_port, B(16) => OP_B_16_port, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n50, B(3) => n49, B(2) => n48, 
                           B(1) => n47, B(0) => n46, S(3) => OP_COMPARE_3_port,
                           S(2) => OP_COMPARE_2_port, S(1) => OP_COMPARE_1_port
                           , S(0) => OP_COMPARE_0_port, Y(31) => n_1275, Y(30) 
                           => n_1276, Y(29) => n_1277, Y(28) => n_1278, Y(27) 
                           => n_1279, Y(26) => n_1280, Y(25) => n_1281, Y(24) 
                           => n_1282, Y(23) => n_1283, Y(22) => n_1284, Y(21) 
                           => n_1285, Y(20) => n_1286, Y(19) => n_1287, Y(18) 
                           => n_1288, Y(17) => n_1289, Y(16) => n_1290, Y(15) 
                           => n_1291, Y(14) => n_1292, Y(13) => n_1293, Y(12) 
                           => n_1294, Y(11) => n_1295, Y(10) => n_1296, Y(9) =>
                           n_1297, Y(8) => n_1298, Y(7) => n_1299, Y(6) => 
                           n_1300, Y(5) => n_1301, Y(4) => n_1302, Y(3) => 
                           n_1303, Y(2) => n_1304, Y(1) => n_1305, Y(0) => 
                           Y_COMPARE_0_port);
   ZDET : ZERO_DETECTOR_N32_0 port map( A(31) => Y_31_port, A(30) => Y_30_port,
                           A(29) => Y_29_port, A(28) => Y_28_port, A(27) => 
                           Y_27_port, A(26) => Y_26_port, A(25) => Y_25_port, 
                           A(24) => Y_24_port, A(23) => Y_23_port, A(22) => 
                           Y_22_port, A(21) => Y_21_port, A(20) => Y_20_port, 
                           A(19) => Y_19_port, A(18) => Y_18_port, A(17) => 
                           Y_17_port, A(16) => Y_16_port, A(15) => Y_15_port, 
                           A(14) => Y_14_port, A(13) => Y_13_port, A(12) => 
                           Y_12_port, A(11) => Y_11_port, A(10) => Y_10_port, 
                           A(9) => Y_9_port, A(8) => Y_8_port, A(7) => Y_7_port
                           , A(6) => Y_6_port, A(5) => Y_5_port, A(4) => 
                           Y_4_port, A(3) => Y_3_port, A(2) => Y_2_port, A(1) 
                           => Y_1_port, A(0) => Y_0_port, Y => Z);
   U3 : NOR3_X1 port map( A1 => OPC(5), A2 => OPC(4), A3 => n298, ZN => n191);
   U4 : NOR3_X1 port map( A1 => n298, A2 => OPC(4), A3 => n297, ZN => n213);
   U5 : BUF_X1 port map( A => n45, Z => n42);
   U6 : BUF_X1 port map( A => n45, Z => n43);
   U7 : BUF_X1 port map( A => N281, Z => n31);
   U8 : BUF_X1 port map( A => N246, Z => n45);
   U9 : BUF_X1 port map( A => n1, Z => n34);
   U10 : BUF_X1 port map( A => n62, Z => n15);
   U11 : BUF_X1 port map( A => n59, Z => n27);
   U12 : BUF_X1 port map( A => n60, Z => n23);
   U13 : BUF_X1 port map( A => n202, Z => n8);
   U14 : BUF_X1 port map( A => OP_A_1_port, Z => n52);
   U15 : BUF_X1 port map( A => OP_A_2_port, Z => n53);
   U16 : BUF_X1 port map( A => OP_A_5_port, Z => n235);
   U17 : BUF_X1 port map( A => OP_A_6_port, Z => n236);
   U18 : BUF_X1 port map( A => OP_A_9_port, Z => n239);
   U19 : BUF_X1 port map( A => OP_A_10_port, Z => n240);
   U20 : BUF_X1 port map( A => OP_A_13_port, Z => n243);
   U21 : BUF_X1 port map( A => OP_A_14_port, Z => n244);
   U22 : BUF_X1 port map( A => OP_B_2_port, Z => n48);
   U23 : BUF_X1 port map( A => OP_A_4_port, Z => n234);
   U24 : BUF_X1 port map( A => OP_A_8_port, Z => n238);
   U25 : BUF_X1 port map( A => OP_A_12_port, Z => n242);
   U26 : BUF_X1 port map( A => OP_B_1_port, Z => n47);
   U27 : BUF_X1 port map( A => OP_A_3_port, Z => n54);
   U28 : BUF_X1 port map( A => OP_A_7_port, Z => n237);
   U29 : BUF_X1 port map( A => OP_A_11_port, Z => n241);
   U30 : BUF_X1 port map( A => OP_A_15_port, Z => n245);
   U31 : BUF_X1 port map( A => n61, Z => n19);
   U32 : BUF_X1 port map( A => OP_B_4_port, Z => n50);
   U33 : BUF_X1 port map( A => OP_B_3_port, Z => n49);
   U34 : BUF_X1 port map( A => OP_B_0_port, Z => n46);
   U35 : BUF_X1 port map( A => OP_A_0_port, Z => n51);
   U36 : BUF_X1 port map( A => n42, Z => n40);
   U37 : BUF_X1 port map( A => n42, Z => n39);
   U38 : BUF_X1 port map( A => n43, Z => n38);
   U39 : BUF_X1 port map( A => n43, Z => n37);
   U40 : BUF_X1 port map( A => n43, Z => n36);
   U41 : BUF_X1 port map( A => n42, Z => n41);
   U42 : BUF_X1 port map( A => n31, Z => n28);
   U43 : BUF_X1 port map( A => n279, Z => n5);
   U44 : BUF_X1 port map( A => n279, Z => n6);
   U45 : BUF_X1 port map( A => n31, Z => n29);
   U46 : BUF_X1 port map( A => n278_port, Z => n2);
   U47 : BUF_X1 port map( A => n278_port, Z => n3);
   U48 : INV_X1 port map( A => n34, ZN => n33);
   U49 : INV_X1 port map( A => n34, ZN => n32);
   U50 : BUF_X1 port map( A => n31, Z => n30);
   U51 : BUF_X1 port map( A => n278_port, Z => n4);
   U52 : BUF_X1 port map( A => n279, Z => n7);
   U53 : BUF_X1 port map( A => n44, Z => n35);
   U54 : BUF_X1 port map( A => n45, Z => n44);
   U55 : NOR4_X1 port map( A1 => n14, A2 => n18, A3 => n221, A4 => n28, ZN => 
                           n203);
   U56 : OR2_X1 port map( A1 => N285, A2 => n7, ZN => n221);
   U57 : INV_X1 port map( A => n214, ZN => n280_port);
   U58 : INV_X1 port map( A => n189, ZN => n292);
   U59 : INV_X1 port map( A => n188, ZN => n285_port);
   U60 : NAND4_X1 port map( A1 => n198, A2 => n195, A3 => n196, A4 => n199, ZN 
                           => N287);
   U61 : NAND4_X1 port map( A1 => n194, A2 => n195, A3 => n196, A4 => n197, ZN 
                           => N288);
   U62 : AOI22_X1 port map( A1 => n291, A2 => n285_port, B1 => n218, B2 => 
                           n280_port, ZN => n222);
   U63 : NAND2_X1 port map( A1 => n192, A2 => n193, ZN => N289);
   U64 : NAND2_X1 port map( A1 => n203, A2 => n1, ZN => N246);
   U65 : INV_X1 port map( A => n225, ZN => n279);
   U66 : INV_X1 port map( A => N280, ZN => n278_port);
   U67 : INV_X1 port map( A => n200, ZN => n282);
   U68 : INV_X1 port map( A => n201, ZN => n283);
   U69 : BUF_X1 port map( A => n27, Z => n24);
   U70 : BUF_X1 port map( A => n27, Z => n25);
   U71 : BUF_X1 port map( A => n15, Z => n13);
   U72 : BUF_X1 port map( A => n15, Z => n12);
   U73 : BUF_X1 port map( A => n23, Z => n20);
   U74 : BUF_X1 port map( A => n23, Z => n21);
   U75 : BUF_X1 port map( A => n8, Z => n9);
   U76 : BUF_X1 port map( A => n8, Z => n10);
   U77 : BUF_X1 port map( A => n8, Z => n11);
   U78 : BUF_X1 port map( A => n15, Z => n14);
   U79 : BUF_X1 port map( A => n27, Z => n26);
   U80 : BUF_X1 port map( A => n23, Z => n22);
   U81 : NOR3_X1 port map( A1 => n294, A2 => n298, A3 => n297, ZN => n218);
   U82 : AOI221_X1 port map( B1 => n280_port, B2 => n191, C1 => n288_port, C2 
                           => n213, A => N96, ZN => n225);
   U83 : AOI22_X1 port map( A1 => n223, A2 => n207, B1 => n191, B2 => n220, ZN 
                           => n195);
   U84 : AND2_X1 port map( A1 => n216, A2 => n224, ZN => n223);
   U85 : OAI22_X1 port map( A1 => n226, A2 => n214, B1 => n190, B2 => n293, ZN 
                           => N96);
   U86 : INV_X1 port map( A => n211, ZN => n293);
   U87 : AOI22_X1 port map( A1 => n288_port, A2 => n218, B1 => n211, B2 => n223
                           , ZN => n198);
   U88 : AOI22_X1 port map( A1 => n223, A2 => n218, B1 => n291, B2 => n220, ZN 
                           => n192);
   U89 : AOI22_X1 port map( A1 => n296, A2 => n223, B1 => n292, B2 => n220, ZN 
                           => n194);
   U90 : NAND4_X1 port map( A1 => n194, A2 => n195, A3 => n198, A4 => n227, ZN 
                           => N285);
   U91 : AOI211_X1 port map( C1 => n223, C2 => n291, A => n228, B => N286, ZN 
                           => n227);
   U92 : OAI21_X1 port map( B1 => n190, B2 => n187, A => n192, ZN => n228);
   U93 : AOI22_X1 port map( A1 => n285_port, A2 => n213, B1 => n292, B2 => n223
                           , ZN => n201);
   U94 : AOI22_X1 port map( A1 => n285_port, A2 => n211, B1 => n223, B2 => n191
                           , ZN => n200);
   U95 : INV_X1 port map( A => n226, ZN => n291);
   U96 : NAND2_X1 port map( A1 => n213, A2 => n230, ZN => n193);
   U97 : AOI22_X1 port map( A1 => OP1(0), A2 => n24, B1 => OP2(0), B2 => n20, 
                           ZN => n186);
   U98 : AOI22_X1 port map( A1 => OP1(1), A2 => n24, B1 => OP2(1), B2 => n20, 
                           ZN => n142);
   U99 : AOI22_X1 port map( A1 => OP1(2), A2 => n25, B1 => OP2(2), B2 => n21, 
                           ZN => n98);
   U100 : AOI22_X1 port map( A1 => OP1(3), A2 => n26, B1 => OP2(3), B2 => n22, 
                           ZN => n86);
   U101 : AOI22_X1 port map( A1 => OP1(4), A2 => n26, B1 => OP2(4), B2 => n22, 
                           ZN => n82);
   U102 : AOI22_X1 port map( A1 => OP1(5), A2 => n26, B1 => OP2(5), B2 => n22, 
                           ZN => n78);
   U103 : AOI22_X1 port map( A1 => OP1(6), A2 => n26, B1 => OP2(6), B2 => n22, 
                           ZN => n74);
   U104 : AOI22_X1 port map( A1 => OP1(7), A2 => n26, B1 => OP2(7), B2 => n22, 
                           ZN => n70);
   U105 : AOI22_X1 port map( A1 => OP1(8), A2 => n26, B1 => OP2(8), B2 => n22, 
                           ZN => n66);
   U106 : AOI22_X1 port map( A1 => OP1(9), A2 => n26, B1 => OP2(9), B2 => n22, 
                           ZN => n58);
   U107 : AOI22_X1 port map( A1 => OP1(10), A2 => n24, B1 => OP2(10), B2 => n20
                           , ZN => n182);
   U108 : AOI22_X1 port map( A1 => OP1(11), A2 => n24, B1 => OP2(11), B2 => n20
                           , ZN => n178);
   U109 : AOI22_X1 port map( A1 => OP1(12), A2 => n24, B1 => OP2(12), B2 => n20
                           , ZN => n174);
   U110 : AOI22_X1 port map( A1 => OP1(13), A2 => n24, B1 => OP2(13), B2 => n20
                           , ZN => n170);
   U111 : AOI22_X1 port map( A1 => OP1(14), A2 => n24, B1 => OP2(14), B2 => n20
                           , ZN => n166);
   U112 : AOI22_X1 port map( A1 => OP1(15), A2 => n24, B1 => OP2(15), B2 => n20
                           , ZN => n162);
   U113 : AOI22_X1 port map( A1 => OP1(16), A2 => n24, B1 => OP2(16), B2 => n20
                           , ZN => n158);
   U114 : AOI22_X1 port map( A1 => OP1(17), A2 => n24, B1 => OP2(17), B2 => n20
                           , ZN => n154);
   U115 : AOI22_X1 port map( A1 => OP1(18), A2 => n24, B1 => OP2(18), B2 => n20
                           , ZN => n150);
   U116 : AOI22_X1 port map( A1 => OP1(19), A2 => n24, B1 => OP2(19), B2 => n20
                           , ZN => n146);
   U117 : AOI22_X1 port map( A1 => OP1(20), A2 => n25, B1 => OP2(20), B2 => n21
                           , ZN => n138);
   U118 : AOI22_X1 port map( A1 => OP1(21), A2 => n25, B1 => OP2(21), B2 => n21
                           , ZN => n134);
   U119 : AOI22_X1 port map( A1 => OP1(22), A2 => n25, B1 => OP2(22), B2 => n21
                           , ZN => n130);
   U120 : AOI22_X1 port map( A1 => OP1(23), A2 => n25, B1 => OP2(23), B2 => n21
                           , ZN => n126);
   U121 : AOI22_X1 port map( A1 => OP1(24), A2 => n25, B1 => OP2(24), B2 => n21
                           , ZN => n122);
   U122 : AOI22_X1 port map( A1 => OP1(25), A2 => n25, B1 => OP2(25), B2 => n21
                           , ZN => n118);
   U123 : AOI22_X1 port map( A1 => OP1(26), A2 => n25, B1 => OP2(26), B2 => n21
                           , ZN => n114);
   U124 : AOI22_X1 port map( A1 => OP1(27), A2 => n25, B1 => OP2(27), B2 => n21
                           , ZN => n110);
   U125 : AOI22_X1 port map( A1 => OP1(28), A2 => n25, B1 => OP2(28), B2 => n21
                           , ZN => n106);
   U126 : AOI22_X1 port map( A1 => OP1(29), A2 => n25, B1 => OP2(29), B2 => n21
                           , ZN => n102);
   U127 : AOI22_X1 port map( A1 => OP1(30), A2 => n25, B1 => OP2(30), B2 => n21
                           , ZN => n94);
   U128 : AOI22_X1 port map( A1 => OP1(31), A2 => n26, B1 => OP2(31), B2 => n22
                           , ZN => n90);
   U129 : NAND2_X1 port map( A1 => n191, A2 => n230, ZN => n197);
   U130 : OAI22_X1 port map( A1 => OP2(0), A2 => n2, B1 => n9, B2 => n246_port,
                           ZN => N247);
   U131 : INV_X1 port map( A => OP2(0), ZN => n246_port);
   U132 : OAI22_X1 port map( A1 => OP2(1), A2 => n2, B1 => n9, B2 => n247_port,
                           ZN => N248);
   U133 : INV_X1 port map( A => OP2(1), ZN => n247_port);
   U134 : OAI22_X1 port map( A1 => OP2(2), A2 => n2, B1 => n9, B2 => n248_port,
                           ZN => N249);
   U135 : INV_X1 port map( A => OP2(2), ZN => n248_port);
   U136 : OAI22_X1 port map( A1 => OP2(3), A2 => n2, B1 => n9, B2 => n249_port,
                           ZN => N250);
   U137 : INV_X1 port map( A => OP2(3), ZN => n249_port);
   U138 : OAI22_X1 port map( A1 => OP2(4), A2 => n2, B1 => n9, B2 => n250_port,
                           ZN => N251);
   U139 : INV_X1 port map( A => OP2(4), ZN => n250_port);
   U140 : OAI22_X1 port map( A1 => OP2(5), A2 => n2, B1 => n9, B2 => n251_port,
                           ZN => N252);
   U141 : INV_X1 port map( A => OP2(5), ZN => n251_port);
   U142 : OAI22_X1 port map( A1 => OP2(6), A2 => n2, B1 => n9, B2 => n252_port,
                           ZN => N253);
   U143 : INV_X1 port map( A => OP2(6), ZN => n252_port);
   U144 : OAI22_X1 port map( A1 => OP2(7), A2 => n2, B1 => n9, B2 => n253_port,
                           ZN => N254);
   U145 : INV_X1 port map( A => OP2(7), ZN => n253_port);
   U146 : OAI22_X1 port map( A1 => OP2(8), A2 => n2, B1 => n9, B2 => n254_port,
                           ZN => N255);
   U147 : INV_X1 port map( A => OP2(8), ZN => n254_port);
   U148 : OAI22_X1 port map( A1 => OP2(9), A2 => n2, B1 => n9, B2 => n255_port,
                           ZN => N256);
   U149 : INV_X1 port map( A => OP2(9), ZN => n255_port);
   U150 : OAI22_X1 port map( A1 => OP2(10), A2 => n2, B1 => n9, B2 => n256_port
                           , ZN => N257);
   U151 : INV_X1 port map( A => OP2(10), ZN => n256_port);
   U152 : OAI22_X1 port map( A1 => OP2(11), A2 => n3, B1 => n10, B2 => 
                           n257_port, ZN => N258);
   U153 : INV_X1 port map( A => OP2(11), ZN => n257_port);
   U154 : OAI22_X1 port map( A1 => OP2(12), A2 => n3, B1 => n10, B2 => 
                           n258_port, ZN => N259);
   U155 : INV_X1 port map( A => OP2(12), ZN => n258_port);
   U156 : OAI22_X1 port map( A1 => OP2(13), A2 => n3, B1 => n10, B2 => 
                           n259_port, ZN => N260);
   U157 : INV_X1 port map( A => OP2(13), ZN => n259_port);
   U158 : OAI22_X1 port map( A1 => OP2(14), A2 => n3, B1 => n10, B2 => 
                           n260_port, ZN => N261);
   U159 : INV_X1 port map( A => OP2(14), ZN => n260_port);
   U160 : OAI22_X1 port map( A1 => OP2(15), A2 => n3, B1 => n10, B2 => 
                           n261_port, ZN => N262);
   U161 : INV_X1 port map( A => OP2(15), ZN => n261_port);
   U162 : OAI22_X1 port map( A1 => OP2(16), A2 => n3, B1 => n10, B2 => 
                           n262_port, ZN => N263);
   U163 : INV_X1 port map( A => OP2(16), ZN => n262_port);
   U164 : OAI22_X1 port map( A1 => OP2(17), A2 => n3, B1 => n10, B2 => 
                           n263_port, ZN => N264);
   U165 : INV_X1 port map( A => OP2(17), ZN => n263_port);
   U166 : OAI22_X1 port map( A1 => OP2(18), A2 => n3, B1 => n10, B2 => 
                           n264_port, ZN => N265);
   U167 : INV_X1 port map( A => OP2(18), ZN => n264_port);
   U168 : OAI22_X1 port map( A1 => OP2(19), A2 => n3, B1 => n10, B2 => 
                           n265_port, ZN => N266);
   U169 : INV_X1 port map( A => OP2(19), ZN => n265_port);
   U170 : OAI22_X1 port map( A1 => OP2(20), A2 => n3, B1 => n10, B2 => 
                           n266_port, ZN => N267);
   U171 : INV_X1 port map( A => OP2(20), ZN => n266_port);
   U172 : OAI22_X1 port map( A1 => OP2(21), A2 => n3, B1 => n10, B2 => 
                           n267_port, ZN => N268);
   U173 : INV_X1 port map( A => OP2(21), ZN => n267_port);
   U174 : OAI22_X1 port map( A1 => OP2(22), A2 => n3, B1 => n11, B2 => 
                           n268_port, ZN => N269);
   U175 : INV_X1 port map( A => OP2(22), ZN => n268_port);
   U176 : OAI22_X1 port map( A1 => OP2(23), A2 => n4, B1 => n11, B2 => 
                           n269_port, ZN => N270);
   U177 : INV_X1 port map( A => OP2(23), ZN => n269_port);
   U178 : OAI22_X1 port map( A1 => OP2(24), A2 => n4, B1 => n11, B2 => 
                           n270_port, ZN => N271);
   U179 : INV_X1 port map( A => OP2(24), ZN => n270_port);
   U180 : OAI22_X1 port map( A1 => OP2(25), A2 => n4, B1 => n11, B2 => 
                           n271_port, ZN => N272);
   U181 : INV_X1 port map( A => OP2(25), ZN => n271_port);
   U182 : OAI22_X1 port map( A1 => OP2(26), A2 => n4, B1 => n11, B2 => 
                           n272_port, ZN => N273);
   U183 : INV_X1 port map( A => OP2(26), ZN => n272_port);
   U184 : OAI22_X1 port map( A1 => OP2(27), A2 => n4, B1 => n11, B2 => 
                           n273_port, ZN => N274);
   U185 : INV_X1 port map( A => OP2(27), ZN => n273_port);
   U186 : OAI22_X1 port map( A1 => OP2(28), A2 => n4, B1 => n11, B2 => 
                           n274_port, ZN => N275);
   U187 : INV_X1 port map( A => OP2(28), ZN => n274_port);
   U188 : OAI22_X1 port map( A1 => OP2(29), A2 => n4, B1 => n11, B2 => 
                           n275_port, ZN => N276);
   U189 : INV_X1 port map( A => OP2(29), ZN => n275_port);
   U190 : OAI22_X1 port map( A1 => OP2(30), A2 => n4, B1 => n11, B2 => 
                           n276_port, ZN => N277);
   U191 : INV_X1 port map( A => OP2(30), ZN => n276_port);
   U192 : OAI22_X1 port map( A1 => OP2(31), A2 => n4, B1 => n11, B2 => 
                           n277_port, ZN => N278);
   U193 : INV_X1 port map( A => OP2(31), ZN => n277_port);
   U194 : NAND4_X1 port map( A1 => n183, A2 => n184, A3 => n185, A4 => n186, ZN
                           => Y_0_port);
   U195 : AOI22_X1 port map( A1 => Y_SHIFTR_0_port, A2 => n5, B1 => 
                           Y_COMPARE_0_port, B2 => N285, ZN => n183);
   U196 : AOI22_X1 port map( A1 => Y_SUM_0_port, A2 => n33, B1 => 
                           Y_LOGIC_0_port, B2 => n30, ZN => n184);
   U197 : AOI22_X1 port map( A1 => Y_MUL_0_port, A2 => n18, B1 => 
                           Y_SHIFTL_0_port, B2 => n14, ZN => n185);
   U198 : NAND4_X1 port map( A1 => n139, A2 => n140, A3 => n141, A4 => n142, ZN
                           => Y_1_port);
   U199 : NAND2_X1 port map( A1 => Y_SHIFTR_1_port, A2 => n5, ZN => n139);
   U200 : AOI22_X1 port map( A1 => Y_SUM_1_port, A2 => n33, B1 => 
                           Y_LOGIC_1_port, B2 => n29, ZN => n140);
   U201 : AOI22_X1 port map( A1 => Y_MUL_1_port, A2 => n17, B1 => 
                           Y_SHIFTL_1_port, B2 => n13, ZN => n141);
   U202 : NAND4_X1 port map( A1 => n95, A2 => n96_port, A3 => n97, A4 => n98, 
                           ZN => Y_2_port);
   U203 : NAND2_X1 port map( A1 => Y_SHIFTR_2_port, A2 => n5, ZN => n95);
   U204 : AOI22_X1 port map( A1 => Y_SUM_2_port, A2 => n32, B1 => 
                           Y_LOGIC_2_port, B2 => n28, ZN => n96_port);
   U205 : AOI22_X1 port map( A1 => Y_MUL_2_port, A2 => n16, B1 => 
                           Y_SHIFTL_2_port, B2 => n12, ZN => n97);
   U206 : NAND4_X1 port map( A1 => n83, A2 => n84, A3 => n85, A4 => n86, ZN => 
                           Y_3_port);
   U207 : NAND2_X1 port map( A1 => Y_SHIFTR_3_port, A2 => n5, ZN => n83);
   U208 : AOI22_X1 port map( A1 => Y_SUM_3_port, A2 => n32, B1 => 
                           Y_LOGIC_3_port, B2 => n28, ZN => n84);
   U209 : AOI22_X1 port map( A1 => Y_MUL_3_port, A2 => n16, B1 => 
                           Y_SHIFTL_3_port, B2 => n12, ZN => n85);
   U210 : NAND4_X1 port map( A1 => n79, A2 => n80, A3 => n81, A4 => n82, ZN => 
                           Y_4_port);
   U211 : NAND2_X1 port map( A1 => Y_SHIFTR_4_port, A2 => n5, ZN => n79);
   U212 : AOI22_X1 port map( A1 => Y_SUM_4_port, A2 => n32, B1 => 
                           Y_LOGIC_4_port, B2 => n28, ZN => n80);
   U213 : AOI22_X1 port map( A1 => Y_MUL_4_port, A2 => n16, B1 => 
                           Y_SHIFTL_4_port, B2 => n12, ZN => n81);
   U214 : NAND4_X1 port map( A1 => n75, A2 => n76, A3 => n77, A4 => n78, ZN => 
                           Y_5_port);
   U215 : NAND2_X1 port map( A1 => Y_SHIFTR_5_port, A2 => n5, ZN => n75);
   U216 : AOI22_X1 port map( A1 => Y_SUM_5_port, A2 => n32, B1 => 
                           Y_LOGIC_5_port, B2 => n28, ZN => n76);
   U217 : AOI22_X1 port map( A1 => Y_MUL_5_port, A2 => n16, B1 => 
                           Y_SHIFTL_5_port, B2 => n12, ZN => n77);
   U218 : NAND4_X1 port map( A1 => n71, A2 => n72, A3 => n73, A4 => n74, ZN => 
                           Y_6_port);
   U219 : NAND2_X1 port map( A1 => Y_SHIFTR_6_port, A2 => n5, ZN => n71);
   U220 : AOI22_X1 port map( A1 => Y_SUM_6_port, A2 => n32, B1 => 
                           Y_LOGIC_6_port, B2 => n28, ZN => n72);
   U221 : AOI22_X1 port map( A1 => Y_MUL_6_port, A2 => n16, B1 => 
                           Y_SHIFTL_6_port, B2 => n12, ZN => n73);
   U222 : NAND4_X1 port map( A1 => n67, A2 => n68, A3 => n69, A4 => n70, ZN => 
                           Y_7_port);
   U223 : NAND2_X1 port map( A1 => Y_SHIFTR_7_port, A2 => n6, ZN => n67);
   U224 : AOI22_X1 port map( A1 => Y_SUM_7_port, A2 => n32, B1 => 
                           Y_LOGIC_7_port, B2 => n28, ZN => n68);
   U225 : AOI22_X1 port map( A1 => Y_MUL_7_port, A2 => n16, B1 => 
                           Y_SHIFTL_7_port, B2 => n12, ZN => n69);
   U226 : NAND4_X1 port map( A1 => n63, A2 => n64, A3 => n65, A4 => n66, ZN => 
                           Y_8_port);
   U227 : NAND2_X1 port map( A1 => Y_SHIFTR_8_port, A2 => n5, ZN => n63);
   U228 : AOI22_X1 port map( A1 => Y_SUM_8_port, A2 => n32, B1 => 
                           Y_LOGIC_8_port, B2 => n28, ZN => n64);
   U229 : AOI22_X1 port map( A1 => Y_MUL_8_port, A2 => n16, B1 => 
                           Y_SHIFTL_8_port, B2 => n12, ZN => n65);
   U230 : NAND4_X1 port map( A1 => n55, A2 => n56, A3 => n57, A4 => n58, ZN => 
                           Y_9_port);
   U231 : NAND2_X1 port map( A1 => Y_SHIFTR_9_port, A2 => n5, ZN => n55);
   U232 : AOI22_X1 port map( A1 => Y_SUM_9_port, A2 => n32, B1 => 
                           Y_LOGIC_9_port, B2 => n29, ZN => n56);
   U233 : AOI22_X1 port map( A1 => Y_MUL_9_port, A2 => n16, B1 => 
                           Y_SHIFTL_9_port, B2 => n12, ZN => n57);
   U234 : NAND4_X1 port map( A1 => n179, A2 => n180, A3 => n181, A4 => n182, ZN
                           => Y_10_port);
   U235 : NAND2_X1 port map( A1 => Y_SHIFTR_10_port, A2 => n5, ZN => n179);
   U236 : AOI22_X1 port map( A1 => Y_SUM_10_port, A2 => n32, B1 => 
                           Y_LOGIC_10_port, B2 => n30, ZN => n180);
   U237 : AOI22_X1 port map( A1 => Y_MUL_10_port, A2 => n18, B1 => 
                           Y_SHIFTL_10_port, B2 => n14, ZN => n181);
   U238 : NAND4_X1 port map( A1 => n175, A2 => n176, A3 => n177, A4 => n178, ZN
                           => Y_11_port);
   U239 : NAND2_X1 port map( A1 => Y_SHIFTR_11_port, A2 => n5, ZN => n175);
   U240 : AOI22_X1 port map( A1 => Y_SUM_11_port, A2 => n33, B1 => 
                           Y_LOGIC_11_port, B2 => n30, ZN => n176);
   U241 : AOI22_X1 port map( A1 => Y_MUL_11_port, A2 => n18, B1 => 
                           Y_SHIFTL_11_port, B2 => n14, ZN => n177);
   U242 : NAND4_X1 port map( A1 => n171, A2 => n172, A3 => n173, A4 => n174, ZN
                           => Y_12_port);
   U243 : NAND2_X1 port map( A1 => Y_SHIFTR_12_port, A2 => n6, ZN => n171);
   U244 : AOI22_X1 port map( A1 => Y_SUM_12_port, A2 => n32, B1 => 
                           Y_LOGIC_12_port, B2 => n30, ZN => n172);
   U245 : AOI22_X1 port map( A1 => Y_MUL_12_port, A2 => n18, B1 => 
                           Y_SHIFTL_12_port, B2 => n14, ZN => n173);
   U246 : NAND4_X1 port map( A1 => n167, A2 => n168, A3 => n169, A4 => n170, ZN
                           => Y_13_port);
   U247 : NAND2_X1 port map( A1 => Y_SHIFTR_13_port, A2 => n6, ZN => n167);
   U248 : AOI22_X1 port map( A1 => Y_SUM_13_port, A2 => n33, B1 => 
                           Y_LOGIC_13_port, B2 => n30, ZN => n168);
   U249 : AOI22_X1 port map( A1 => Y_MUL_13_port, A2 => n18, B1 => 
                           Y_SHIFTL_13_port, B2 => n14, ZN => n169);
   U250 : NAND4_X1 port map( A1 => n163, A2 => n164, A3 => n165, A4 => n166, ZN
                           => Y_14_port);
   U251 : NAND2_X1 port map( A1 => Y_SHIFTR_14_port, A2 => n6, ZN => n163);
   U252 : AOI22_X1 port map( A1 => Y_SUM_14_port, A2 => n32, B1 => 
                           Y_LOGIC_14_port, B2 => n30, ZN => n164);
   U253 : AOI22_X1 port map( A1 => Y_MUL_14_port, A2 => n18, B1 => 
                           Y_SHIFTL_14_port, B2 => n14, ZN => n165);
   U254 : NAND4_X1 port map( A1 => n159, A2 => n160, A3 => n161, A4 => n162, ZN
                           => Y_15_port);
   U255 : NAND2_X1 port map( A1 => Y_SHIFTR_15_port, A2 => n6, ZN => n159);
   U256 : AOI22_X1 port map( A1 => Y_SUM_15_port, A2 => n33, B1 => 
                           Y_LOGIC_15_port, B2 => n30, ZN => n160);
   U257 : AOI22_X1 port map( A1 => Y_MUL_15_port, A2 => n18, B1 => 
                           Y_SHIFTL_15_port, B2 => n14, ZN => n161);
   U258 : NAND4_X1 port map( A1 => n155, A2 => n156, A3 => n157, A4 => n158, ZN
                           => Y_16_port);
   U259 : NAND2_X1 port map( A1 => Y_SHIFTR_16_port, A2 => n6, ZN => n155);
   U260 : AOI22_X1 port map( A1 => Y_SUM_16_port, A2 => n32, B1 => 
                           Y_LOGIC_16_port, B2 => n30, ZN => n156);
   U261 : AOI22_X1 port map( A1 => Y_MUL_16_port, A2 => n18, B1 => 
                           Y_SHIFTL_16_port, B2 => n14, ZN => n157);
   U262 : NAND4_X1 port map( A1 => n151, A2 => n152, A3 => n153, A4 => n154, ZN
                           => Y_17_port);
   U263 : NAND2_X1 port map( A1 => Y_SHIFTR_17_port, A2 => n6, ZN => n151);
   U264 : AOI22_X1 port map( A1 => Y_SUM_17_port, A2 => n33, B1 => 
                           Y_LOGIC_17_port, B2 => n30, ZN => n152);
   U265 : AOI22_X1 port map( A1 => Y_MUL_17_port, A2 => n17, B1 => 
                           Y_SHIFTL_17_port, B2 => n13, ZN => n153);
   U266 : NAND4_X1 port map( A1 => n147, A2 => n148, A3 => n149, A4 => n150, ZN
                           => Y_18_port);
   U267 : NAND2_X1 port map( A1 => Y_SHIFTR_18_port, A2 => n6, ZN => n147);
   U268 : AOI22_X1 port map( A1 => Y_SUM_18_port, A2 => n33, B1 => 
                           Y_LOGIC_18_port, B2 => n29, ZN => n148);
   U269 : AOI22_X1 port map( A1 => Y_MUL_18_port, A2 => n17, B1 => 
                           Y_SHIFTL_18_port, B2 => n13, ZN => n149);
   U270 : NAND4_X1 port map( A1 => n143, A2 => n144, A3 => n145, A4 => n146, ZN
                           => Y_19_port);
   U271 : NAND2_X1 port map( A1 => Y_SHIFTR_19_port, A2 => n6, ZN => n143);
   U272 : AOI22_X1 port map( A1 => Y_SUM_19_port, A2 => n33, B1 => 
                           Y_LOGIC_19_port, B2 => n29, ZN => n144);
   U273 : AOI22_X1 port map( A1 => Y_MUL_19_port, A2 => n17, B1 => 
                           Y_SHIFTL_19_port, B2 => n13, ZN => n145);
   U274 : NAND4_X1 port map( A1 => n135, A2 => n136, A3 => n137, A4 => n138, ZN
                           => Y_20_port);
   U275 : NAND2_X1 port map( A1 => Y_SHIFTR_20_port, A2 => n6, ZN => n135);
   U276 : AOI22_X1 port map( A1 => Y_SUM_20_port, A2 => n33, B1 => 
                           Y_LOGIC_20_port, B2 => n29, ZN => n136);
   U277 : AOI22_X1 port map( A1 => Y_MUL_20_port, A2 => n17, B1 => 
                           Y_SHIFTL_20_port, B2 => n13, ZN => n137);
   U278 : NAND4_X1 port map( A1 => n131, A2 => n132, A3 => n133, A4 => n134, ZN
                           => Y_21_port);
   U279 : NAND2_X1 port map( A1 => Y_SHIFTR_21_port, A2 => n6, ZN => n131);
   U280 : AOI22_X1 port map( A1 => Y_SUM_21_port, A2 => n33, B1 => 
                           Y_LOGIC_21_port, B2 => n29, ZN => n132);
   U281 : AOI22_X1 port map( A1 => Y_MUL_21_port, A2 => n17, B1 => 
                           Y_SHIFTL_21_port, B2 => n13, ZN => n133);
   U282 : NAND4_X1 port map( A1 => n127, A2 => n128, A3 => n129, A4 => n130, ZN
                           => Y_22_port);
   U283 : NAND2_X1 port map( A1 => Y_SHIFTR_22_port, A2 => n6, ZN => n127);
   U284 : AOI22_X1 port map( A1 => Y_SUM_22_port, A2 => n33, B1 => 
                           Y_LOGIC_22_port, B2 => n29, ZN => n128);
   U285 : AOI22_X1 port map( A1 => Y_MUL_22_port, A2 => n17, B1 => 
                           Y_SHIFTL_22_port, B2 => n13, ZN => n129);
   U286 : NAND4_X1 port map( A1 => n123, A2 => n124, A3 => n125, A4 => n126, ZN
                           => Y_23_port);
   U287 : NAND2_X1 port map( A1 => Y_SHIFTR_23_port, A2 => n7, ZN => n123);
   U288 : AOI22_X1 port map( A1 => Y_SUM_23_port, A2 => n33, B1 => 
                           Y_LOGIC_23_port, B2 => n29, ZN => n124);
   U289 : AOI22_X1 port map( A1 => Y_MUL_23_port, A2 => n17, B1 => 
                           Y_SHIFTL_23_port, B2 => n13, ZN => n125);
   U290 : NAND4_X1 port map( A1 => n119, A2 => n120, A3 => n121, A4 => n122, ZN
                           => Y_24_port);
   U291 : NAND2_X1 port map( A1 => Y_SHIFTR_24_port, A2 => n7, ZN => n119);
   U292 : AOI22_X1 port map( A1 => Y_SUM_24_port, A2 => n33, B1 => 
                           Y_LOGIC_24_port, B2 => n29, ZN => n120);
   U293 : AOI22_X1 port map( A1 => Y_MUL_24_port, A2 => n17, B1 => 
                           Y_SHIFTL_24_port, B2 => n13, ZN => n121);
   U294 : NAND4_X1 port map( A1 => n115, A2 => n116, A3 => n117, A4 => n118, ZN
                           => Y_25_port);
   U295 : NAND2_X1 port map( A1 => Y_SHIFTR_25_port, A2 => n7, ZN => n115);
   U296 : AOI22_X1 port map( A1 => Y_SUM_25_port, A2 => n33, B1 => 
                           Y_LOGIC_25_port, B2 => n29, ZN => n116);
   U297 : AOI22_X1 port map( A1 => Y_MUL_25_port, A2 => n17, B1 => 
                           Y_SHIFTL_25_port, B2 => n13, ZN => n117);
   U298 : NAND4_X1 port map( A1 => n111, A2 => n112, A3 => n113, A4 => n114, ZN
                           => Y_26_port);
   U299 : NAND2_X1 port map( A1 => Y_SHIFTR_26_port, A2 => n7, ZN => n111);
   U300 : AOI22_X1 port map( A1 => Y_SUM_26_port, A2 => n33, B1 => 
                           Y_LOGIC_26_port, B2 => n29, ZN => n112);
   U310 : AOI22_X1 port map( A1 => Y_MUL_26_port, A2 => n17, B1 => 
                           Y_SHIFTL_26_port, B2 => n13, ZN => n113);
   U311 : NAND4_X1 port map( A1 => n107, A2 => n108, A3 => n109, A4 => n110, ZN
                           => Y_27_port);
   U312 : NAND2_X1 port map( A1 => Y_SHIFTR_27_port, A2 => n7, ZN => n107);
   U313 : AOI22_X1 port map( A1 => Y_SUM_27_port, A2 => n33, B1 => 
                           Y_LOGIC_27_port, B2 => n29, ZN => n108);
   U314 : AOI22_X1 port map( A1 => Y_MUL_27_port, A2 => n17, B1 => 
                           Y_SHIFTL_27_port, B2 => n13, ZN => n109);
   U315 : NAND4_X1 port map( A1 => n103, A2 => n104, A3 => n105, A4 => n106, ZN
                           => Y_28_port);
   U316 : NAND2_X1 port map( A1 => Y_SHIFTR_28_port, A2 => n7, ZN => n103);
   U317 : AOI22_X1 port map( A1 => Y_SUM_28_port, A2 => n32, B1 => 
                           Y_LOGIC_28_port, B2 => n28, ZN => n104);
   U318 : AOI22_X1 port map( A1 => Y_MUL_28_port, A2 => n16, B1 => 
                           Y_SHIFTL_28_port, B2 => n12, ZN => n105);
   U319 : NAND4_X1 port map( A1 => n99, A2 => n100, A3 => n101, A4 => n102, ZN 
                           => Y_29_port);
   U320 : NAND2_X1 port map( A1 => Y_SHIFTR_29_port, A2 => n7, ZN => n99);
   U321 : AOI22_X1 port map( A1 => Y_SUM_29_port, A2 => n32, B1 => 
                           Y_LOGIC_29_port, B2 => n28, ZN => n100);
   U322 : AOI22_X1 port map( A1 => Y_MUL_29_port, A2 => n16, B1 => 
                           Y_SHIFTL_29_port, B2 => n12, ZN => n101);
   U323 : NAND4_X1 port map( A1 => n91, A2 => n92, A3 => n93, A4 => n94, ZN => 
                           Y_30_port);
   U324 : NAND2_X1 port map( A1 => Y_SHIFTR_30_port, A2 => n7, ZN => n91);
   U325 : AOI22_X1 port map( A1 => Y_SUM_30_port, A2 => n32, B1 => 
                           Y_LOGIC_30_port, B2 => n28, ZN => n92);
   U326 : AOI22_X1 port map( A1 => Y_MUL_30_port, A2 => n16, B1 => 
                           Y_SHIFTL_30_port, B2 => n12, ZN => n93);
   U327 : NAND4_X1 port map( A1 => n87, A2 => n88, A3 => n89, A4 => n90, ZN => 
                           Y_31_port);
   U328 : NAND2_X1 port map( A1 => Y_SHIFTR_31_port, A2 => n5, ZN => n87);
   U329 : AOI22_X1 port map( A1 => Y_SUM_31_port, A2 => n32, B1 => 
                           Y_LOGIC_31_port, B2 => n28, ZN => n88);
   U330 : AOI22_X1 port map( A1 => Y_MUL_31_port, A2 => n16, B1 => 
                           Y_SHIFTL_31_port, B2 => n12, ZN => n89);
   U331 : INV_X1 port map( A => n190, ZN => n288_port);
   U332 : NAND4_X1 port map( A1 => n197, A2 => n199, A3 => n196, A4 => n229, ZN
                           => N286);
   U333 : AOI221_X1 port map( B1 => n207, B2 => n288_port, C1 => n223, C2 => 
                           n213, A => n284, ZN => n229);
   U334 : INV_X1 port map( A => n193, ZN => n284);
   U335 : NAND2_X1 port map( A1 => n291, A2 => n230, ZN => n196);
   U336 : INV_X1 port map( A => n187, ZN => n296);
   U337 : OR4_X1 port map( A1 => n218, A2 => n291, A3 => n207, A4 => n213, ZN 
                           => n217);
   U338 : NAND2_X1 port map( A1 => n292, A2 => n230, ZN => n199);
   U339 : AND2_X1 port map( A1 => n204, A2 => n2, ZN => n1);
   U340 : NAND2_X1 port map( A1 => n286_port, A2 => n224, ZN => n188);
   U341 : NAND2_X1 port map( A1 => n205, A2 => n206, ZN => N280);
   U342 : OAI21_X1 port map( B1 => n296, B2 => n207, A => n280_port, ZN => n205
                           );
   U343 : OAI21_X1 port map( B1 => n191, B2 => n292, A => n285_port, ZN => n206
                           );
   U344 : OAI22_X1 port map( A1 => n190, A2 => n226, B1 => n214, B2 => n189, ZN
                           => n62);
   U345 : INV_X1 port map( A => n219, ZN => n287_port);
   U346 : AOI21_X1 port map( B1 => n295, B2 => n189, A => n190, ZN => n59);
   U347 : INV_X1 port map( A => n191, ZN => n295);
   U348 : NOR2_X1 port map( A1 => n187, A2 => n188, ZN => n60);
   U349 : INV_X1 port map( A => n232, ZN => n286_port);
   U350 : AND2_X1 port map( A1 => n203, A2 => n204, ZN => n202);
   U351 : BUF_X1 port map( A => n19, Z => n17);
   U352 : BUF_X1 port map( A => n19, Z => n16);
   U353 : BUF_X1 port map( A => n19, Z => n18);
   U354 : NOR3_X1 port map( A1 => n294, A2 => OPC(6), A3 => n297, ZN => n207);
   U355 : NOR3_X1 port map( A1 => OPC(6), A2 => OPC(5), A3 => n294, ZN => n211)
                           ;
   U356 : NOR3_X1 port map( A1 => n232, A2 => OPC(2), A3 => n289_port, ZN => 
                           n219);
   U357 : NOR2_X1 port map( A1 => OPC(1), A2 => OPC(2), ZN => n224);
   U358 : NOR2_X1 port map( A1 => n290, A2 => OPC(0), ZN => n216);
   U359 : NAND2_X1 port map( A1 => n287_port, A2 => n231, ZN => n230);
   U360 : AND3_X1 port map( A1 => n286_port, A2 => n289_port, A3 => OPC(2), ZN 
                           => n220);
   U361 : INV_X1 port map( A => OPC(5), ZN => n297);
   U362 : INV_X1 port map( A => OPC(6), ZN => n298);
   U363 : INV_X1 port map( A => OPC(4), ZN => n294);
   U364 : NAND4_X1 port map( A1 => OPC(2), A2 => OPC(0), A3 => OPC(3), A4 => 
                           n289_port, ZN => n215);
   U365 : INV_X1 port map( A => OPC(1), ZN => n289_port);
   U366 : NAND2_X1 port map( A1 => OPC(0), A2 => n290, ZN => n232);
   U367 : INV_X1 port map( A => OPC(3), ZN => n290);
   U368 : AND3_X1 port map( A1 => n208, A2 => n209, A3 => n210, ZN => n204);
   U369 : OAI21_X1 port map( B1 => n219, B2 => n220, A => n296, ZN => n208);
   U370 : NAND4_X1 port map( A1 => n216, A2 => OPC(1), A3 => OPC(2), A4 => n217
                           , ZN => n209);
   U371 : AOI22_X1 port map( A1 => n211, A2 => n212, B1 => n213, B2 => 
                           n280_port, ZN => n210);
   U372 : INV_X1 port map( A => OPC(0), ZN => n281_port);
   U373 : AND4_X1 port map( A1 => OPC(1), A2 => n291, A3 => n233, A4 => 
                           n281_port, ZN => n61);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX41_N32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX41_N32_1;

architecture SYN_BEHAVIORAL of MUX41_N32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n6, Z => n76);
   U2 : BUF_X1 port map( A => n7, Z => n72);
   U3 : BUF_X1 port map( A => n4, Z => n81);
   U4 : BUF_X1 port map( A => n5, Z => n77);
   U5 : INV_X1 port map( A => S(0), ZN => n85);
   U6 : BUF_X1 port map( A => n76, Z => n73);
   U7 : BUF_X1 port map( A => n76, Z => n74);
   U8 : BUF_X1 port map( A => n81, Z => n82);
   U9 : BUF_X1 port map( A => n81, Z => n83);
   U10 : BUF_X1 port map( A => n72, Z => n1);
   U11 : BUF_X1 port map( A => n72, Z => n70);
   U12 : BUF_X1 port map( A => n77, Z => n78);
   U13 : BUF_X1 port map( A => n77, Z => n79);
   U14 : BUF_X1 port map( A => n76, Z => n75);
   U15 : BUF_X1 port map( A => n81, Z => n84);
   U16 : BUF_X1 port map( A => n72, Z => n71);
   U17 : BUF_X1 port map( A => n77, Z => n80);
   U18 : NOR2_X1 port map( A1 => n85, A2 => S(1), ZN => n6);
   U19 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n7);
   U20 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n4);
   U21 : AND2_X1 port map( A1 => S(1), A2 => n85, ZN => n5);
   U22 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Y(0));
   U23 : AOI22_X1 port map( A1 => D(0), A2 => n82, B1 => C(0), B2 => n78, ZN =>
                           n69);
   U24 : AOI22_X1 port map( A1 => B(0), A2 => n73, B1 => A(0), B2 => n1, ZN => 
                           n68);
   U25 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Y(1));
   U26 : AOI22_X1 port map( A1 => D(1), A2 => n82, B1 => C(1), B2 => n78, ZN =>
                           n47);
   U27 : AOI22_X1 port map( A1 => B(1), A2 => n73, B1 => A(1), B2 => n1, ZN => 
                           n46);
   U28 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(2));
   U29 : AOI22_X1 port map( A1 => D(2), A2 => n83, B1 => C(2), B2 => n79, ZN =>
                           n25);
   U30 : AOI22_X1 port map( A1 => B(2), A2 => n74, B1 => A(2), B2 => n70, ZN =>
                           n24);
   U31 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(3));
   U32 : AOI22_X1 port map( A1 => D(3), A2 => n84, B1 => C(3), B2 => n80, ZN =>
                           n19);
   U33 : AOI22_X1 port map( A1 => B(3), A2 => n75, B1 => A(3), B2 => n71, ZN =>
                           n18);
   U34 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(4));
   U35 : AOI22_X1 port map( A1 => D(4), A2 => n84, B1 => C(4), B2 => n80, ZN =>
                           n17);
   U36 : AOI22_X1 port map( A1 => B(4), A2 => n75, B1 => A(4), B2 => n71, ZN =>
                           n16);
   U37 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(5));
   U38 : AOI22_X1 port map( A1 => D(5), A2 => n84, B1 => C(5), B2 => n80, ZN =>
                           n15);
   U39 : AOI22_X1 port map( A1 => B(5), A2 => n75, B1 => A(5), B2 => n71, ZN =>
                           n14);
   U40 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Y(6));
   U41 : AOI22_X1 port map( A1 => D(6), A2 => n84, B1 => C(6), B2 => n80, ZN =>
                           n13);
   U42 : AOI22_X1 port map( A1 => B(6), A2 => n75, B1 => A(6), B2 => n71, ZN =>
                           n12);
   U43 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Y(7));
   U44 : AOI22_X1 port map( A1 => D(7), A2 => n84, B1 => C(7), B2 => n80, ZN =>
                           n11);
   U45 : AOI22_X1 port map( A1 => B(7), A2 => n75, B1 => A(7), B2 => n71, ZN =>
                           n10);
   U46 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Y(8));
   U47 : AOI22_X1 port map( A1 => D(8), A2 => n84, B1 => C(8), B2 => n80, ZN =>
                           n9);
   U48 : AOI22_X1 port map( A1 => B(8), A2 => n75, B1 => A(8), B2 => n71, ZN =>
                           n8);
   U49 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Y(9));
   U50 : AOI22_X1 port map( A1 => D(9), A2 => n84, B1 => C(9), B2 => n80, ZN =>
                           n3);
   U51 : AOI22_X1 port map( A1 => B(9), A2 => n75, B1 => A(9), B2 => n71, ZN =>
                           n2);
   U52 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Y(10));
   U53 : AOI22_X1 port map( A1 => D(10), A2 => n82, B1 => C(10), B2 => n78, ZN 
                           => n67);
   U54 : AOI22_X1 port map( A1 => B(10), A2 => n73, B1 => A(10), B2 => n1, ZN 
                           => n66);
   U55 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Y(11));
   U56 : AOI22_X1 port map( A1 => D(11), A2 => n82, B1 => C(11), B2 => n78, ZN 
                           => n65);
   U57 : AOI22_X1 port map( A1 => B(11), A2 => n73, B1 => A(11), B2 => n1, ZN 
                           => n64);
   U58 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Y(12));
   U59 : AOI22_X1 port map( A1 => D(12), A2 => n82, B1 => C(12), B2 => n78, ZN 
                           => n63);
   U60 : AOI22_X1 port map( A1 => B(12), A2 => n73, B1 => A(12), B2 => n1, ZN 
                           => n62);
   U61 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Y(13));
   U62 : AOI22_X1 port map( A1 => D(13), A2 => n82, B1 => C(13), B2 => n78, ZN 
                           => n61);
   U63 : AOI22_X1 port map( A1 => B(13), A2 => n73, B1 => A(13), B2 => n1, ZN 
                           => n60);
   U64 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Y(14));
   U65 : AOI22_X1 port map( A1 => D(14), A2 => n82, B1 => C(14), B2 => n78, ZN 
                           => n59);
   U66 : AOI22_X1 port map( A1 => B(14), A2 => n73, B1 => A(14), B2 => n1, ZN 
                           => n58);
   U67 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Y(15));
   U68 : AOI22_X1 port map( A1 => D(15), A2 => n82, B1 => C(15), B2 => n78, ZN 
                           => n57);
   U69 : AOI22_X1 port map( A1 => B(15), A2 => n73, B1 => A(15), B2 => n1, ZN 
                           => n56);
   U70 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Y(16));
   U71 : AOI22_X1 port map( A1 => D(16), A2 => n82, B1 => C(16), B2 => n78, ZN 
                           => n55);
   U72 : AOI22_X1 port map( A1 => B(16), A2 => n73, B1 => A(16), B2 => n1, ZN 
                           => n54);
   U73 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Y(17));
   U74 : AOI22_X1 port map( A1 => D(17), A2 => n82, B1 => C(17), B2 => n78, ZN 
                           => n53);
   U75 : AOI22_X1 port map( A1 => B(17), A2 => n73, B1 => A(17), B2 => n1, ZN 
                           => n52);
   U76 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Y(18));
   U77 : AOI22_X1 port map( A1 => D(18), A2 => n82, B1 => C(18), B2 => n78, ZN 
                           => n51);
   U78 : AOI22_X1 port map( A1 => B(18), A2 => n73, B1 => A(18), B2 => n1, ZN 
                           => n50);
   U79 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Y(19));
   U80 : AOI22_X1 port map( A1 => D(19), A2 => n82, B1 => C(19), B2 => n78, ZN 
                           => n49);
   U81 : AOI22_X1 port map( A1 => B(19), A2 => n73, B1 => A(19), B2 => n1, ZN 
                           => n48);
   U82 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Y(20));
   U83 : AOI22_X1 port map( A1 => D(20), A2 => n83, B1 => C(20), B2 => n79, ZN 
                           => n45);
   U84 : AOI22_X1 port map( A1 => B(20), A2 => n74, B1 => A(20), B2 => n70, ZN 
                           => n44);
   U85 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Y(21));
   U86 : AOI22_X1 port map( A1 => D(21), A2 => n83, B1 => C(21), B2 => n79, ZN 
                           => n43);
   U87 : AOI22_X1 port map( A1 => B(21), A2 => n74, B1 => A(21), B2 => n70, ZN 
                           => n42);
   U88 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Y(22));
   U89 : AOI22_X1 port map( A1 => D(22), A2 => n83, B1 => C(22), B2 => n79, ZN 
                           => n41);
   U90 : AOI22_X1 port map( A1 => B(22), A2 => n74, B1 => A(22), B2 => n70, ZN 
                           => n40);
   U91 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Y(23));
   U92 : AOI22_X1 port map( A1 => D(23), A2 => n83, B1 => C(23), B2 => n79, ZN 
                           => n39);
   U93 : AOI22_X1 port map( A1 => B(23), A2 => n74, B1 => A(23), B2 => n70, ZN 
                           => n38);
   U94 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Y(24));
   U95 : AOI22_X1 port map( A1 => D(24), A2 => n83, B1 => C(24), B2 => n79, ZN 
                           => n37);
   U96 : AOI22_X1 port map( A1 => B(24), A2 => n74, B1 => A(24), B2 => n70, ZN 
                           => n36);
   U97 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Y(25));
   U98 : AOI22_X1 port map( A1 => D(25), A2 => n83, B1 => C(25), B2 => n79, ZN 
                           => n35);
   U99 : AOI22_X1 port map( A1 => B(25), A2 => n74, B1 => A(25), B2 => n70, ZN 
                           => n34);
   U100 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Y(26));
   U101 : AOI22_X1 port map( A1 => D(26), A2 => n83, B1 => C(26), B2 => n79, ZN
                           => n33);
   U102 : AOI22_X1 port map( A1 => B(26), A2 => n74, B1 => A(26), B2 => n70, ZN
                           => n32);
   U103 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(27));
   U104 : AOI22_X1 port map( A1 => D(27), A2 => n83, B1 => C(27), B2 => n79, ZN
                           => n31);
   U105 : AOI22_X1 port map( A1 => B(27), A2 => n74, B1 => A(27), B2 => n70, ZN
                           => n30);
   U106 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Y(28));
   U107 : AOI22_X1 port map( A1 => D(28), A2 => n83, B1 => C(28), B2 => n79, ZN
                           => n29);
   U108 : AOI22_X1 port map( A1 => B(28), A2 => n74, B1 => A(28), B2 => n70, ZN
                           => n28);
   U109 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Y(29));
   U110 : AOI22_X1 port map( A1 => D(29), A2 => n83, B1 => C(29), B2 => n79, ZN
                           => n27);
   U111 : AOI22_X1 port map( A1 => B(29), A2 => n74, B1 => A(29), B2 => n70, ZN
                           => n26);
   U112 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Y(30));
   U113 : AOI22_X1 port map( A1 => D(30), A2 => n83, B1 => C(30), B2 => n79, ZN
                           => n23);
   U114 : AOI22_X1 port map( A1 => B(30), A2 => n74, B1 => A(30), B2 => n70, ZN
                           => n22);
   U115 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Y(31));
   U116 : AOI22_X1 port map( A1 => D(31), A2 => n84, B1 => C(31), B2 => n80, ZN
                           => n21);
   U117 : AOI22_X1 port map( A1 => B(31), A2 => n75, B1 => A(31), B2 => n71, ZN
                           => n20);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REGADDR_N32_OPC6_REG5 is

   port( INSTR : in std_logic_vector (31 downto 0);  RS1, RS2, RD : out 
         std_logic_vector (4 downto 0));

end REGADDR_N32_OPC6_REG5;

architecture SYN_BEHAVIORAL of REGADDR_N32_OPC6_REG5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n16, n23, n24, n25, n26, n27, net24608, net24609, net24616, net31033,
      net39258, net39347, net39721, net39703, net39746, net39757, net40157, 
      net40115, net40113, net40102, n29, net40276, net40137, net40133, net40127
      , net40125, net40107, net40103, net40098, net40092, net40080, net39686, 
      net39315, net24613, net39750, net39747, net39726, net39724, net39618, 
      net39298, net39249, net38954, net24619, net24618, net24614, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14 : std_logic;

begin
   
   U46 : NAND3_X1 port map( A1 => n27, A2 => n24, A3 => n26, ZN => n23);
   U3 : NAND2_X1 port map( A1 => net40103, A2 => n8, ZN => n1);
   U4 : CLKBUF_X1 port map( A => INSTR(26), Z => net40115);
   U5 : OR3_X2 port map( A1 => net39721, A2 => n6, A3 => net40127, ZN => 
                           net40103);
   U6 : OR2_X1 port map( A1 => INSTR(29), A2 => INSTR(31), ZN => net39315);
   U7 : BUF_X1 port map( A => net24619, Z => net39618);
   U8 : AND2_X1 port map( A1 => net40157, A2 => net39703, ZN => net39746);
   U9 : NAND4_X1 port map( A1 => net40133, A2 => net40276, A3 => n29, A4 => 
                           net31033, ZN => n2);
   U10 : NAND2_X1 port map( A1 => net39746, A2 => net39618, ZN => n3);
   U11 : AND2_X1 port map( A1 => INSTR(21), A2 => n3, ZN => RS1(0));
   U12 : CLKBUF_X1 port map( A => INSTR(26), Z => n4);
   U13 : BUF_X1 port map( A => INSTR(28), Z => n5);
   U14 : NAND2_X1 port map( A1 => net40080, A2 => INSTR(29), ZN => net40107);
   U15 : NAND4_X1 port map( A1 => net39258, A2 => net24616, A3 => net24619, A4 
                           => net39721, ZN => n24);
   U16 : INV_X1 port map( A => n4, ZN => n6);
   U17 : AND2_X1 port map( A1 => net39726, A2 => net39747, ZN => RS2(3));
   U18 : AND2_X1 port map( A1 => n7, A2 => INSTR(19), ZN => net39747);
   U19 : INV_X1 port map( A => INSTR(19), ZN => net24614);
   U20 : OAI221_X1 port map( B1 => net24614, B2 => net39757, C1 => net39347, C2
                           => net24609, A => n25, ZN => RD(3));
   U21 : AND2_X1 port map( A1 => net40092, A2 => net39686, ZN => net39726);
   U22 : AND2_X1 port map( A1 => net39726, A2 => net39750, ZN => RS2(2));
   U23 : AND2_X1 port map( A1 => net24618, A2 => net39618, ZN => n7);
   U24 : AND2_X1 port map( A1 => n7, A2 => INSTR(18), ZN => net39750);
   U25 : AND2_X1 port map( A1 => net39618, A2 => net24618, ZN => net38954);
   U26 : INV_X1 port map( A => INSTR(30), ZN => net24619);
   U27 : AND3_X1 port map( A1 => net40113, A2 => net24619, A3 => net39298, ZN 
                           => n29);
   U28 : INV_X1 port map( A => net39249, ZN => net24618);
   U29 : INV_X1 port map( A => net39298, ZN => net39249);
   U30 : INV_X1 port map( A => INSTR(28), ZN => net39298);
   U31 : NAND2_X1 port map( A1 => n1, A2 => net39724, ZN => n16);
   U32 : AND2_X1 port map( A1 => net38954, A2 => net39686, ZN => net39724);
   U33 : NOR2_X1 port map( A1 => net39315, A2 => n5, ZN => net40157);
   U34 : NOR2_X1 port map( A1 => net39315, A2 => n5, ZN => net39258);
   U35 : INV_X1 port map( A => INSTR(18), ZN => net24613);
   U36 : OAI221_X1 port map( B1 => n23, B2 => net24613, C1 => net39347, C2 => 
                           net24608, A => n25, ZN => RD(2));
   U37 : NAND2_X1 port map( A1 => net40103, A2 => n8, ZN => net40092);
   U38 : MUX2_X1 port map( A => net40107, B => net39315, S => net40098, Z => n8
                           );
   U39 : BUF_X1 port map( A => net40080, Z => net40125);
   U40 : INV_X1 port map( A => net40125, ZN => net40133);
   U41 : NAND2_X1 port map( A1 => net40125, A2 => net40137, ZN => net39686);
   U42 : INV_X1 port map( A => INSTR(31), ZN => net40080);
   U43 : INV_X1 port map( A => net40127, ZN => net40276);
   U44 : NAND4_X1 port map( A1 => net40133, A2 => net40276, A3 => n29, A4 => 
                           net31033, ZN => n27);
   U45 : INV_X1 port map( A => INSTR(29), ZN => net40127);
   U47 : OAI21_X1 port map( B1 => net40127, B2 => net40098, A => net40102, ZN 
                           => net40137);
   U48 : BUF_X1 port map( A => INSTR(27), Z => net40113);
   U49 : XNOR2_X1 port map( A => INSTR(26), B => INSTR(27), ZN => net40098);
   U50 : NAND2_X1 port map( A1 => net40113, A2 => net40115, ZN => net40102);
   U51 : INV_X1 port map( A => net40115, ZN => net24616);
   U52 : INV_X1 port map( A => net40113, ZN => net39721);
   U53 : INV_X1 port map( A => net24616, ZN => net31033);
   U54 : NAND3_X1 port map( A1 => n2, A2 => n24, A3 => n26, ZN => net39757);
   U55 : NAND2_X1 port map( A1 => net40157, A2 => net39703, ZN => n26);
   U56 : INV_X1 port map( A => net39721, ZN => net39703);
   U57 : BUF_X1 port map( A => n24, Z => net39347);
   U58 : INV_X1 port map( A => INSTR(11), ZN => n14);
   U59 : INV_X1 port map( A => INSTR(12), ZN => n13);
   U60 : INV_X1 port map( A => INSTR(13), ZN => net24608);
   U61 : INV_X1 port map( A => INSTR(14), ZN => net24609);
   U62 : INV_X1 port map( A => INSTR(15), ZN => n12);
   U63 : AND2_X1 port map( A1 => INSTR(25), A2 => n3, ZN => RS1(4));
   U64 : AND2_X1 port map( A1 => INSTR(23), A2 => n3, ZN => RS1(2));
   U65 : AND2_X1 port map( A1 => INSTR(22), A2 => n3, ZN => RS1(1));
   U66 : AND2_X1 port map( A1 => INSTR(24), A2 => n3, ZN => RS1(3));
   U67 : INV_X1 port map( A => INSTR(17), ZN => n10);
   U68 : INV_X1 port map( A => INSTR(16), ZN => n11);
   U69 : INV_X1 port map( A => INSTR(20), ZN => n9);
   U70 : OAI221_X1 port map( B1 => n23, B2 => n9, C1 => net39347, C2 => n12, A 
                           => n25, ZN => RD(4));
   U71 : OAI221_X1 port map( B1 => n10, B2 => net39757, C1 => net39347, C2 => 
                           n13, A => n25, ZN => RD(1));
   U72 : OAI221_X1 port map( B1 => n23, B2 => n11, C1 => net39347, C2 => n14, A
                           => n25, ZN => RD(0));
   U73 : NOR2_X1 port map( A1 => n16, A2 => n11, ZN => RS2(0));
   U74 : NOR2_X1 port map( A1 => n16, A2 => n10, ZN => RS2(1));
   U75 : NOR2_X1 port map( A1 => n16, A2 => n9, ZN => RS2(4));
   U76 : NAND2_X1 port map( A1 => net39746, A2 => net31033, ZN => n25);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SIGNEX_N32_OPC6_REG5 is

   port( INSTR : in std_logic_vector (31 downto 0);  IMM : out std_logic_vector
         (31 downto 0));

end SIGNEX_N32_OPC6_REG5;

architecture SYN_BEHAVIORAL of SIGNEX_N32_OPC6_REG5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n1, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24 : std_logic;

begin
   
   U82 : NAND3_X1 port map( A1 => n47, A2 => n3, A3 => INSTR(26), ZN => n43);
   U83 : OAI33_X1 port map( A1 => n5, A2 => INSTR(30), A3 => INSTR(28), B1 => 
                           n48, B2 => INSTR(29), B3 => n7, ZN => n47);
   U2 : NAND2_X1 port map( A1 => n29, A2 => n27, ZN => n25);
   U3 : INV_X1 port map( A => n45, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n32, A2 => n27, ZN => n34);
   U5 : AND2_X1 port map( A1 => n28, A2 => n29, ZN => n32);
   U6 : INV_X1 port map( A => INSTR(26), ZN => n8);
   U7 : OAI21_X1 port map( B1 => n29, B2 => n10, A => n30, ZN => IMM(30));
   U8 : OAI21_X1 port map( B1 => n29, B2 => n11, A => n30, ZN => IMM(29));
   U9 : OAI21_X1 port map( B1 => n29, B2 => n12, A => n30, ZN => IMM(28));
   U10 : OAI21_X1 port map( B1 => n29, B2 => n13, A => n30, ZN => IMM(27));
   U11 : OAI21_X1 port map( B1 => n29, B2 => n14, A => n30, ZN => IMM(26));
   U12 : OAI21_X1 port map( B1 => n15, B2 => n29, A => n30, ZN => IMM(25));
   U13 : NOR2_X1 port map( A1 => n25, A2 => n10, ZN => IMM(14));
   U14 : NOR2_X1 port map( A1 => n25, A2 => n11, ZN => IMM(13));
   U15 : NOR2_X1 port map( A1 => n25, A2 => n12, ZN => IMM(12));
   U16 : NOR2_X1 port map( A1 => n25, A2 => n13, ZN => IMM(11));
   U17 : NOR2_X1 port map( A1 => n25, A2 => n14, ZN => IMM(10));
   U18 : NOR2_X1 port map( A1 => n25, A2 => n15, ZN => IMM(9));
   U19 : NOR2_X1 port map( A1 => n25, A2 => n16, ZN => IMM(8));
   U20 : NOR2_X1 port map( A1 => n25, A2 => n17, ZN => IMM(7));
   U21 : NOR2_X1 port map( A1 => n25, A2 => n18, ZN => IMM(6));
   U22 : NOR2_X1 port map( A1 => n25, A2 => n19, ZN => IMM(5));
   U23 : NOR2_X1 port map( A1 => n25, A2 => n20, ZN => IMM(4));
   U24 : NOR2_X1 port map( A1 => n25, A2 => n21, ZN => IMM(3));
   U25 : NOR2_X1 port map( A1 => n25, A2 => n22, ZN => IMM(2));
   U26 : NOR2_X1 port map( A1 => n25, A2 => n23, ZN => IMM(1));
   U27 : NOR2_X1 port map( A1 => n25, A2 => n24, ZN => IMM(0));
   U28 : NAND4_X1 port map( A1 => n7, A2 => n6, A3 => n8, A4 => n50, ZN => n27)
                           ;
   U29 : NAND2_X1 port map( A1 => n1, A2 => n27, ZN => n30);
   U30 : INV_X1 port map( A => n31, ZN => n1);
   U31 : AOI21_X1 port map( B1 => n4, B2 => INSTR(25), A => n32, ZN => n31);
   U32 : INV_X1 port map( A => INSTR(28), ZN => n6);
   U33 : INV_X1 port map( A => INSTR(29), ZN => n5);
   U34 : INV_X1 port map( A => INSTR(14), ZN => n10);
   U35 : INV_X1 port map( A => INSTR(13), ZN => n11);
   U36 : INV_X1 port map( A => INSTR(12), ZN => n12);
   U37 : INV_X1 port map( A => INSTR(11), ZN => n13);
   U38 : INV_X1 port map( A => INSTR(10), ZN => n14);
   U39 : INV_X1 port map( A => INSTR(2), ZN => n22);
   U40 : INV_X1 port map( A => INSTR(1), ZN => n23);
   U41 : INV_X1 port map( A => INSTR(0), ZN => n24);
   U42 : AND4_X1 port map( A1 => INSTR(15), A2 => n43, A3 => n44, A4 => n45, ZN
                           => n28);
   U43 : INV_X1 port map( A => INSTR(31), ZN => n3);
   U44 : INV_X1 port map( A => INSTR(9), ZN => n15);
   U45 : INV_X1 port map( A => INSTR(8), ZN => n16);
   U46 : INV_X1 port map( A => INSTR(7), ZN => n17);
   U47 : INV_X1 port map( A => INSTR(6), ZN => n18);
   U48 : INV_X1 port map( A => INSTR(5), ZN => n19);
   U49 : INV_X1 port map( A => INSTR(4), ZN => n20);
   U50 : INV_X1 port map( A => INSTR(3), ZN => n21);
   U51 : OAI211_X1 port map( C1 => n29, C2 => n22, A => n40, B => n34, ZN => 
                           IMM(18));
   U52 : NAND2_X1 port map( A1 => INSTR(18), A2 => n4, ZN => n40);
   U53 : OAI211_X1 port map( C1 => n29, C2 => n23, A => n41, B => n34, ZN => 
                           IMM(17));
   U54 : NAND2_X1 port map( A1 => INSTR(17), A2 => n4, ZN => n41);
   U55 : OAI211_X1 port map( C1 => n29, C2 => n24, A => n42, B => n34, ZN => 
                           IMM(16));
   U56 : NAND2_X1 port map( A1 => INSTR(16), A2 => n4, ZN => n42);
   U57 : OAI211_X1 port map( C1 => n16, C2 => n29, A => n33, B => n34, ZN => 
                           IMM(24));
   U58 : NAND2_X1 port map( A1 => INSTR(24), A2 => n4, ZN => n33);
   U59 : OAI211_X1 port map( C1 => n17, C2 => n29, A => n35, B => n34, ZN => 
                           IMM(23));
   U60 : NAND2_X1 port map( A1 => INSTR(23), A2 => n4, ZN => n35);
   U61 : OAI211_X1 port map( C1 => n18, C2 => n29, A => n36, B => n34, ZN => 
                           IMM(22));
   U62 : NAND2_X1 port map( A1 => INSTR(22), A2 => n4, ZN => n36);
   U63 : OAI211_X1 port map( C1 => n19, C2 => n29, A => n37, B => n34, ZN => 
                           IMM(21));
   U64 : NAND2_X1 port map( A1 => INSTR(21), A2 => n4, ZN => n37);
   U65 : OAI211_X1 port map( C1 => n20, C2 => n29, A => n38, B => n34, ZN => 
                           IMM(20));
   U66 : NAND2_X1 port map( A1 => INSTR(20), A2 => n4, ZN => n38);
   U67 : OAI211_X1 port map( C1 => n21, C2 => n29, A => n39, B => n34, ZN => 
                           IMM(19));
   U68 : NAND2_X1 port map( A1 => INSTR(19), A2 => n4, ZN => n39);
   U69 : NOR2_X1 port map( A1 => n25, A2 => n9, ZN => IMM(15));
   U70 : INV_X1 port map( A => INSTR(15), ZN => n9);
   U71 : INV_X1 port map( A => n26, ZN => IMM(31));
   U72 : AOI22_X1 port map( A1 => n4, A2 => INSTR(25), B1 => n27, B2 => n28, ZN
                           => n26);
   U73 : NAND4_X1 port map( A1 => INSTR(31), A2 => INSTR(30), A3 => INSTR(29), 
                           A4 => n46, ZN => n44);
   U74 : NAND2_X1 port map( A1 => INSTR(30), A2 => INSTR(28), ZN => n48);
   U75 : NOR2_X1 port map( A1 => INSTR(31), A2 => INSTR(30), ZN => n49);
   U76 : NOR3_X1 port map( A1 => INSTR(29), A2 => INSTR(31), A3 => INSTR(30), 
                           ZN => n50);
   U77 : NOR3_X1 port map( A1 => n8, A2 => INSTR(31), A3 => INSTR(30), ZN => 
                           n51);
   U78 : XNOR2_X1 port map( A => n6, B => INSTR(27), ZN => n46);
   U79 : NAND4_X1 port map( A1 => INSTR(27), A2 => n6, A3 => n49, A4 => n5, ZN 
                           => n45);
   U80 : INV_X1 port map( A => INSTR(27), ZN => n7);
   U81 : NAND4_X1 port map( A1 => INSTR(28), A2 => INSTR(27), A3 => INSTR(29), 
                           A4 => n51, ZN => n29);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RF_N32_NA5 is

   port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
         ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_N32_NA5;

architecture SYN_BEHAVIORAL of RF_N32_NA5 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REG_0_31_port, REG_0_30_port, REG_0_29_port, REG_0_28_port, 
      REG_0_27_port, REG_0_26_port, REG_0_25_port, REG_0_24_port, REG_0_23_port
      , REG_0_22_port, REG_0_21_port, REG_0_20_port, REG_0_19_port, 
      REG_0_18_port, REG_0_17_port, REG_0_16_port, REG_0_15_port, REG_0_14_port
      , REG_0_13_port, REG_0_12_port, REG_0_11_port, REG_0_10_port, 
      REG_0_9_port, REG_0_8_port, REG_0_7_port, REG_0_6_port, REG_0_5_port, 
      REG_0_4_port, REG_0_3_port, REG_0_2_port, REG_0_1_port, REG_0_0_port, 
      REG_1_31_port, REG_1_30_port, REG_1_29_port, REG_1_28_port, REG_1_27_port
      , REG_1_26_port, REG_1_25_port, REG_1_24_port, REG_1_23_port, 
      REG_1_22_port, REG_1_21_port, REG_1_20_port, REG_1_19_port, REG_1_18_port
      , REG_1_17_port, REG_1_16_port, REG_1_15_port, REG_1_14_port, 
      REG_1_13_port, REG_1_12_port, REG_1_11_port, REG_1_10_port, REG_1_9_port,
      REG_1_8_port, REG_1_7_port, REG_1_6_port, REG_1_5_port, REG_1_4_port, 
      REG_1_3_port, REG_1_2_port, REG_1_1_port, REG_1_0_port, REG_2_31_port, 
      REG_2_30_port, REG_2_29_port, REG_2_28_port, REG_2_27_port, REG_2_26_port
      , REG_2_25_port, REG_2_24_port, REG_2_23_port, REG_2_22_port, 
      REG_2_21_port, REG_2_20_port, REG_2_19_port, REG_2_18_port, REG_2_17_port
      , REG_2_16_port, REG_2_15_port, REG_2_14_port, REG_2_13_port, 
      REG_2_12_port, REG_2_11_port, REG_2_10_port, REG_2_9_port, REG_2_8_port, 
      REG_2_7_port, REG_2_6_port, REG_2_5_port, REG_2_4_port, REG_2_3_port, 
      REG_2_2_port, REG_2_1_port, REG_2_0_port, REG_3_31_port, REG_3_30_port, 
      REG_3_29_port, REG_3_28_port, REG_3_27_port, REG_3_26_port, REG_3_25_port
      , REG_3_24_port, REG_3_23_port, REG_3_22_port, REG_3_21_port, 
      REG_3_20_port, REG_3_19_port, REG_3_18_port, REG_3_17_port, REG_3_16_port
      , REG_3_15_port, REG_3_14_port, REG_3_13_port, REG_3_12_port, 
      REG_3_11_port, REG_3_10_port, REG_3_9_port, REG_3_8_port, REG_3_7_port, 
      REG_3_6_port, REG_3_5_port, REG_3_4_port, REG_3_3_port, REG_3_2_port, 
      REG_3_1_port, REG_3_0_port, REG_4_31_port, REG_4_30_port, REG_4_29_port, 
      REG_4_28_port, REG_4_27_port, REG_4_26_port, REG_4_25_port, REG_4_24_port
      , REG_4_23_port, REG_4_22_port, REG_4_21_port, REG_4_20_port, 
      REG_4_19_port, REG_4_18_port, REG_4_17_port, REG_4_16_port, REG_4_15_port
      , REG_4_14_port, REG_4_13_port, REG_4_12_port, REG_4_11_port, 
      REG_4_10_port, REG_4_9_port, REG_4_8_port, REG_4_7_port, REG_4_6_port, 
      REG_4_5_port, REG_4_4_port, REG_4_3_port, REG_4_2_port, REG_4_1_port, 
      REG_4_0_port, REG_5_31_port, REG_5_30_port, REG_5_29_port, REG_5_28_port,
      REG_5_27_port, REG_5_26_port, REG_5_25_port, REG_5_24_port, REG_5_23_port
      , REG_5_22_port, REG_5_21_port, REG_5_20_port, REG_5_19_port, 
      REG_5_18_port, REG_5_17_port, REG_5_16_port, REG_5_15_port, REG_5_14_port
      , REG_5_13_port, REG_5_12_port, REG_5_11_port, REG_5_10_port, 
      REG_5_9_port, REG_5_8_port, REG_5_7_port, REG_5_6_port, REG_5_5_port, 
      REG_5_4_port, REG_5_3_port, REG_5_2_port, REG_5_1_port, REG_5_0_port, 
      REG_6_31_port, REG_6_30_port, REG_6_29_port, REG_6_28_port, REG_6_27_port
      , REG_6_26_port, REG_6_25_port, REG_6_24_port, REG_6_23_port, 
      REG_6_22_port, REG_6_21_port, REG_6_20_port, REG_6_19_port, REG_6_18_port
      , REG_6_17_port, REG_6_16_port, REG_6_15_port, REG_6_14_port, 
      REG_6_13_port, REG_6_12_port, REG_6_11_port, REG_6_10_port, REG_6_9_port,
      REG_6_8_port, REG_6_7_port, REG_6_6_port, REG_6_5_port, REG_6_4_port, 
      REG_6_3_port, REG_6_2_port, REG_6_1_port, REG_6_0_port, REG_7_31_port, 
      REG_7_30_port, REG_7_29_port, REG_7_28_port, REG_7_27_port, REG_7_26_port
      , REG_7_25_port, REG_7_24_port, REG_7_23_port, REG_7_22_port, 
      REG_7_21_port, REG_7_20_port, REG_7_19_port, REG_7_18_port, REG_7_17_port
      , REG_7_16_port, REG_7_15_port, REG_7_14_port, REG_7_13_port, 
      REG_7_12_port, REG_7_11_port, REG_7_10_port, REG_7_9_port, REG_7_8_port, 
      REG_7_7_port, REG_7_6_port, REG_7_5_port, REG_7_4_port, REG_7_3_port, 
      REG_7_2_port, REG_7_1_port, REG_7_0_port, REG_8_31_port, REG_8_30_port, 
      REG_8_29_port, REG_8_28_port, REG_8_27_port, REG_8_26_port, REG_8_25_port
      , REG_8_24_port, REG_8_23_port, REG_8_22_port, REG_8_21_port, 
      REG_8_20_port, REG_8_19_port, REG_8_18_port, REG_8_17_port, REG_8_16_port
      , REG_8_15_port, REG_8_14_port, REG_8_13_port, REG_8_12_port, 
      REG_8_11_port, REG_8_10_port, REG_8_9_port, REG_8_8_port, REG_8_7_port, 
      REG_8_6_port, REG_8_5_port, REG_8_4_port, REG_8_3_port, REG_8_2_port, 
      REG_8_1_port, REG_8_0_port, REG_9_31_port, REG_9_30_port, REG_9_29_port, 
      REG_9_28_port, REG_9_27_port, REG_9_26_port, REG_9_25_port, REG_9_24_port
      , REG_9_23_port, REG_9_22_port, REG_9_21_port, REG_9_20_port, 
      REG_9_19_port, REG_9_18_port, REG_9_17_port, REG_9_16_port, REG_9_15_port
      , REG_9_14_port, REG_9_13_port, REG_9_12_port, REG_9_11_port, 
      REG_9_10_port, REG_9_9_port, REG_9_8_port, REG_9_7_port, REG_9_6_port, 
      REG_9_5_port, REG_9_4_port, REG_9_3_port, REG_9_2_port, REG_9_1_port, 
      REG_9_0_port, REG_10_31_port, REG_10_30_port, REG_10_29_port, 
      REG_10_28_port, REG_10_27_port, REG_10_26_port, REG_10_25_port, 
      REG_10_24_port, REG_10_23_port, REG_10_22_port, REG_10_21_port, 
      REG_10_20_port, REG_10_19_port, REG_10_18_port, REG_10_17_port, 
      REG_10_16_port, REG_10_15_port, REG_10_14_port, REG_10_13_port, 
      REG_10_12_port, REG_10_11_port, REG_10_10_port, REG_10_9_port, 
      REG_10_8_port, REG_10_7_port, REG_10_6_port, REG_10_5_port, REG_10_4_port
      , REG_10_3_port, REG_10_2_port, REG_10_1_port, REG_10_0_port, 
      REG_11_31_port, REG_11_30_port, REG_11_29_port, REG_11_28_port, 
      REG_11_27_port, REG_11_26_port, REG_11_25_port, REG_11_24_port, 
      REG_11_23_port, REG_11_22_port, REG_11_21_port, REG_11_20_port, 
      REG_11_19_port, REG_11_18_port, REG_11_17_port, REG_11_16_port, 
      REG_11_15_port, REG_11_14_port, REG_11_13_port, REG_11_12_port, 
      REG_11_11_port, REG_11_10_port, REG_11_9_port, REG_11_8_port, 
      REG_11_7_port, REG_11_6_port, REG_11_5_port, REG_11_4_port, REG_11_3_port
      , REG_11_2_port, REG_11_1_port, REG_11_0_port, REG_12_31_port, 
      REG_12_30_port, REG_12_29_port, REG_12_28_port, REG_12_27_port, 
      REG_12_26_port, REG_12_25_port, REG_12_24_port, REG_12_23_port, 
      REG_12_22_port, REG_12_21_port, REG_12_20_port, REG_12_19_port, 
      REG_12_18_port, REG_12_17_port, REG_12_16_port, REG_12_15_port, 
      REG_12_14_port, REG_12_13_port, REG_12_12_port, REG_12_11_port, 
      REG_12_10_port, REG_12_9_port, REG_12_8_port, REG_12_7_port, 
      REG_12_6_port, REG_12_5_port, REG_12_4_port, REG_12_3_port, REG_12_2_port
      , REG_12_1_port, REG_12_0_port, REG_13_31_port, REG_13_30_port, 
      REG_13_29_port, REG_13_28_port, REG_13_27_port, REG_13_26_port, 
      REG_13_25_port, REG_13_24_port, REG_13_23_port, REG_13_22_port, 
      REG_13_21_port, REG_13_20_port, REG_13_19_port, REG_13_18_port, 
      REG_13_17_port, REG_13_16_port, REG_13_15_port, REG_13_14_port, 
      REG_13_13_port, REG_13_12_port, REG_13_11_port, REG_13_10_port, 
      REG_13_9_port, REG_13_8_port, REG_13_7_port, REG_13_6_port, REG_13_5_port
      , REG_13_4_port, REG_13_3_port, REG_13_2_port, REG_13_1_port, 
      REG_13_0_port, REG_14_31_port, REG_14_30_port, REG_14_29_port, 
      REG_14_28_port, REG_14_27_port, REG_14_26_port, REG_14_25_port, 
      REG_14_24_port, REG_14_23_port, REG_14_22_port, REG_14_21_port, 
      REG_14_20_port, REG_14_19_port, REG_14_18_port, REG_14_17_port, 
      REG_14_16_port, REG_14_15_port, REG_14_14_port, REG_14_13_port, 
      REG_14_12_port, REG_14_11_port, REG_14_10_port, REG_14_9_port, 
      REG_14_8_port, REG_14_7_port, REG_14_6_port, REG_14_5_port, REG_14_4_port
      , REG_14_3_port, REG_14_2_port, REG_14_1_port, REG_14_0_port, 
      REG_15_31_port, REG_15_30_port, REG_15_29_port, REG_15_28_port, 
      REG_15_27_port, REG_15_26_port, REG_15_25_port, REG_15_24_port, 
      REG_15_23_port, REG_15_22_port, REG_15_21_port, REG_15_20_port, 
      REG_15_19_port, REG_15_18_port, REG_15_17_port, REG_15_16_port, 
      REG_15_15_port, REG_15_14_port, REG_15_13_port, REG_15_12_port, 
      REG_15_11_port, REG_15_10_port, REG_15_9_port, REG_15_8_port, 
      REG_15_7_port, REG_15_6_port, REG_15_5_port, REG_15_4_port, REG_15_3_port
      , REG_15_2_port, REG_15_1_port, REG_15_0_port, REG_16_31_port, 
      REG_16_30_port, REG_16_29_port, REG_16_28_port, REG_16_27_port, 
      REG_16_26_port, REG_16_25_port, REG_16_24_port, REG_16_23_port, 
      REG_16_22_port, REG_16_21_port, REG_16_20_port, REG_16_19_port, 
      REG_16_18_port, REG_16_17_port, REG_16_16_port, REG_16_15_port, 
      REG_16_14_port, REG_16_13_port, REG_16_12_port, REG_16_11_port, 
      REG_16_10_port, REG_16_9_port, REG_16_8_port, REG_16_7_port, 
      REG_16_6_port, REG_16_5_port, REG_16_4_port, REG_16_3_port, REG_16_2_port
      , REG_16_1_port, REG_16_0_port, REG_17_31_port, REG_17_30_port, 
      REG_17_29_port, REG_17_28_port, REG_17_27_port, REG_17_26_port, 
      REG_17_25_port, REG_17_24_port, REG_17_23_port, REG_17_22_port, 
      REG_17_21_port, REG_17_20_port, REG_17_19_port, REG_17_18_port, 
      REG_17_17_port, REG_17_16_port, REG_17_15_port, REG_17_14_port, 
      REG_17_13_port, REG_17_12_port, REG_17_11_port, REG_17_10_port, 
      REG_17_9_port, REG_17_8_port, REG_17_7_port, REG_17_6_port, REG_17_5_port
      , REG_17_4_port, REG_17_3_port, REG_17_2_port, REG_17_1_port, 
      REG_17_0_port, REG_18_31_port, REG_18_30_port, REG_18_29_port, 
      REG_18_28_port, REG_18_27_port, REG_18_26_port, REG_18_25_port, 
      REG_18_24_port, REG_18_23_port, REG_18_22_port, REG_18_21_port, 
      REG_18_20_port, REG_18_19_port, REG_18_18_port, REG_18_17_port, 
      REG_18_16_port, REG_18_15_port, REG_18_14_port, REG_18_13_port, 
      REG_18_12_port, REG_18_11_port, REG_18_10_port, REG_18_9_port, 
      REG_18_8_port, REG_18_7_port, REG_18_6_port, REG_18_5_port, REG_18_4_port
      , REG_18_3_port, REG_18_2_port, REG_18_1_port, REG_18_0_port, 
      REG_19_31_port, REG_19_30_port, REG_19_29_port, REG_19_28_port, 
      REG_19_27_port, REG_19_26_port, REG_19_25_port, REG_19_24_port, 
      REG_19_23_port, REG_19_22_port, REG_19_21_port, REG_19_20_port, 
      REG_19_19_port, REG_19_18_port, REG_19_17_port, REG_19_16_port, 
      REG_19_15_port, REG_19_14_port, REG_19_13_port, REG_19_12_port, 
      REG_19_11_port, REG_19_10_port, REG_19_9_port, REG_19_8_port, 
      REG_19_7_port, REG_19_6_port, REG_19_5_port, REG_19_4_port, REG_19_3_port
      , REG_19_2_port, REG_19_1_port, REG_19_0_port, REG_20_31_port, 
      REG_20_30_port, REG_20_29_port, REG_20_28_port, REG_20_27_port, 
      REG_20_26_port, REG_20_25_port, REG_20_24_port, REG_20_23_port, 
      REG_20_22_port, REG_20_21_port, REG_20_20_port, REG_20_19_port, 
      REG_20_18_port, REG_20_17_port, REG_20_16_port, REG_20_15_port, 
      REG_20_14_port, REG_20_13_port, REG_20_12_port, REG_20_11_port, 
      REG_20_10_port, REG_20_9_port, REG_20_8_port, REG_20_7_port, 
      REG_20_6_port, REG_20_5_port, REG_20_4_port, REG_20_3_port, REG_20_2_port
      , REG_20_1_port, REG_20_0_port, REG_21_31_port, REG_21_30_port, 
      REG_21_29_port, REG_21_28_port, REG_21_27_port, REG_21_26_port, 
      REG_21_25_port, REG_21_24_port, REG_21_23_port, REG_21_22_port, 
      REG_21_21_port, REG_21_20_port, REG_21_19_port, REG_21_18_port, 
      REG_21_17_port, REG_21_16_port, REG_21_15_port, REG_21_14_port, 
      REG_21_13_port, REG_21_12_port, REG_21_11_port, REG_21_10_port, 
      REG_21_9_port, REG_21_8_port, REG_21_7_port, REG_21_6_port, REG_21_5_port
      , REG_21_4_port, REG_21_3_port, REG_21_2_port, REG_21_1_port, 
      REG_21_0_port, REG_22_31_port, REG_22_30_port, REG_22_29_port, 
      REG_22_28_port, REG_22_27_port, REG_22_26_port, REG_22_25_port, 
      REG_22_24_port, REG_22_23_port, REG_22_22_port, REG_22_21_port, 
      REG_22_20_port, REG_22_19_port, REG_22_18_port, REG_22_17_port, 
      REG_22_16_port, REG_22_15_port, REG_22_14_port, REG_22_13_port, 
      REG_22_12_port, REG_22_11_port, REG_22_10_port, REG_22_9_port, 
      REG_22_8_port, REG_22_7_port, REG_22_6_port, REG_22_5_port, REG_22_4_port
      , REG_22_3_port, REG_22_2_port, REG_22_1_port, REG_22_0_port, 
      REG_23_31_port, REG_23_30_port, REG_23_29_port, REG_23_28_port, 
      REG_23_27_port, REG_23_26_port, REG_23_25_port, REG_23_24_port, 
      REG_23_23_port, REG_23_22_port, REG_23_21_port, REG_23_20_port, 
      REG_23_19_port, REG_23_18_port, REG_23_17_port, REG_23_16_port, 
      REG_23_15_port, REG_23_14_port, REG_23_13_port, REG_23_12_port, 
      REG_23_11_port, REG_23_10_port, REG_23_9_port, REG_23_8_port, 
      REG_23_7_port, REG_23_6_port, REG_23_5_port, REG_23_4_port, REG_23_3_port
      , REG_23_2_port, REG_23_1_port, REG_23_0_port, REG_24_31_port, 
      REG_24_30_port, REG_24_29_port, REG_24_28_port, REG_24_27_port, 
      REG_24_26_port, REG_24_25_port, REG_24_24_port, REG_24_23_port, 
      REG_24_22_port, REG_24_21_port, REG_24_20_port, REG_24_19_port, 
      REG_24_18_port, REG_24_17_port, REG_24_16_port, REG_24_15_port, 
      REG_24_14_port, REG_24_13_port, REG_24_12_port, REG_24_11_port, 
      REG_24_10_port, REG_24_9_port, REG_24_8_port, REG_24_7_port, 
      REG_24_6_port, REG_24_5_port, REG_24_4_port, REG_24_3_port, REG_24_2_port
      , REG_24_1_port, REG_24_0_port, REG_25_31_port, REG_25_30_port, 
      REG_25_29_port, REG_25_28_port, REG_25_27_port, REG_25_26_port, 
      REG_25_25_port, REG_25_24_port, REG_25_23_port, REG_25_22_port, 
      REG_25_21_port, REG_25_20_port, REG_25_19_port, REG_25_18_port, 
      REG_25_17_port, REG_25_16_port, REG_25_15_port, REG_25_14_port, 
      REG_25_13_port, REG_25_12_port, REG_25_11_port, REG_25_10_port, 
      REG_25_9_port, REG_25_8_port, REG_25_7_port, REG_25_6_port, REG_25_5_port
      , REG_25_4_port, REG_25_3_port, REG_25_2_port, REG_25_1_port, 
      REG_25_0_port, REG_26_31_port, REG_26_30_port, REG_26_29_port, 
      REG_26_28_port, REG_26_27_port, REG_26_26_port, REG_26_25_port, 
      REG_26_24_port, REG_26_23_port, REG_26_22_port, REG_26_21_port, 
      REG_26_20_port, REG_26_19_port, REG_26_18_port, REG_26_17_port, 
      REG_26_16_port, REG_26_15_port, REG_26_14_port, REG_26_13_port, 
      REG_26_12_port, REG_26_11_port, REG_26_10_port, REG_26_9_port, 
      REG_26_8_port, REG_26_7_port, REG_26_6_port, REG_26_5_port, REG_26_4_port
      , REG_26_3_port, REG_26_2_port, REG_26_1_port, REG_26_0_port, 
      REG_27_31_port, REG_27_30_port, REG_27_29_port, REG_27_28_port, 
      REG_27_27_port, REG_27_26_port, REG_27_25_port, REG_27_24_port, 
      REG_27_23_port, REG_27_22_port, REG_27_21_port, REG_27_20_port, 
      REG_27_19_port, REG_27_18_port, REG_27_17_port, REG_27_16_port, 
      REG_27_15_port, REG_27_14_port, REG_27_13_port, REG_27_12_port, 
      REG_27_11_port, REG_27_10_port, REG_27_9_port, REG_27_8_port, 
      REG_27_7_port, REG_27_6_port, REG_27_5_port, REG_27_4_port, REG_27_3_port
      , REG_27_2_port, REG_27_1_port, REG_27_0_port, REG_28_31_port, 
      REG_28_30_port, REG_28_29_port, REG_28_28_port, REG_28_27_port, 
      REG_28_26_port, REG_28_25_port, REG_28_24_port, REG_28_23_port, 
      REG_28_22_port, REG_28_21_port, REG_28_20_port, REG_28_19_port, 
      REG_28_18_port, REG_28_17_port, REG_28_16_port, REG_28_15_port, 
      REG_28_14_port, REG_28_13_port, REG_28_12_port, REG_28_11_port, 
      REG_28_10_port, REG_28_9_port, REG_28_8_port, REG_28_7_port, 
      REG_28_6_port, REG_28_5_port, REG_28_4_port, REG_28_3_port, REG_28_2_port
      , REG_28_1_port, REG_28_0_port, REG_29_31_port, REG_29_30_port, 
      REG_29_29_port, REG_29_28_port, REG_29_27_port, REG_29_26_port, 
      REG_29_25_port, REG_29_24_port, REG_29_23_port, REG_29_22_port, 
      REG_29_21_port, REG_29_20_port, REG_29_19_port, REG_29_18_port, 
      REG_29_17_port, REG_29_16_port, REG_29_15_port, REG_29_14_port, 
      REG_29_13_port, REG_29_12_port, REG_29_11_port, REG_29_10_port, 
      REG_29_9_port, REG_29_8_port, REG_29_7_port, REG_29_6_port, REG_29_5_port
      , REG_29_4_port, REG_29_3_port, REG_29_2_port, REG_29_1_port, 
      REG_29_0_port, REG_30_31_port, REG_30_30_port, REG_30_29_port, 
      REG_30_28_port, REG_30_27_port, REG_30_26_port, REG_30_25_port, 
      REG_30_24_port, REG_30_23_port, REG_30_22_port, REG_30_21_port, 
      REG_30_20_port, REG_30_19_port, REG_30_18_port, REG_30_17_port, 
      REG_30_16_port, REG_30_15_port, REG_30_14_port, REG_30_13_port, 
      REG_30_12_port, REG_30_11_port, REG_30_10_port, REG_30_9_port, 
      REG_30_8_port, REG_30_7_port, REG_30_6_port, REG_30_5_port, REG_30_4_port
      , REG_30_3_port, REG_30_2_port, REG_30_1_port, REG_30_0_port, 
      REG_31_31_port, REG_31_30_port, REG_31_29_port, REG_31_28_port, 
      REG_31_27_port, REG_31_26_port, REG_31_25_port, REG_31_24_port, 
      REG_31_23_port, REG_31_22_port, REG_31_21_port, REG_31_20_port, 
      REG_31_19_port, REG_31_18_port, REG_31_17_port, REG_31_16_port, 
      REG_31_15_port, REG_31_14_port, REG_31_13_port, REG_31_12_port, 
      REG_31_11_port, REG_31_10_port, REG_31_9_port, REG_31_8_port, 
      REG_31_7_port, REG_31_6_port, REG_31_5_port, REG_31_4_port, REG_31_3_port
      , REG_31_2_port, REG_31_1_port, REG_31_0_port, N155, N188, N189, N190, 
      N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, 
      N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, 
      N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, 
      N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, 
      N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, 
      N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, 
      N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, 
      N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, 
      N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, 
      N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, 
      N312, N313, N314, N315, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155_port, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188_port, n189_port, n190_port, n191_port,
      n192_port, n193_port, n194_port, n195_port, n196_port, n197_port, 
      n198_port, n199_port, n200_port, n201_port, n202_port, n203_port, 
      n204_port, n205_port, n206_port, n207_port, n208_port, n209_port, 
      n210_port, n211_port, n212_port, n213_port, n214_port, n215_port, 
      n216_port, n217_port, n218_port, n219_port, n220_port, n221_port, 
      n222_port, n223_port, n224_port, n225_port, n226_port, n227_port, 
      n228_port, n229_port, n230_port, n231_port, n232_port, n233_port, 
      n234_port, n235_port, n236_port, n237_port, n238_port, n239_port, 
      n240_port, n241_port, n242_port, n243_port, n244_port, n245_port, 
      n246_port, n247_port, n248_port, n249_port, n250_port, n251, n252_port, 
      n253_port, n254_port, n255_port, n256_port, n257_port, n258_port, 
      n259_port, n260_port, n261_port, n262_port, n263_port, n264_port, 
      n265_port, n266_port, n267_port, n268_port, n269_port, n270_port, 
      n271_port, n272_port, n273_port, n274_port, n275_port, n276_port, 
      n277_port, n278_port, n279_port, n280_port, n281_port, n282_port, 
      n283_port, n284_port, n285_port, n286_port, n287_port, n288_port, 
      n289_port, n290_port, n291_port, n292_port, n293_port, n294_port, 
      n295_port, n296_port, n297_port, n298_port, n299_port, n300_port, 
      n301_port, n302_port, n303_port, n304_port, n305_port, n306_port, 
      n307_port, n308_port, n309_port, n310_port, n311_port, n312_port, 
      n313_port, n314_port, n315_port, n316, n317, n318, n319, n320, n321, n322
      , n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
      n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
      n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, 
      n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, 
      n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, 
      n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, 
      n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, 
      n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
      n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
      n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, 
      n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, 
      n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, 
      n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
      n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
      n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, 
      n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
      n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, 
      n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, 
      n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, 
      n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, 
      n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
      n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, 
      n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, 
      n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, 
      n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, 
      n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, 
      n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, 
      n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, 
      n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, 
      n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, 
      n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, 
      n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, 
      n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, 
      n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, 
      n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, 
      n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, 
      n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, 
      n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, 
      n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, 
      n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, 
      n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, 
      n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, 
      n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, 
      n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, 
      n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, 
      n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, 
      n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, 
      n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
      n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, 
      n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, 
      n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, 
      n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, 
      n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, 
      n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, 
      n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, 
      n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, 
      n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, 
      n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, 
      n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, 
      n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, 
      n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, 
      n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, 
      n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, 
      n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, 
      n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
      n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, 
      n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
      n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, 
      n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
      n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, 
      n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
      n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, 
      n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, 
      n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, 
      n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, 
      n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, 
      n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, 
      n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, 
      n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, 
      n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, 
      n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, 
      n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, 
      n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, 
      n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
      n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, 
      n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, 
      n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, 
      n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, 
      n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, 
      n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, 
      n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, 
      n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, 
      n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, 
      n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, 
      n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, 
      n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, 
      n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, 
      n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, 
      n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, 
      n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, 
      n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, 
      n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, 
      n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, 
      n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, 
      n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, 
      n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, 
      n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, 
      n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, 
      n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
      n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, 
      n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, 
      n2096, n2097 : std_logic;

begin
   
   REG_reg_0_31_inst : DLH_X1 port map( G => n1839, D => N250, Q => 
                           REG_0_31_port);
   REG_reg_0_30_inst : DLH_X1 port map( G => n1839, D => N249, Q => 
                           REG_0_30_port);
   REG_reg_0_29_inst : DLH_X1 port map( G => n1838, D => N248, Q => 
                           REG_0_29_port);
   REG_reg_0_28_inst : DLH_X1 port map( G => n1838, D => N247, Q => 
                           REG_0_28_port);
   REG_reg_0_27_inst : DLH_X1 port map( G => n1838, D => N246, Q => 
                           REG_0_27_port);
   REG_reg_0_26_inst : DLH_X1 port map( G => n1838, D => N245, Q => 
                           REG_0_26_port);
   REG_reg_0_25_inst : DLH_X1 port map( G => n1838, D => N244, Q => 
                           REG_0_25_port);
   REG_reg_0_24_inst : DLH_X1 port map( G => n1838, D => N243, Q => 
                           REG_0_24_port);
   REG_reg_0_23_inst : DLH_X1 port map( G => n1838, D => N242, Q => 
                           REG_0_23_port);
   REG_reg_0_22_inst : DLH_X1 port map( G => n1838, D => N241, Q => 
                           REG_0_22_port);
   REG_reg_0_21_inst : DLH_X1 port map( G => n1838, D => N240, Q => 
                           REG_0_21_port);
   REG_reg_0_20_inst : DLH_X1 port map( G => n1838, D => N239, Q => 
                           REG_0_20_port);
   REG_reg_0_19_inst : DLH_X1 port map( G => n1837, D => N238, Q => 
                           REG_0_19_port);
   REG_reg_0_18_inst : DLH_X1 port map( G => n1837, D => N237, Q => 
                           REG_0_18_port);
   REG_reg_0_17_inst : DLH_X1 port map( G => n1837, D => N236, Q => 
                           REG_0_17_port);
   REG_reg_0_16_inst : DLH_X1 port map( G => n1837, D => N235, Q => 
                           REG_0_16_port);
   REG_reg_0_15_inst : DLH_X1 port map( G => n1837, D => N234, Q => 
                           REG_0_15_port);
   REG_reg_0_14_inst : DLH_X1 port map( G => n1837, D => N233, Q => 
                           REG_0_14_port);
   REG_reg_0_13_inst : DLH_X1 port map( G => n1837, D => N232, Q => 
                           REG_0_13_port);
   REG_reg_0_12_inst : DLH_X1 port map( G => n1837, D => N231, Q => 
                           REG_0_12_port);
   REG_reg_0_11_inst : DLH_X1 port map( G => n1837, D => N230, Q => 
                           REG_0_11_port);
   REG_reg_0_10_inst : DLH_X1 port map( G => n1837, D => N229, Q => 
                           REG_0_10_port);
   REG_reg_0_9_inst : DLH_X1 port map( G => n1836, D => N228, Q => REG_0_9_port
                           );
   REG_reg_0_8_inst : DLH_X1 port map( G => n1836, D => N227, Q => REG_0_8_port
                           );
   REG_reg_0_7_inst : DLH_X1 port map( G => n1836, D => N226, Q => REG_0_7_port
                           );
   REG_reg_0_6_inst : DLH_X1 port map( G => n1836, D => N225, Q => REG_0_6_port
                           );
   REG_reg_0_5_inst : DLH_X1 port map( G => n1836, D => N224, Q => REG_0_5_port
                           );
   REG_reg_0_4_inst : DLH_X1 port map( G => n1836, D => N223, Q => REG_0_4_port
                           );
   REG_reg_0_3_inst : DLH_X1 port map( G => n1836, D => N222, Q => REG_0_3_port
                           );
   REG_reg_0_2_inst : DLH_X1 port map( G => n1836, D => N221, Q => REG_0_2_port
                           );
   REG_reg_0_1_inst : DLH_X1 port map( G => n1836, D => N220, Q => REG_0_1_port
                           );
   REG_reg_0_0_inst : DLH_X1 port map( G => n1836, D => N219, Q => REG_0_0_port
                           );
   REG_reg_1_31_inst : DLH_X1 port map( G => n1846, D => n1629, Q => 
                           REG_1_31_port);
   REG_reg_1_30_inst : DLH_X1 port map( G => n1846, D => n1635, Q => 
                           REG_1_30_port);
   REG_reg_1_29_inst : DLH_X1 port map( G => n1845, D => n1641, Q => 
                           REG_1_29_port);
   REG_reg_1_28_inst : DLH_X1 port map( G => n1845, D => n1647, Q => 
                           REG_1_28_port);
   REG_reg_1_27_inst : DLH_X1 port map( G => n1845, D => n1653, Q => 
                           REG_1_27_port);
   REG_reg_1_26_inst : DLH_X1 port map( G => n1845, D => n1659, Q => 
                           REG_1_26_port);
   REG_reg_1_25_inst : DLH_X1 port map( G => n1845, D => n1665, Q => 
                           REG_1_25_port);
   REG_reg_1_24_inst : DLH_X1 port map( G => n1845, D => n1671, Q => 
                           REG_1_24_port);
   REG_reg_1_23_inst : DLH_X1 port map( G => n1845, D => n1677, Q => 
                           REG_1_23_port);
   REG_reg_1_22_inst : DLH_X1 port map( G => n1845, D => n1683, Q => 
                           REG_1_22_port);
   REG_reg_1_21_inst : DLH_X1 port map( G => n1845, D => n1689, Q => 
                           REG_1_21_port);
   REG_reg_1_20_inst : DLH_X1 port map( G => n1845, D => n1695, Q => 
                           REG_1_20_port);
   REG_reg_1_19_inst : DLH_X1 port map( G => n1844, D => n1701, Q => 
                           REG_1_19_port);
   REG_reg_1_18_inst : DLH_X1 port map( G => n1844, D => n1707, Q => 
                           REG_1_18_port);
   REG_reg_1_17_inst : DLH_X1 port map( G => n1844, D => n1713, Q => 
                           REG_1_17_port);
   REG_reg_1_16_inst : DLH_X1 port map( G => n1844, D => n1719, Q => 
                           REG_1_16_port);
   REG_reg_1_15_inst : DLH_X1 port map( G => n1844, D => n1725, Q => 
                           REG_1_15_port);
   REG_reg_1_14_inst : DLH_X1 port map( G => n1844, D => n1731, Q => 
                           REG_1_14_port);
   REG_reg_1_13_inst : DLH_X1 port map( G => n1844, D => n1737, Q => 
                           REG_1_13_port);
   REG_reg_1_12_inst : DLH_X1 port map( G => n1844, D => n1743, Q => 
                           REG_1_12_port);
   REG_reg_1_11_inst : DLH_X1 port map( G => n1844, D => n1749, Q => 
                           REG_1_11_port);
   REG_reg_1_10_inst : DLH_X1 port map( G => n1844, D => n1755, Q => 
                           REG_1_10_port);
   REG_reg_1_9_inst : DLH_X1 port map( G => n1843, D => n1761, Q => 
                           REG_1_9_port);
   REG_reg_1_8_inst : DLH_X1 port map( G => n1843, D => n1767, Q => 
                           REG_1_8_port);
   REG_reg_1_7_inst : DLH_X1 port map( G => n1843, D => n1773, Q => 
                           REG_1_7_port);
   REG_reg_1_6_inst : DLH_X1 port map( G => n1843, D => n1779, Q => 
                           REG_1_6_port);
   REG_reg_1_5_inst : DLH_X1 port map( G => n1843, D => n1785, Q => 
                           REG_1_5_port);
   REG_reg_1_4_inst : DLH_X1 port map( G => n1843, D => n1791, Q => 
                           REG_1_4_port);
   REG_reg_1_3_inst : DLH_X1 port map( G => n1843, D => n1797, Q => 
                           REG_1_3_port);
   REG_reg_1_2_inst : DLH_X1 port map( G => n1843, D => n1803, Q => 
                           REG_1_2_port);
   REG_reg_1_1_inst : DLH_X1 port map( G => n1843, D => n1809, Q => 
                           REG_1_1_port);
   REG_reg_1_0_inst : DLH_X1 port map( G => n1843, D => n1815, Q => 
                           REG_1_0_port);
   REG_reg_2_31_inst : DLH_X1 port map( G => n1853, D => n1629, Q => 
                           REG_2_31_port);
   REG_reg_2_30_inst : DLH_X1 port map( G => n1853, D => n1635, Q => 
                           REG_2_30_port);
   REG_reg_2_29_inst : DLH_X1 port map( G => n1852, D => n1641, Q => 
                           REG_2_29_port);
   REG_reg_2_28_inst : DLH_X1 port map( G => n1852, D => n1647, Q => 
                           REG_2_28_port);
   REG_reg_2_27_inst : DLH_X1 port map( G => n1852, D => n1653, Q => 
                           REG_2_27_port);
   REG_reg_2_26_inst : DLH_X1 port map( G => n1852, D => n1659, Q => 
                           REG_2_26_port);
   REG_reg_2_25_inst : DLH_X1 port map( G => n1852, D => n1665, Q => 
                           REG_2_25_port);
   REG_reg_2_24_inst : DLH_X1 port map( G => n1852, D => n1671, Q => 
                           REG_2_24_port);
   REG_reg_2_23_inst : DLH_X1 port map( G => n1852, D => n1677, Q => 
                           REG_2_23_port);
   REG_reg_2_22_inst : DLH_X1 port map( G => n1852, D => n1683, Q => 
                           REG_2_22_port);
   REG_reg_2_21_inst : DLH_X1 port map( G => n1852, D => n1689, Q => 
                           REG_2_21_port);
   REG_reg_2_20_inst : DLH_X1 port map( G => n1852, D => n1695, Q => 
                           REG_2_20_port);
   REG_reg_2_19_inst : DLH_X1 port map( G => n1851, D => n1701, Q => 
                           REG_2_19_port);
   REG_reg_2_18_inst : DLH_X1 port map( G => n1851, D => n1707, Q => 
                           REG_2_18_port);
   REG_reg_2_17_inst : DLH_X1 port map( G => n1851, D => n1713, Q => 
                           REG_2_17_port);
   REG_reg_2_16_inst : DLH_X1 port map( G => n1851, D => n1719, Q => 
                           REG_2_16_port);
   REG_reg_2_15_inst : DLH_X1 port map( G => n1851, D => n1725, Q => 
                           REG_2_15_port);
   REG_reg_2_14_inst : DLH_X1 port map( G => n1851, D => n1731, Q => 
                           REG_2_14_port);
   REG_reg_2_13_inst : DLH_X1 port map( G => n1851, D => n1737, Q => 
                           REG_2_13_port);
   REG_reg_2_12_inst : DLH_X1 port map( G => n1851, D => n1743, Q => 
                           REG_2_12_port);
   REG_reg_2_11_inst : DLH_X1 port map( G => n1851, D => n1749, Q => 
                           REG_2_11_port);
   REG_reg_2_10_inst : DLH_X1 port map( G => n1851, D => n1755, Q => 
                           REG_2_10_port);
   REG_reg_2_9_inst : DLH_X1 port map( G => n1850, D => n1761, Q => 
                           REG_2_9_port);
   REG_reg_2_8_inst : DLH_X1 port map( G => n1850, D => n1767, Q => 
                           REG_2_8_port);
   REG_reg_2_7_inst : DLH_X1 port map( G => n1850, D => n1773, Q => 
                           REG_2_7_port);
   REG_reg_2_6_inst : DLH_X1 port map( G => n1850, D => n1779, Q => 
                           REG_2_6_port);
   REG_reg_2_5_inst : DLH_X1 port map( G => n1850, D => n1785, Q => 
                           REG_2_5_port);
   REG_reg_2_4_inst : DLH_X1 port map( G => n1850, D => n1791, Q => 
                           REG_2_4_port);
   REG_reg_2_3_inst : DLH_X1 port map( G => n1850, D => n1797, Q => 
                           REG_2_3_port);
   REG_reg_2_2_inst : DLH_X1 port map( G => n1850, D => n1803, Q => 
                           REG_2_2_port);
   REG_reg_2_1_inst : DLH_X1 port map( G => n1850, D => n1809, Q => 
                           REG_2_1_port);
   REG_reg_2_0_inst : DLH_X1 port map( G => n1850, D => n1815, Q => 
                           REG_2_0_port);
   REG_reg_3_31_inst : DLH_X1 port map( G => n1860, D => n1629, Q => 
                           REG_3_31_port);
   REG_reg_3_30_inst : DLH_X1 port map( G => n1860, D => n1635, Q => 
                           REG_3_30_port);
   REG_reg_3_29_inst : DLH_X1 port map( G => n1859, D => n1641, Q => 
                           REG_3_29_port);
   REG_reg_3_28_inst : DLH_X1 port map( G => n1859, D => n1647, Q => 
                           REG_3_28_port);
   REG_reg_3_27_inst : DLH_X1 port map( G => n1859, D => n1653, Q => 
                           REG_3_27_port);
   REG_reg_3_26_inst : DLH_X1 port map( G => n1859, D => n1659, Q => 
                           REG_3_26_port);
   REG_reg_3_25_inst : DLH_X1 port map( G => n1859, D => n1665, Q => 
                           REG_3_25_port);
   REG_reg_3_24_inst : DLH_X1 port map( G => n1859, D => n1671, Q => 
                           REG_3_24_port);
   REG_reg_3_23_inst : DLH_X1 port map( G => n1859, D => n1677, Q => 
                           REG_3_23_port);
   REG_reg_3_22_inst : DLH_X1 port map( G => n1859, D => n1683, Q => 
                           REG_3_22_port);
   REG_reg_3_21_inst : DLH_X1 port map( G => n1859, D => n1689, Q => 
                           REG_3_21_port);
   REG_reg_3_20_inst : DLH_X1 port map( G => n1859, D => n1695, Q => 
                           REG_3_20_port);
   REG_reg_3_19_inst : DLH_X1 port map( G => n1858, D => n1701, Q => 
                           REG_3_19_port);
   REG_reg_3_18_inst : DLH_X1 port map( G => n1858, D => n1707, Q => 
                           REG_3_18_port);
   REG_reg_3_17_inst : DLH_X1 port map( G => n1858, D => n1713, Q => 
                           REG_3_17_port);
   REG_reg_3_16_inst : DLH_X1 port map( G => n1858, D => n1719, Q => 
                           REG_3_16_port);
   REG_reg_3_15_inst : DLH_X1 port map( G => n1858, D => n1725, Q => 
                           REG_3_15_port);
   REG_reg_3_14_inst : DLH_X1 port map( G => n1858, D => n1731, Q => 
                           REG_3_14_port);
   REG_reg_3_13_inst : DLH_X1 port map( G => n1858, D => n1737, Q => 
                           REG_3_13_port);
   REG_reg_3_12_inst : DLH_X1 port map( G => n1858, D => n1743, Q => 
                           REG_3_12_port);
   REG_reg_3_11_inst : DLH_X1 port map( G => n1858, D => n1749, Q => 
                           REG_3_11_port);
   REG_reg_3_10_inst : DLH_X1 port map( G => n1858, D => n1755, Q => 
                           REG_3_10_port);
   REG_reg_3_9_inst : DLH_X1 port map( G => n1857, D => n1761, Q => 
                           REG_3_9_port);
   REG_reg_3_8_inst : DLH_X1 port map( G => n1857, D => n1767, Q => 
                           REG_3_8_port);
   REG_reg_3_7_inst : DLH_X1 port map( G => n1857, D => n1773, Q => 
                           REG_3_7_port);
   REG_reg_3_6_inst : DLH_X1 port map( G => n1857, D => n1779, Q => 
                           REG_3_6_port);
   REG_reg_3_5_inst : DLH_X1 port map( G => n1857, D => n1785, Q => 
                           REG_3_5_port);
   REG_reg_3_4_inst : DLH_X1 port map( G => n1857, D => n1791, Q => 
                           REG_3_4_port);
   REG_reg_3_3_inst : DLH_X1 port map( G => n1857, D => n1797, Q => 
                           REG_3_3_port);
   REG_reg_3_2_inst : DLH_X1 port map( G => n1857, D => n1803, Q => 
                           REG_3_2_port);
   REG_reg_3_1_inst : DLH_X1 port map( G => n1857, D => n1809, Q => 
                           REG_3_1_port);
   REG_reg_3_0_inst : DLH_X1 port map( G => n1857, D => n1815, Q => 
                           REG_3_0_port);
   REG_reg_4_31_inst : DLH_X1 port map( G => n1867, D => n1629, Q => 
                           REG_4_31_port);
   REG_reg_4_30_inst : DLH_X1 port map( G => n1867, D => n1635, Q => 
                           REG_4_30_port);
   REG_reg_4_29_inst : DLH_X1 port map( G => n1866, D => n1641, Q => 
                           REG_4_29_port);
   REG_reg_4_28_inst : DLH_X1 port map( G => n1866, D => n1647, Q => 
                           REG_4_28_port);
   REG_reg_4_27_inst : DLH_X1 port map( G => n1866, D => n1653, Q => 
                           REG_4_27_port);
   REG_reg_4_26_inst : DLH_X1 port map( G => n1866, D => n1659, Q => 
                           REG_4_26_port);
   REG_reg_4_25_inst : DLH_X1 port map( G => n1866, D => n1665, Q => 
                           REG_4_25_port);
   REG_reg_4_24_inst : DLH_X1 port map( G => n1866, D => n1671, Q => 
                           REG_4_24_port);
   REG_reg_4_23_inst : DLH_X1 port map( G => n1866, D => n1677, Q => 
                           REG_4_23_port);
   REG_reg_4_22_inst : DLH_X1 port map( G => n1866, D => n1683, Q => 
                           REG_4_22_port);
   REG_reg_4_21_inst : DLH_X1 port map( G => n1866, D => n1689, Q => 
                           REG_4_21_port);
   REG_reg_4_20_inst : DLH_X1 port map( G => n1866, D => n1695, Q => 
                           REG_4_20_port);
   REG_reg_4_19_inst : DLH_X1 port map( G => n1865, D => n1701, Q => 
                           REG_4_19_port);
   REG_reg_4_18_inst : DLH_X1 port map( G => n1865, D => n1707, Q => 
                           REG_4_18_port);
   REG_reg_4_17_inst : DLH_X1 port map( G => n1865, D => n1713, Q => 
                           REG_4_17_port);
   REG_reg_4_16_inst : DLH_X1 port map( G => n1865, D => n1719, Q => 
                           REG_4_16_port);
   REG_reg_4_15_inst : DLH_X1 port map( G => n1865, D => n1725, Q => 
                           REG_4_15_port);
   REG_reg_4_14_inst : DLH_X1 port map( G => n1865, D => n1731, Q => 
                           REG_4_14_port);
   REG_reg_4_13_inst : DLH_X1 port map( G => n1865, D => n1737, Q => 
                           REG_4_13_port);
   REG_reg_4_12_inst : DLH_X1 port map( G => n1865, D => n1743, Q => 
                           REG_4_12_port);
   REG_reg_4_11_inst : DLH_X1 port map( G => n1865, D => n1749, Q => 
                           REG_4_11_port);
   REG_reg_4_10_inst : DLH_X1 port map( G => n1865, D => n1755, Q => 
                           REG_4_10_port);
   REG_reg_4_9_inst : DLH_X1 port map( G => n1864, D => n1761, Q => 
                           REG_4_9_port);
   REG_reg_4_8_inst : DLH_X1 port map( G => n1864, D => n1767, Q => 
                           REG_4_8_port);
   REG_reg_4_7_inst : DLH_X1 port map( G => n1864, D => n1773, Q => 
                           REG_4_7_port);
   REG_reg_4_6_inst : DLH_X1 port map( G => n1864, D => n1779, Q => 
                           REG_4_6_port);
   REG_reg_4_5_inst : DLH_X1 port map( G => n1864, D => n1785, Q => 
                           REG_4_5_port);
   REG_reg_4_4_inst : DLH_X1 port map( G => n1864, D => n1791, Q => 
                           REG_4_4_port);
   REG_reg_4_3_inst : DLH_X1 port map( G => n1864, D => n1797, Q => 
                           REG_4_3_port);
   REG_reg_4_2_inst : DLH_X1 port map( G => n1864, D => n1803, Q => 
                           REG_4_2_port);
   REG_reg_4_1_inst : DLH_X1 port map( G => n1864, D => n1809, Q => 
                           REG_4_1_port);
   REG_reg_4_0_inst : DLH_X1 port map( G => n1864, D => n1815, Q => 
                           REG_4_0_port);
   REG_reg_5_31_inst : DLH_X1 port map( G => n1874, D => n1629, Q => 
                           REG_5_31_port);
   REG_reg_5_30_inst : DLH_X1 port map( G => n1874, D => n1635, Q => 
                           REG_5_30_port);
   REG_reg_5_29_inst : DLH_X1 port map( G => n1873, D => n1641, Q => 
                           REG_5_29_port);
   REG_reg_5_28_inst : DLH_X1 port map( G => n1873, D => n1647, Q => 
                           REG_5_28_port);
   REG_reg_5_27_inst : DLH_X1 port map( G => n1873, D => n1653, Q => 
                           REG_5_27_port);
   REG_reg_5_26_inst : DLH_X1 port map( G => n1873, D => n1659, Q => 
                           REG_5_26_port);
   REG_reg_5_25_inst : DLH_X1 port map( G => n1873, D => n1665, Q => 
                           REG_5_25_port);
   REG_reg_5_24_inst : DLH_X1 port map( G => n1873, D => n1671, Q => 
                           REG_5_24_port);
   REG_reg_5_23_inst : DLH_X1 port map( G => n1873, D => n1677, Q => 
                           REG_5_23_port);
   REG_reg_5_22_inst : DLH_X1 port map( G => n1873, D => n1683, Q => 
                           REG_5_22_port);
   REG_reg_5_21_inst : DLH_X1 port map( G => n1873, D => n1689, Q => 
                           REG_5_21_port);
   REG_reg_5_20_inst : DLH_X1 port map( G => n1873, D => n1695, Q => 
                           REG_5_20_port);
   REG_reg_5_19_inst : DLH_X1 port map( G => n1872, D => n1701, Q => 
                           REG_5_19_port);
   REG_reg_5_18_inst : DLH_X1 port map( G => n1872, D => n1707, Q => 
                           REG_5_18_port);
   REG_reg_5_17_inst : DLH_X1 port map( G => n1872, D => n1713, Q => 
                           REG_5_17_port);
   REG_reg_5_16_inst : DLH_X1 port map( G => n1872, D => n1719, Q => 
                           REG_5_16_port);
   REG_reg_5_15_inst : DLH_X1 port map( G => n1872, D => n1725, Q => 
                           REG_5_15_port);
   REG_reg_5_14_inst : DLH_X1 port map( G => n1872, D => n1731, Q => 
                           REG_5_14_port);
   REG_reg_5_13_inst : DLH_X1 port map( G => n1872, D => n1737, Q => 
                           REG_5_13_port);
   REG_reg_5_12_inst : DLH_X1 port map( G => n1872, D => n1743, Q => 
                           REG_5_12_port);
   REG_reg_5_11_inst : DLH_X1 port map( G => n1872, D => n1749, Q => 
                           REG_5_11_port);
   REG_reg_5_10_inst : DLH_X1 port map( G => n1872, D => n1755, Q => 
                           REG_5_10_port);
   REG_reg_5_9_inst : DLH_X1 port map( G => n1871, D => n1761, Q => 
                           REG_5_9_port);
   REG_reg_5_8_inst : DLH_X1 port map( G => n1871, D => n1767, Q => 
                           REG_5_8_port);
   REG_reg_5_7_inst : DLH_X1 port map( G => n1871, D => n1773, Q => 
                           REG_5_7_port);
   REG_reg_5_6_inst : DLH_X1 port map( G => n1871, D => n1779, Q => 
                           REG_5_6_port);
   REG_reg_5_5_inst : DLH_X1 port map( G => n1871, D => n1785, Q => 
                           REG_5_5_port);
   REG_reg_5_4_inst : DLH_X1 port map( G => n1871, D => n1791, Q => 
                           REG_5_4_port);
   REG_reg_5_3_inst : DLH_X1 port map( G => n1871, D => n1797, Q => 
                           REG_5_3_port);
   REG_reg_5_2_inst : DLH_X1 port map( G => n1871, D => n1803, Q => 
                           REG_5_2_port);
   REG_reg_5_1_inst : DLH_X1 port map( G => n1871, D => n1809, Q => 
                           REG_5_1_port);
   REG_reg_5_0_inst : DLH_X1 port map( G => n1871, D => n1815, Q => 
                           REG_5_0_port);
   REG_reg_6_31_inst : DLH_X1 port map( G => n1881, D => n1629, Q => 
                           REG_6_31_port);
   REG_reg_6_30_inst : DLH_X1 port map( G => n1881, D => n1635, Q => 
                           REG_6_30_port);
   REG_reg_6_29_inst : DLH_X1 port map( G => n1880, D => n1641, Q => 
                           REG_6_29_port);
   REG_reg_6_28_inst : DLH_X1 port map( G => n1880, D => n1647, Q => 
                           REG_6_28_port);
   REG_reg_6_27_inst : DLH_X1 port map( G => n1880, D => n1653, Q => 
                           REG_6_27_port);
   REG_reg_6_26_inst : DLH_X1 port map( G => n1880, D => n1659, Q => 
                           REG_6_26_port);
   REG_reg_6_25_inst : DLH_X1 port map( G => n1880, D => n1665, Q => 
                           REG_6_25_port);
   REG_reg_6_24_inst : DLH_X1 port map( G => n1880, D => n1671, Q => 
                           REG_6_24_port);
   REG_reg_6_23_inst : DLH_X1 port map( G => n1880, D => n1677, Q => 
                           REG_6_23_port);
   REG_reg_6_22_inst : DLH_X1 port map( G => n1880, D => n1683, Q => 
                           REG_6_22_port);
   REG_reg_6_21_inst : DLH_X1 port map( G => n1880, D => n1689, Q => 
                           REG_6_21_port);
   REG_reg_6_20_inst : DLH_X1 port map( G => n1880, D => n1695, Q => 
                           REG_6_20_port);
   REG_reg_6_19_inst : DLH_X1 port map( G => n1879, D => n1701, Q => 
                           REG_6_19_port);
   REG_reg_6_18_inst : DLH_X1 port map( G => n1879, D => n1707, Q => 
                           REG_6_18_port);
   REG_reg_6_17_inst : DLH_X1 port map( G => n1879, D => n1713, Q => 
                           REG_6_17_port);
   REG_reg_6_16_inst : DLH_X1 port map( G => n1879, D => n1719, Q => 
                           REG_6_16_port);
   REG_reg_6_15_inst : DLH_X1 port map( G => n1879, D => n1725, Q => 
                           REG_6_15_port);
   REG_reg_6_14_inst : DLH_X1 port map( G => n1879, D => n1731, Q => 
                           REG_6_14_port);
   REG_reg_6_13_inst : DLH_X1 port map( G => n1879, D => n1737, Q => 
                           REG_6_13_port);
   REG_reg_6_12_inst : DLH_X1 port map( G => n1879, D => n1743, Q => 
                           REG_6_12_port);
   REG_reg_6_11_inst : DLH_X1 port map( G => n1879, D => n1749, Q => 
                           REG_6_11_port);
   REG_reg_6_10_inst : DLH_X1 port map( G => n1879, D => n1755, Q => 
                           REG_6_10_port);
   REG_reg_6_9_inst : DLH_X1 port map( G => n1878, D => n1761, Q => 
                           REG_6_9_port);
   REG_reg_6_8_inst : DLH_X1 port map( G => n1878, D => n1767, Q => 
                           REG_6_8_port);
   REG_reg_6_7_inst : DLH_X1 port map( G => n1878, D => n1773, Q => 
                           REG_6_7_port);
   REG_reg_6_6_inst : DLH_X1 port map( G => n1878, D => n1779, Q => 
                           REG_6_6_port);
   REG_reg_6_5_inst : DLH_X1 port map( G => n1878, D => n1785, Q => 
                           REG_6_5_port);
   REG_reg_6_4_inst : DLH_X1 port map( G => n1878, D => n1791, Q => 
                           REG_6_4_port);
   REG_reg_6_3_inst : DLH_X1 port map( G => n1878, D => n1797, Q => 
                           REG_6_3_port);
   REG_reg_6_2_inst : DLH_X1 port map( G => n1878, D => n1803, Q => 
                           REG_6_2_port);
   REG_reg_6_1_inst : DLH_X1 port map( G => n1878, D => n1809, Q => 
                           REG_6_1_port);
   REG_reg_6_0_inst : DLH_X1 port map( G => n1878, D => n1815, Q => 
                           REG_6_0_port);
   REG_reg_7_31_inst : DLH_X1 port map( G => n1888, D => n1629, Q => 
                           REG_7_31_port);
   REG_reg_7_30_inst : DLH_X1 port map( G => n1888, D => n1635, Q => 
                           REG_7_30_port);
   REG_reg_7_29_inst : DLH_X1 port map( G => n1887, D => n1641, Q => 
                           REG_7_29_port);
   REG_reg_7_28_inst : DLH_X1 port map( G => n1887, D => n1647, Q => 
                           REG_7_28_port);
   REG_reg_7_27_inst : DLH_X1 port map( G => n1887, D => n1653, Q => 
                           REG_7_27_port);
   REG_reg_7_26_inst : DLH_X1 port map( G => n1887, D => n1659, Q => 
                           REG_7_26_port);
   REG_reg_7_25_inst : DLH_X1 port map( G => n1887, D => n1665, Q => 
                           REG_7_25_port);
   REG_reg_7_24_inst : DLH_X1 port map( G => n1887, D => n1671, Q => 
                           REG_7_24_port);
   REG_reg_7_23_inst : DLH_X1 port map( G => n1887, D => n1677, Q => 
                           REG_7_23_port);
   REG_reg_7_22_inst : DLH_X1 port map( G => n1887, D => n1683, Q => 
                           REG_7_22_port);
   REG_reg_7_21_inst : DLH_X1 port map( G => n1887, D => n1689, Q => 
                           REG_7_21_port);
   REG_reg_7_20_inst : DLH_X1 port map( G => n1887, D => n1695, Q => 
                           REG_7_20_port);
   REG_reg_7_19_inst : DLH_X1 port map( G => n1886, D => n1701, Q => 
                           REG_7_19_port);
   REG_reg_7_18_inst : DLH_X1 port map( G => n1886, D => n1707, Q => 
                           REG_7_18_port);
   REG_reg_7_17_inst : DLH_X1 port map( G => n1886, D => n1713, Q => 
                           REG_7_17_port);
   REG_reg_7_16_inst : DLH_X1 port map( G => n1886, D => n1719, Q => 
                           REG_7_16_port);
   REG_reg_7_15_inst : DLH_X1 port map( G => n1886, D => n1725, Q => 
                           REG_7_15_port);
   REG_reg_7_14_inst : DLH_X1 port map( G => n1886, D => n1731, Q => 
                           REG_7_14_port);
   REG_reg_7_13_inst : DLH_X1 port map( G => n1886, D => n1737, Q => 
                           REG_7_13_port);
   REG_reg_7_12_inst : DLH_X1 port map( G => n1886, D => n1743, Q => 
                           REG_7_12_port);
   REG_reg_7_11_inst : DLH_X1 port map( G => n1886, D => n1749, Q => 
                           REG_7_11_port);
   REG_reg_7_10_inst : DLH_X1 port map( G => n1886, D => n1755, Q => 
                           REG_7_10_port);
   REG_reg_7_9_inst : DLH_X1 port map( G => n1885, D => n1761, Q => 
                           REG_7_9_port);
   REG_reg_7_8_inst : DLH_X1 port map( G => n1885, D => n1767, Q => 
                           REG_7_8_port);
   REG_reg_7_7_inst : DLH_X1 port map( G => n1885, D => n1773, Q => 
                           REG_7_7_port);
   REG_reg_7_6_inst : DLH_X1 port map( G => n1885, D => n1779, Q => 
                           REG_7_6_port);
   REG_reg_7_5_inst : DLH_X1 port map( G => n1885, D => n1785, Q => 
                           REG_7_5_port);
   REG_reg_7_4_inst : DLH_X1 port map( G => n1885, D => n1791, Q => 
                           REG_7_4_port);
   REG_reg_7_3_inst : DLH_X1 port map( G => n1885, D => n1797, Q => 
                           REG_7_3_port);
   REG_reg_7_2_inst : DLH_X1 port map( G => n1885, D => n1803, Q => 
                           REG_7_2_port);
   REG_reg_7_1_inst : DLH_X1 port map( G => n1885, D => n1809, Q => 
                           REG_7_1_port);
   REG_reg_7_0_inst : DLH_X1 port map( G => n1885, D => n1815, Q => 
                           REG_7_0_port);
   REG_reg_8_31_inst : DLH_X1 port map( G => n1895, D => n1629, Q => 
                           REG_8_31_port);
   REG_reg_8_30_inst : DLH_X1 port map( G => n1895, D => n1635, Q => 
                           REG_8_30_port);
   REG_reg_8_29_inst : DLH_X1 port map( G => n1894, D => n1641, Q => 
                           REG_8_29_port);
   REG_reg_8_28_inst : DLH_X1 port map( G => n1894, D => n1647, Q => 
                           REG_8_28_port);
   REG_reg_8_27_inst : DLH_X1 port map( G => n1894, D => n1653, Q => 
                           REG_8_27_port);
   REG_reg_8_26_inst : DLH_X1 port map( G => n1894, D => n1659, Q => 
                           REG_8_26_port);
   REG_reg_8_25_inst : DLH_X1 port map( G => n1894, D => n1665, Q => 
                           REG_8_25_port);
   REG_reg_8_24_inst : DLH_X1 port map( G => n1894, D => n1671, Q => 
                           REG_8_24_port);
   REG_reg_8_23_inst : DLH_X1 port map( G => n1894, D => n1677, Q => 
                           REG_8_23_port);
   REG_reg_8_22_inst : DLH_X1 port map( G => n1894, D => n1683, Q => 
                           REG_8_22_port);
   REG_reg_8_21_inst : DLH_X1 port map( G => n1894, D => n1689, Q => 
                           REG_8_21_port);
   REG_reg_8_20_inst : DLH_X1 port map( G => n1894, D => n1695, Q => 
                           REG_8_20_port);
   REG_reg_8_19_inst : DLH_X1 port map( G => n1893, D => n1701, Q => 
                           REG_8_19_port);
   REG_reg_8_18_inst : DLH_X1 port map( G => n1893, D => n1707, Q => 
                           REG_8_18_port);
   REG_reg_8_17_inst : DLH_X1 port map( G => n1893, D => n1713, Q => 
                           REG_8_17_port);
   REG_reg_8_16_inst : DLH_X1 port map( G => n1893, D => n1719, Q => 
                           REG_8_16_port);
   REG_reg_8_15_inst : DLH_X1 port map( G => n1893, D => n1725, Q => 
                           REG_8_15_port);
   REG_reg_8_14_inst : DLH_X1 port map( G => n1893, D => n1731, Q => 
                           REG_8_14_port);
   REG_reg_8_13_inst : DLH_X1 port map( G => n1893, D => n1737, Q => 
                           REG_8_13_port);
   REG_reg_8_12_inst : DLH_X1 port map( G => n1893, D => n1743, Q => 
                           REG_8_12_port);
   REG_reg_8_11_inst : DLH_X1 port map( G => n1893, D => n1749, Q => 
                           REG_8_11_port);
   REG_reg_8_10_inst : DLH_X1 port map( G => n1893, D => n1755, Q => 
                           REG_8_10_port);
   REG_reg_8_9_inst : DLH_X1 port map( G => n1892, D => n1761, Q => 
                           REG_8_9_port);
   REG_reg_8_8_inst : DLH_X1 port map( G => n1892, D => n1767, Q => 
                           REG_8_8_port);
   REG_reg_8_7_inst : DLH_X1 port map( G => n1892, D => n1773, Q => 
                           REG_8_7_port);
   REG_reg_8_6_inst : DLH_X1 port map( G => n1892, D => n1779, Q => 
                           REG_8_6_port);
   REG_reg_8_5_inst : DLH_X1 port map( G => n1892, D => n1785, Q => 
                           REG_8_5_port);
   REG_reg_8_4_inst : DLH_X1 port map( G => n1892, D => n1791, Q => 
                           REG_8_4_port);
   REG_reg_8_3_inst : DLH_X1 port map( G => n1892, D => n1797, Q => 
                           REG_8_3_port);
   REG_reg_8_2_inst : DLH_X1 port map( G => n1892, D => n1803, Q => 
                           REG_8_2_port);
   REG_reg_8_1_inst : DLH_X1 port map( G => n1892, D => n1809, Q => 
                           REG_8_1_port);
   REG_reg_8_0_inst : DLH_X1 port map( G => n1892, D => n1815, Q => 
                           REG_8_0_port);
   REG_reg_9_31_inst : DLH_X1 port map( G => n1902, D => n1629, Q => 
                           REG_9_31_port);
   REG_reg_9_30_inst : DLH_X1 port map( G => n1902, D => n1635, Q => 
                           REG_9_30_port);
   REG_reg_9_29_inst : DLH_X1 port map( G => n1901, D => n1641, Q => 
                           REG_9_29_port);
   REG_reg_9_28_inst : DLH_X1 port map( G => n1901, D => n1647, Q => 
                           REG_9_28_port);
   REG_reg_9_27_inst : DLH_X1 port map( G => n1901, D => n1653, Q => 
                           REG_9_27_port);
   REG_reg_9_26_inst : DLH_X1 port map( G => n1901, D => n1659, Q => 
                           REG_9_26_port);
   REG_reg_9_25_inst : DLH_X1 port map( G => n1901, D => n1665, Q => 
                           REG_9_25_port);
   REG_reg_9_24_inst : DLH_X1 port map( G => n1901, D => n1671, Q => 
                           REG_9_24_port);
   REG_reg_9_23_inst : DLH_X1 port map( G => n1901, D => n1677, Q => 
                           REG_9_23_port);
   REG_reg_9_22_inst : DLH_X1 port map( G => n1901, D => n1683, Q => 
                           REG_9_22_port);
   REG_reg_9_21_inst : DLH_X1 port map( G => n1901, D => n1689, Q => 
                           REG_9_21_port);
   REG_reg_9_20_inst : DLH_X1 port map( G => n1901, D => n1695, Q => 
                           REG_9_20_port);
   REG_reg_9_19_inst : DLH_X1 port map( G => n1900, D => n1701, Q => 
                           REG_9_19_port);
   REG_reg_9_18_inst : DLH_X1 port map( G => n1900, D => n1707, Q => 
                           REG_9_18_port);
   REG_reg_9_17_inst : DLH_X1 port map( G => n1900, D => n1713, Q => 
                           REG_9_17_port);
   REG_reg_9_16_inst : DLH_X1 port map( G => n1900, D => n1719, Q => 
                           REG_9_16_port);
   REG_reg_9_15_inst : DLH_X1 port map( G => n1900, D => n1725, Q => 
                           REG_9_15_port);
   REG_reg_9_14_inst : DLH_X1 port map( G => n1900, D => n1731, Q => 
                           REG_9_14_port);
   REG_reg_9_13_inst : DLH_X1 port map( G => n1900, D => n1737, Q => 
                           REG_9_13_port);
   REG_reg_9_12_inst : DLH_X1 port map( G => n1900, D => n1743, Q => 
                           REG_9_12_port);
   REG_reg_9_11_inst : DLH_X1 port map( G => n1900, D => n1749, Q => 
                           REG_9_11_port);
   REG_reg_9_10_inst : DLH_X1 port map( G => n1900, D => n1755, Q => 
                           REG_9_10_port);
   REG_reg_9_9_inst : DLH_X1 port map( G => n1899, D => n1761, Q => 
                           REG_9_9_port);
   REG_reg_9_8_inst : DLH_X1 port map( G => n1899, D => n1767, Q => 
                           REG_9_8_port);
   REG_reg_9_7_inst : DLH_X1 port map( G => n1899, D => n1773, Q => 
                           REG_9_7_port);
   REG_reg_9_6_inst : DLH_X1 port map( G => n1899, D => n1779, Q => 
                           REG_9_6_port);
   REG_reg_9_5_inst : DLH_X1 port map( G => n1899, D => n1785, Q => 
                           REG_9_5_port);
   REG_reg_9_4_inst : DLH_X1 port map( G => n1899, D => n1791, Q => 
                           REG_9_4_port);
   REG_reg_9_3_inst : DLH_X1 port map( G => n1899, D => n1797, Q => 
                           REG_9_3_port);
   REG_reg_9_2_inst : DLH_X1 port map( G => n1899, D => n1803, Q => 
                           REG_9_2_port);
   REG_reg_9_1_inst : DLH_X1 port map( G => n1899, D => n1809, Q => 
                           REG_9_1_port);
   REG_reg_9_0_inst : DLH_X1 port map( G => n1899, D => n1815, Q => 
                           REG_9_0_port);
   REG_reg_10_31_inst : DLH_X1 port map( G => n1909, D => n1629, Q => 
                           REG_10_31_port);
   REG_reg_10_30_inst : DLH_X1 port map( G => n1909, D => n1635, Q => 
                           REG_10_30_port);
   REG_reg_10_29_inst : DLH_X1 port map( G => n1908, D => n1641, Q => 
                           REG_10_29_port);
   REG_reg_10_28_inst : DLH_X1 port map( G => n1908, D => n1647, Q => 
                           REG_10_28_port);
   REG_reg_10_27_inst : DLH_X1 port map( G => n1908, D => n1653, Q => 
                           REG_10_27_port);
   REG_reg_10_26_inst : DLH_X1 port map( G => n1908, D => n1659, Q => 
                           REG_10_26_port);
   REG_reg_10_25_inst : DLH_X1 port map( G => n1908, D => n1665, Q => 
                           REG_10_25_port);
   REG_reg_10_24_inst : DLH_X1 port map( G => n1908, D => n1671, Q => 
                           REG_10_24_port);
   REG_reg_10_23_inst : DLH_X1 port map( G => n1908, D => n1677, Q => 
                           REG_10_23_port);
   REG_reg_10_22_inst : DLH_X1 port map( G => n1908, D => n1683, Q => 
                           REG_10_22_port);
   REG_reg_10_21_inst : DLH_X1 port map( G => n1908, D => n1689, Q => 
                           REG_10_21_port);
   REG_reg_10_20_inst : DLH_X1 port map( G => n1908, D => n1695, Q => 
                           REG_10_20_port);
   REG_reg_10_19_inst : DLH_X1 port map( G => n1907, D => n1701, Q => 
                           REG_10_19_port);
   REG_reg_10_18_inst : DLH_X1 port map( G => n1907, D => n1707, Q => 
                           REG_10_18_port);
   REG_reg_10_17_inst : DLH_X1 port map( G => n1907, D => n1713, Q => 
                           REG_10_17_port);
   REG_reg_10_16_inst : DLH_X1 port map( G => n1907, D => n1719, Q => 
                           REG_10_16_port);
   REG_reg_10_15_inst : DLH_X1 port map( G => n1907, D => n1725, Q => 
                           REG_10_15_port);
   REG_reg_10_14_inst : DLH_X1 port map( G => n1907, D => n1731, Q => 
                           REG_10_14_port);
   REG_reg_10_13_inst : DLH_X1 port map( G => n1907, D => n1737, Q => 
                           REG_10_13_port);
   REG_reg_10_12_inst : DLH_X1 port map( G => n1907, D => n1743, Q => 
                           REG_10_12_port);
   REG_reg_10_11_inst : DLH_X1 port map( G => n1907, D => n1749, Q => 
                           REG_10_11_port);
   REG_reg_10_10_inst : DLH_X1 port map( G => n1907, D => n1755, Q => 
                           REG_10_10_port);
   REG_reg_10_9_inst : DLH_X1 port map( G => n1906, D => n1761, Q => 
                           REG_10_9_port);
   REG_reg_10_8_inst : DLH_X1 port map( G => n1906, D => n1767, Q => 
                           REG_10_8_port);
   REG_reg_10_7_inst : DLH_X1 port map( G => n1906, D => n1773, Q => 
                           REG_10_7_port);
   REG_reg_10_6_inst : DLH_X1 port map( G => n1906, D => n1779, Q => 
                           REG_10_6_port);
   REG_reg_10_5_inst : DLH_X1 port map( G => n1906, D => n1785, Q => 
                           REG_10_5_port);
   REG_reg_10_4_inst : DLH_X1 port map( G => n1906, D => n1791, Q => 
                           REG_10_4_port);
   REG_reg_10_3_inst : DLH_X1 port map( G => n1906, D => n1797, Q => 
                           REG_10_3_port);
   REG_reg_10_2_inst : DLH_X1 port map( G => n1906, D => n1803, Q => 
                           REG_10_2_port);
   REG_reg_10_1_inst : DLH_X1 port map( G => n1906, D => n1809, Q => 
                           REG_10_1_port);
   REG_reg_10_0_inst : DLH_X1 port map( G => n1906, D => n1815, Q => 
                           REG_10_0_port);
   REG_reg_11_31_inst : DLH_X1 port map( G => n1916, D => n1630, Q => 
                           REG_11_31_port);
   REG_reg_11_30_inst : DLH_X1 port map( G => n1916, D => n1636, Q => 
                           REG_11_30_port);
   REG_reg_11_29_inst : DLH_X1 port map( G => n1915, D => n1642, Q => 
                           REG_11_29_port);
   REG_reg_11_28_inst : DLH_X1 port map( G => n1915, D => n1648, Q => 
                           REG_11_28_port);
   REG_reg_11_27_inst : DLH_X1 port map( G => n1915, D => n1654, Q => 
                           REG_11_27_port);
   REG_reg_11_26_inst : DLH_X1 port map( G => n1915, D => n1660, Q => 
                           REG_11_26_port);
   REG_reg_11_25_inst : DLH_X1 port map( G => n1915, D => n1666, Q => 
                           REG_11_25_port);
   REG_reg_11_24_inst : DLH_X1 port map( G => n1915, D => n1672, Q => 
                           REG_11_24_port);
   REG_reg_11_23_inst : DLH_X1 port map( G => n1915, D => n1678, Q => 
                           REG_11_23_port);
   REG_reg_11_22_inst : DLH_X1 port map( G => n1915, D => n1684, Q => 
                           REG_11_22_port);
   REG_reg_11_21_inst : DLH_X1 port map( G => n1915, D => n1690, Q => 
                           REG_11_21_port);
   REG_reg_11_20_inst : DLH_X1 port map( G => n1915, D => n1696, Q => 
                           REG_11_20_port);
   REG_reg_11_19_inst : DLH_X1 port map( G => n1914, D => n1702, Q => 
                           REG_11_19_port);
   REG_reg_11_18_inst : DLH_X1 port map( G => n1914, D => n1708, Q => 
                           REG_11_18_port);
   REG_reg_11_17_inst : DLH_X1 port map( G => n1914, D => n1714, Q => 
                           REG_11_17_port);
   REG_reg_11_16_inst : DLH_X1 port map( G => n1914, D => n1720, Q => 
                           REG_11_16_port);
   REG_reg_11_15_inst : DLH_X1 port map( G => n1914, D => n1726, Q => 
                           REG_11_15_port);
   REG_reg_11_14_inst : DLH_X1 port map( G => n1914, D => n1732, Q => 
                           REG_11_14_port);
   REG_reg_11_13_inst : DLH_X1 port map( G => n1914, D => n1738, Q => 
                           REG_11_13_port);
   REG_reg_11_12_inst : DLH_X1 port map( G => n1914, D => n1744, Q => 
                           REG_11_12_port);
   REG_reg_11_11_inst : DLH_X1 port map( G => n1914, D => n1750, Q => 
                           REG_11_11_port);
   REG_reg_11_10_inst : DLH_X1 port map( G => n1914, D => n1756, Q => 
                           REG_11_10_port);
   REG_reg_11_9_inst : DLH_X1 port map( G => n1913, D => n1762, Q => 
                           REG_11_9_port);
   REG_reg_11_8_inst : DLH_X1 port map( G => n1913, D => n1768, Q => 
                           REG_11_8_port);
   REG_reg_11_7_inst : DLH_X1 port map( G => n1913, D => n1774, Q => 
                           REG_11_7_port);
   REG_reg_11_6_inst : DLH_X1 port map( G => n1913, D => n1780, Q => 
                           REG_11_6_port);
   REG_reg_11_5_inst : DLH_X1 port map( G => n1913, D => n1786, Q => 
                           REG_11_5_port);
   REG_reg_11_4_inst : DLH_X1 port map( G => n1913, D => n1792, Q => 
                           REG_11_4_port);
   REG_reg_11_3_inst : DLH_X1 port map( G => n1913, D => n1798, Q => 
                           REG_11_3_port);
   REG_reg_11_2_inst : DLH_X1 port map( G => n1913, D => n1804, Q => 
                           REG_11_2_port);
   REG_reg_11_1_inst : DLH_X1 port map( G => n1913, D => n1810, Q => 
                           REG_11_1_port);
   REG_reg_11_0_inst : DLH_X1 port map( G => n1913, D => n1816, Q => 
                           REG_11_0_port);
   REG_reg_12_31_inst : DLH_X1 port map( G => n1923, D => n1630, Q => 
                           REG_12_31_port);
   REG_reg_12_30_inst : DLH_X1 port map( G => n1923, D => n1636, Q => 
                           REG_12_30_port);
   REG_reg_12_29_inst : DLH_X1 port map( G => n1922, D => n1642, Q => 
                           REG_12_29_port);
   REG_reg_12_28_inst : DLH_X1 port map( G => n1922, D => n1648, Q => 
                           REG_12_28_port);
   REG_reg_12_27_inst : DLH_X1 port map( G => n1922, D => n1654, Q => 
                           REG_12_27_port);
   REG_reg_12_26_inst : DLH_X1 port map( G => n1922, D => n1660, Q => 
                           REG_12_26_port);
   REG_reg_12_25_inst : DLH_X1 port map( G => n1922, D => n1666, Q => 
                           REG_12_25_port);
   REG_reg_12_24_inst : DLH_X1 port map( G => n1922, D => n1672, Q => 
                           REG_12_24_port);
   REG_reg_12_23_inst : DLH_X1 port map( G => n1922, D => n1678, Q => 
                           REG_12_23_port);
   REG_reg_12_22_inst : DLH_X1 port map( G => n1922, D => n1684, Q => 
                           REG_12_22_port);
   REG_reg_12_21_inst : DLH_X1 port map( G => n1922, D => n1690, Q => 
                           REG_12_21_port);
   REG_reg_12_20_inst : DLH_X1 port map( G => n1922, D => n1696, Q => 
                           REG_12_20_port);
   REG_reg_12_19_inst : DLH_X1 port map( G => n1921, D => n1702, Q => 
                           REG_12_19_port);
   REG_reg_12_18_inst : DLH_X1 port map( G => n1921, D => n1708, Q => 
                           REG_12_18_port);
   REG_reg_12_17_inst : DLH_X1 port map( G => n1921, D => n1714, Q => 
                           REG_12_17_port);
   REG_reg_12_16_inst : DLH_X1 port map( G => n1921, D => n1720, Q => 
                           REG_12_16_port);
   REG_reg_12_15_inst : DLH_X1 port map( G => n1921, D => n1726, Q => 
                           REG_12_15_port);
   REG_reg_12_14_inst : DLH_X1 port map( G => n1921, D => n1732, Q => 
                           REG_12_14_port);
   REG_reg_12_13_inst : DLH_X1 port map( G => n1921, D => n1738, Q => 
                           REG_12_13_port);
   REG_reg_12_12_inst : DLH_X1 port map( G => n1921, D => n1744, Q => 
                           REG_12_12_port);
   REG_reg_12_11_inst : DLH_X1 port map( G => n1921, D => n1750, Q => 
                           REG_12_11_port);
   REG_reg_12_10_inst : DLH_X1 port map( G => n1921, D => n1756, Q => 
                           REG_12_10_port);
   REG_reg_12_9_inst : DLH_X1 port map( G => n1920, D => n1762, Q => 
                           REG_12_9_port);
   REG_reg_12_8_inst : DLH_X1 port map( G => n1920, D => n1768, Q => 
                           REG_12_8_port);
   REG_reg_12_7_inst : DLH_X1 port map( G => n1920, D => n1774, Q => 
                           REG_12_7_port);
   REG_reg_12_6_inst : DLH_X1 port map( G => n1920, D => n1780, Q => 
                           REG_12_6_port);
   REG_reg_12_5_inst : DLH_X1 port map( G => n1920, D => n1786, Q => 
                           REG_12_5_port);
   REG_reg_12_4_inst : DLH_X1 port map( G => n1920, D => n1792, Q => 
                           REG_12_4_port);
   REG_reg_12_3_inst : DLH_X1 port map( G => n1920, D => n1798, Q => 
                           REG_12_3_port);
   REG_reg_12_2_inst : DLH_X1 port map( G => n1920, D => n1804, Q => 
                           REG_12_2_port);
   REG_reg_12_1_inst : DLH_X1 port map( G => n1920, D => n1810, Q => 
                           REG_12_1_port);
   REG_reg_12_0_inst : DLH_X1 port map( G => n1920, D => n1816, Q => 
                           REG_12_0_port);
   REG_reg_13_31_inst : DLH_X1 port map( G => n1930, D => n1630, Q => 
                           REG_13_31_port);
   REG_reg_13_30_inst : DLH_X1 port map( G => n1930, D => n1636, Q => 
                           REG_13_30_port);
   REG_reg_13_29_inst : DLH_X1 port map( G => n1929, D => n1642, Q => 
                           REG_13_29_port);
   REG_reg_13_28_inst : DLH_X1 port map( G => n1929, D => n1648, Q => 
                           REG_13_28_port);
   REG_reg_13_27_inst : DLH_X1 port map( G => n1929, D => n1654, Q => 
                           REG_13_27_port);
   REG_reg_13_26_inst : DLH_X1 port map( G => n1929, D => n1660, Q => 
                           REG_13_26_port);
   REG_reg_13_25_inst : DLH_X1 port map( G => n1929, D => n1666, Q => 
                           REG_13_25_port);
   REG_reg_13_24_inst : DLH_X1 port map( G => n1929, D => n1672, Q => 
                           REG_13_24_port);
   REG_reg_13_23_inst : DLH_X1 port map( G => n1929, D => n1678, Q => 
                           REG_13_23_port);
   REG_reg_13_22_inst : DLH_X1 port map( G => n1929, D => n1684, Q => 
                           REG_13_22_port);
   REG_reg_13_21_inst : DLH_X1 port map( G => n1929, D => n1690, Q => 
                           REG_13_21_port);
   REG_reg_13_20_inst : DLH_X1 port map( G => n1929, D => n1696, Q => 
                           REG_13_20_port);
   REG_reg_13_19_inst : DLH_X1 port map( G => n1928, D => n1702, Q => 
                           REG_13_19_port);
   REG_reg_13_18_inst : DLH_X1 port map( G => n1928, D => n1708, Q => 
                           REG_13_18_port);
   REG_reg_13_17_inst : DLH_X1 port map( G => n1928, D => n1714, Q => 
                           REG_13_17_port);
   REG_reg_13_16_inst : DLH_X1 port map( G => n1928, D => n1720, Q => 
                           REG_13_16_port);
   REG_reg_13_15_inst : DLH_X1 port map( G => n1928, D => n1726, Q => 
                           REG_13_15_port);
   REG_reg_13_14_inst : DLH_X1 port map( G => n1928, D => n1732, Q => 
                           REG_13_14_port);
   REG_reg_13_13_inst : DLH_X1 port map( G => n1928, D => n1738, Q => 
                           REG_13_13_port);
   REG_reg_13_12_inst : DLH_X1 port map( G => n1928, D => n1744, Q => 
                           REG_13_12_port);
   REG_reg_13_11_inst : DLH_X1 port map( G => n1928, D => n1750, Q => 
                           REG_13_11_port);
   REG_reg_13_10_inst : DLH_X1 port map( G => n1928, D => n1756, Q => 
                           REG_13_10_port);
   REG_reg_13_9_inst : DLH_X1 port map( G => n1927, D => n1762, Q => 
                           REG_13_9_port);
   REG_reg_13_8_inst : DLH_X1 port map( G => n1927, D => n1768, Q => 
                           REG_13_8_port);
   REG_reg_13_7_inst : DLH_X1 port map( G => n1927, D => n1774, Q => 
                           REG_13_7_port);
   REG_reg_13_6_inst : DLH_X1 port map( G => n1927, D => n1780, Q => 
                           REG_13_6_port);
   REG_reg_13_5_inst : DLH_X1 port map( G => n1927, D => n1786, Q => 
                           REG_13_5_port);
   REG_reg_13_4_inst : DLH_X1 port map( G => n1927, D => n1792, Q => 
                           REG_13_4_port);
   REG_reg_13_3_inst : DLH_X1 port map( G => n1927, D => n1798, Q => 
                           REG_13_3_port);
   REG_reg_13_2_inst : DLH_X1 port map( G => n1927, D => n1804, Q => 
                           REG_13_2_port);
   REG_reg_13_1_inst : DLH_X1 port map( G => n1927, D => n1810, Q => 
                           REG_13_1_port);
   REG_reg_13_0_inst : DLH_X1 port map( G => n1927, D => n1816, Q => 
                           REG_13_0_port);
   REG_reg_14_31_inst : DLH_X1 port map( G => n1937, D => n1630, Q => 
                           REG_14_31_port);
   REG_reg_14_30_inst : DLH_X1 port map( G => n1937, D => n1636, Q => 
                           REG_14_30_port);
   REG_reg_14_29_inst : DLH_X1 port map( G => n1936, D => n1642, Q => 
                           REG_14_29_port);
   REG_reg_14_28_inst : DLH_X1 port map( G => n1936, D => n1648, Q => 
                           REG_14_28_port);
   REG_reg_14_27_inst : DLH_X1 port map( G => n1936, D => n1654, Q => 
                           REG_14_27_port);
   REG_reg_14_26_inst : DLH_X1 port map( G => n1936, D => n1660, Q => 
                           REG_14_26_port);
   REG_reg_14_25_inst : DLH_X1 port map( G => n1936, D => n1666, Q => 
                           REG_14_25_port);
   REG_reg_14_24_inst : DLH_X1 port map( G => n1936, D => n1672, Q => 
                           REG_14_24_port);
   REG_reg_14_23_inst : DLH_X1 port map( G => n1936, D => n1678, Q => 
                           REG_14_23_port);
   REG_reg_14_22_inst : DLH_X1 port map( G => n1936, D => n1684, Q => 
                           REG_14_22_port);
   REG_reg_14_21_inst : DLH_X1 port map( G => n1936, D => n1690, Q => 
                           REG_14_21_port);
   REG_reg_14_20_inst : DLH_X1 port map( G => n1936, D => n1696, Q => 
                           REG_14_20_port);
   REG_reg_14_19_inst : DLH_X1 port map( G => n1935, D => n1702, Q => 
                           REG_14_19_port);
   REG_reg_14_18_inst : DLH_X1 port map( G => n1935, D => n1708, Q => 
                           REG_14_18_port);
   REG_reg_14_17_inst : DLH_X1 port map( G => n1935, D => n1714, Q => 
                           REG_14_17_port);
   REG_reg_14_16_inst : DLH_X1 port map( G => n1935, D => n1720, Q => 
                           REG_14_16_port);
   REG_reg_14_15_inst : DLH_X1 port map( G => n1935, D => n1726, Q => 
                           REG_14_15_port);
   REG_reg_14_14_inst : DLH_X1 port map( G => n1935, D => n1732, Q => 
                           REG_14_14_port);
   REG_reg_14_13_inst : DLH_X1 port map( G => n1935, D => n1738, Q => 
                           REG_14_13_port);
   REG_reg_14_12_inst : DLH_X1 port map( G => n1935, D => n1744, Q => 
                           REG_14_12_port);
   REG_reg_14_11_inst : DLH_X1 port map( G => n1935, D => n1750, Q => 
                           REG_14_11_port);
   REG_reg_14_10_inst : DLH_X1 port map( G => n1935, D => n1756, Q => 
                           REG_14_10_port);
   REG_reg_14_9_inst : DLH_X1 port map( G => n1934, D => n1762, Q => 
                           REG_14_9_port);
   REG_reg_14_8_inst : DLH_X1 port map( G => n1934, D => n1768, Q => 
                           REG_14_8_port);
   REG_reg_14_7_inst : DLH_X1 port map( G => n1934, D => n1774, Q => 
                           REG_14_7_port);
   REG_reg_14_6_inst : DLH_X1 port map( G => n1934, D => n1780, Q => 
                           REG_14_6_port);
   REG_reg_14_5_inst : DLH_X1 port map( G => n1934, D => n1786, Q => 
                           REG_14_5_port);
   REG_reg_14_4_inst : DLH_X1 port map( G => n1934, D => n1792, Q => 
                           REG_14_4_port);
   REG_reg_14_3_inst : DLH_X1 port map( G => n1934, D => n1798, Q => 
                           REG_14_3_port);
   REG_reg_14_2_inst : DLH_X1 port map( G => n1934, D => n1804, Q => 
                           REG_14_2_port);
   REG_reg_14_1_inst : DLH_X1 port map( G => n1934, D => n1810, Q => 
                           REG_14_1_port);
   REG_reg_14_0_inst : DLH_X1 port map( G => n1934, D => n1816, Q => 
                           REG_14_0_port);
   REG_reg_15_31_inst : DLH_X1 port map( G => n1944, D => n1630, Q => 
                           REG_15_31_port);
   REG_reg_15_30_inst : DLH_X1 port map( G => n1944, D => n1636, Q => 
                           REG_15_30_port);
   REG_reg_15_29_inst : DLH_X1 port map( G => n1943, D => n1642, Q => 
                           REG_15_29_port);
   REG_reg_15_28_inst : DLH_X1 port map( G => n1943, D => n1648, Q => 
                           REG_15_28_port);
   REG_reg_15_27_inst : DLH_X1 port map( G => n1943, D => n1654, Q => 
                           REG_15_27_port);
   REG_reg_15_26_inst : DLH_X1 port map( G => n1943, D => n1660, Q => 
                           REG_15_26_port);
   REG_reg_15_25_inst : DLH_X1 port map( G => n1943, D => n1666, Q => 
                           REG_15_25_port);
   REG_reg_15_24_inst : DLH_X1 port map( G => n1943, D => n1672, Q => 
                           REG_15_24_port);
   REG_reg_15_23_inst : DLH_X1 port map( G => n1943, D => n1678, Q => 
                           REG_15_23_port);
   REG_reg_15_22_inst : DLH_X1 port map( G => n1943, D => n1684, Q => 
                           REG_15_22_port);
   REG_reg_15_21_inst : DLH_X1 port map( G => n1943, D => n1690, Q => 
                           REG_15_21_port);
   REG_reg_15_20_inst : DLH_X1 port map( G => n1943, D => n1696, Q => 
                           REG_15_20_port);
   REG_reg_15_19_inst : DLH_X1 port map( G => n1942, D => n1702, Q => 
                           REG_15_19_port);
   REG_reg_15_18_inst : DLH_X1 port map( G => n1942, D => n1708, Q => 
                           REG_15_18_port);
   REG_reg_15_17_inst : DLH_X1 port map( G => n1942, D => n1714, Q => 
                           REG_15_17_port);
   REG_reg_15_16_inst : DLH_X1 port map( G => n1942, D => n1720, Q => 
                           REG_15_16_port);
   REG_reg_15_15_inst : DLH_X1 port map( G => n1942, D => n1726, Q => 
                           REG_15_15_port);
   REG_reg_15_14_inst : DLH_X1 port map( G => n1942, D => n1732, Q => 
                           REG_15_14_port);
   REG_reg_15_13_inst : DLH_X1 port map( G => n1942, D => n1738, Q => 
                           REG_15_13_port);
   REG_reg_15_12_inst : DLH_X1 port map( G => n1942, D => n1744, Q => 
                           REG_15_12_port);
   REG_reg_15_11_inst : DLH_X1 port map( G => n1942, D => n1750, Q => 
                           REG_15_11_port);
   REG_reg_15_10_inst : DLH_X1 port map( G => n1942, D => n1756, Q => 
                           REG_15_10_port);
   REG_reg_15_9_inst : DLH_X1 port map( G => n1941, D => n1762, Q => 
                           REG_15_9_port);
   REG_reg_15_8_inst : DLH_X1 port map( G => n1941, D => n1768, Q => 
                           REG_15_8_port);
   REG_reg_15_7_inst : DLH_X1 port map( G => n1941, D => n1774, Q => 
                           REG_15_7_port);
   REG_reg_15_6_inst : DLH_X1 port map( G => n1941, D => n1780, Q => 
                           REG_15_6_port);
   REG_reg_15_5_inst : DLH_X1 port map( G => n1941, D => n1786, Q => 
                           REG_15_5_port);
   REG_reg_15_4_inst : DLH_X1 port map( G => n1941, D => n1792, Q => 
                           REG_15_4_port);
   REG_reg_15_3_inst : DLH_X1 port map( G => n1941, D => n1798, Q => 
                           REG_15_3_port);
   REG_reg_15_2_inst : DLH_X1 port map( G => n1941, D => n1804, Q => 
                           REG_15_2_port);
   REG_reg_15_1_inst : DLH_X1 port map( G => n1941, D => n1810, Q => 
                           REG_15_1_port);
   REG_reg_15_0_inst : DLH_X1 port map( G => n1941, D => n1816, Q => 
                           REG_15_0_port);
   REG_reg_16_31_inst : DLH_X1 port map( G => n1951, D => n1630, Q => 
                           REG_16_31_port);
   REG_reg_16_30_inst : DLH_X1 port map( G => n1951, D => n1636, Q => 
                           REG_16_30_port);
   REG_reg_16_29_inst : DLH_X1 port map( G => n1950, D => n1642, Q => 
                           REG_16_29_port);
   REG_reg_16_28_inst : DLH_X1 port map( G => n1950, D => n1648, Q => 
                           REG_16_28_port);
   REG_reg_16_27_inst : DLH_X1 port map( G => n1950, D => n1654, Q => 
                           REG_16_27_port);
   REG_reg_16_26_inst : DLH_X1 port map( G => n1950, D => n1660, Q => 
                           REG_16_26_port);
   REG_reg_16_25_inst : DLH_X1 port map( G => n1950, D => n1666, Q => 
                           REG_16_25_port);
   REG_reg_16_24_inst : DLH_X1 port map( G => n1950, D => n1672, Q => 
                           REG_16_24_port);
   REG_reg_16_23_inst : DLH_X1 port map( G => n1950, D => n1678, Q => 
                           REG_16_23_port);
   REG_reg_16_22_inst : DLH_X1 port map( G => n1950, D => n1684, Q => 
                           REG_16_22_port);
   REG_reg_16_21_inst : DLH_X1 port map( G => n1950, D => n1690, Q => 
                           REG_16_21_port);
   REG_reg_16_20_inst : DLH_X1 port map( G => n1950, D => n1696, Q => 
                           REG_16_20_port);
   REG_reg_16_19_inst : DLH_X1 port map( G => n1949, D => n1702, Q => 
                           REG_16_19_port);
   REG_reg_16_18_inst : DLH_X1 port map( G => n1949, D => n1708, Q => 
                           REG_16_18_port);
   REG_reg_16_17_inst : DLH_X1 port map( G => n1949, D => n1714, Q => 
                           REG_16_17_port);
   REG_reg_16_16_inst : DLH_X1 port map( G => n1949, D => n1720, Q => 
                           REG_16_16_port);
   REG_reg_16_15_inst : DLH_X1 port map( G => n1949, D => n1726, Q => 
                           REG_16_15_port);
   REG_reg_16_14_inst : DLH_X1 port map( G => n1949, D => n1732, Q => 
                           REG_16_14_port);
   REG_reg_16_13_inst : DLH_X1 port map( G => n1949, D => n1738, Q => 
                           REG_16_13_port);
   REG_reg_16_12_inst : DLH_X1 port map( G => n1949, D => n1744, Q => 
                           REG_16_12_port);
   REG_reg_16_11_inst : DLH_X1 port map( G => n1949, D => n1750, Q => 
                           REG_16_11_port);
   REG_reg_16_10_inst : DLH_X1 port map( G => n1949, D => n1756, Q => 
                           REG_16_10_port);
   REG_reg_16_9_inst : DLH_X1 port map( G => n1948, D => n1762, Q => 
                           REG_16_9_port);
   REG_reg_16_8_inst : DLH_X1 port map( G => n1948, D => n1768, Q => 
                           REG_16_8_port);
   REG_reg_16_7_inst : DLH_X1 port map( G => n1948, D => n1774, Q => 
                           REG_16_7_port);
   REG_reg_16_6_inst : DLH_X1 port map( G => n1948, D => n1780, Q => 
                           REG_16_6_port);
   REG_reg_16_5_inst : DLH_X1 port map( G => n1948, D => n1786, Q => 
                           REG_16_5_port);
   REG_reg_16_4_inst : DLH_X1 port map( G => n1948, D => n1792, Q => 
                           REG_16_4_port);
   REG_reg_16_3_inst : DLH_X1 port map( G => n1948, D => n1798, Q => 
                           REG_16_3_port);
   REG_reg_16_2_inst : DLH_X1 port map( G => n1948, D => n1804, Q => 
                           REG_16_2_port);
   REG_reg_16_1_inst : DLH_X1 port map( G => n1948, D => n1810, Q => 
                           REG_16_1_port);
   REG_reg_16_0_inst : DLH_X1 port map( G => n1948, D => n1816, Q => 
                           REG_16_0_port);
   REG_reg_17_31_inst : DLH_X1 port map( G => n1958, D => n1630, Q => 
                           REG_17_31_port);
   REG_reg_17_30_inst : DLH_X1 port map( G => n1958, D => n1636, Q => 
                           REG_17_30_port);
   REG_reg_17_29_inst : DLH_X1 port map( G => n1957, D => n1642, Q => 
                           REG_17_29_port);
   REG_reg_17_28_inst : DLH_X1 port map( G => n1957, D => n1648, Q => 
                           REG_17_28_port);
   REG_reg_17_27_inst : DLH_X1 port map( G => n1957, D => n1654, Q => 
                           REG_17_27_port);
   REG_reg_17_26_inst : DLH_X1 port map( G => n1957, D => n1660, Q => 
                           REG_17_26_port);
   REG_reg_17_25_inst : DLH_X1 port map( G => n1957, D => n1666, Q => 
                           REG_17_25_port);
   REG_reg_17_24_inst : DLH_X1 port map( G => n1957, D => n1672, Q => 
                           REG_17_24_port);
   REG_reg_17_23_inst : DLH_X1 port map( G => n1957, D => n1678, Q => 
                           REG_17_23_port);
   REG_reg_17_22_inst : DLH_X1 port map( G => n1957, D => n1684, Q => 
                           REG_17_22_port);
   REG_reg_17_21_inst : DLH_X1 port map( G => n1957, D => n1690, Q => 
                           REG_17_21_port);
   REG_reg_17_20_inst : DLH_X1 port map( G => n1957, D => n1696, Q => 
                           REG_17_20_port);
   REG_reg_17_19_inst : DLH_X1 port map( G => n1956, D => n1702, Q => 
                           REG_17_19_port);
   REG_reg_17_18_inst : DLH_X1 port map( G => n1956, D => n1708, Q => 
                           REG_17_18_port);
   REG_reg_17_17_inst : DLH_X1 port map( G => n1956, D => n1714, Q => 
                           REG_17_17_port);
   REG_reg_17_16_inst : DLH_X1 port map( G => n1956, D => n1720, Q => 
                           REG_17_16_port);
   REG_reg_17_15_inst : DLH_X1 port map( G => n1956, D => n1726, Q => 
                           REG_17_15_port);
   REG_reg_17_14_inst : DLH_X1 port map( G => n1956, D => n1732, Q => 
                           REG_17_14_port);
   REG_reg_17_13_inst : DLH_X1 port map( G => n1956, D => n1738, Q => 
                           REG_17_13_port);
   REG_reg_17_12_inst : DLH_X1 port map( G => n1956, D => n1744, Q => 
                           REG_17_12_port);
   REG_reg_17_11_inst : DLH_X1 port map( G => n1956, D => n1750, Q => 
                           REG_17_11_port);
   REG_reg_17_10_inst : DLH_X1 port map( G => n1956, D => n1756, Q => 
                           REG_17_10_port);
   REG_reg_17_9_inst : DLH_X1 port map( G => n1955, D => n1762, Q => 
                           REG_17_9_port);
   REG_reg_17_8_inst : DLH_X1 port map( G => n1955, D => n1768, Q => 
                           REG_17_8_port);
   REG_reg_17_7_inst : DLH_X1 port map( G => n1955, D => n1774, Q => 
                           REG_17_7_port);
   REG_reg_17_6_inst : DLH_X1 port map( G => n1955, D => n1780, Q => 
                           REG_17_6_port);
   REG_reg_17_5_inst : DLH_X1 port map( G => n1955, D => n1786, Q => 
                           REG_17_5_port);
   REG_reg_17_4_inst : DLH_X1 port map( G => n1955, D => n1792, Q => 
                           REG_17_4_port);
   REG_reg_17_3_inst : DLH_X1 port map( G => n1955, D => n1798, Q => 
                           REG_17_3_port);
   REG_reg_17_2_inst : DLH_X1 port map( G => n1955, D => n1804, Q => 
                           REG_17_2_port);
   REG_reg_17_1_inst : DLH_X1 port map( G => n1955, D => n1810, Q => 
                           REG_17_1_port);
   REG_reg_17_0_inst : DLH_X1 port map( G => n1955, D => n1816, Q => 
                           REG_17_0_port);
   REG_reg_18_31_inst : DLH_X1 port map( G => n1965, D => n1630, Q => 
                           REG_18_31_port);
   REG_reg_18_30_inst : DLH_X1 port map( G => n1965, D => n1636, Q => 
                           REG_18_30_port);
   REG_reg_18_29_inst : DLH_X1 port map( G => n1964, D => n1642, Q => 
                           REG_18_29_port);
   REG_reg_18_28_inst : DLH_X1 port map( G => n1964, D => n1648, Q => 
                           REG_18_28_port);
   REG_reg_18_27_inst : DLH_X1 port map( G => n1964, D => n1654, Q => 
                           REG_18_27_port);
   REG_reg_18_26_inst : DLH_X1 port map( G => n1964, D => n1660, Q => 
                           REG_18_26_port);
   REG_reg_18_25_inst : DLH_X1 port map( G => n1964, D => n1666, Q => 
                           REG_18_25_port);
   REG_reg_18_24_inst : DLH_X1 port map( G => n1964, D => n1672, Q => 
                           REG_18_24_port);
   REG_reg_18_23_inst : DLH_X1 port map( G => n1964, D => n1678, Q => 
                           REG_18_23_port);
   REG_reg_18_22_inst : DLH_X1 port map( G => n1964, D => n1684, Q => 
                           REG_18_22_port);
   REG_reg_18_21_inst : DLH_X1 port map( G => n1964, D => n1690, Q => 
                           REG_18_21_port);
   REG_reg_18_20_inst : DLH_X1 port map( G => n1964, D => n1696, Q => 
                           REG_18_20_port);
   REG_reg_18_19_inst : DLH_X1 port map( G => n1963, D => n1702, Q => 
                           REG_18_19_port);
   REG_reg_18_18_inst : DLH_X1 port map( G => n1963, D => n1708, Q => 
                           REG_18_18_port);
   REG_reg_18_17_inst : DLH_X1 port map( G => n1963, D => n1714, Q => 
                           REG_18_17_port);
   REG_reg_18_16_inst : DLH_X1 port map( G => n1963, D => n1720, Q => 
                           REG_18_16_port);
   REG_reg_18_15_inst : DLH_X1 port map( G => n1963, D => n1726, Q => 
                           REG_18_15_port);
   REG_reg_18_14_inst : DLH_X1 port map( G => n1963, D => n1732, Q => 
                           REG_18_14_port);
   REG_reg_18_13_inst : DLH_X1 port map( G => n1963, D => n1738, Q => 
                           REG_18_13_port);
   REG_reg_18_12_inst : DLH_X1 port map( G => n1963, D => n1744, Q => 
                           REG_18_12_port);
   REG_reg_18_11_inst : DLH_X1 port map( G => n1963, D => n1750, Q => 
                           REG_18_11_port);
   REG_reg_18_10_inst : DLH_X1 port map( G => n1963, D => n1756, Q => 
                           REG_18_10_port);
   REG_reg_18_9_inst : DLH_X1 port map( G => n1962, D => n1762, Q => 
                           REG_18_9_port);
   REG_reg_18_8_inst : DLH_X1 port map( G => n1962, D => n1768, Q => 
                           REG_18_8_port);
   REG_reg_18_7_inst : DLH_X1 port map( G => n1962, D => n1774, Q => 
                           REG_18_7_port);
   REG_reg_18_6_inst : DLH_X1 port map( G => n1962, D => n1780, Q => 
                           REG_18_6_port);
   REG_reg_18_5_inst : DLH_X1 port map( G => n1962, D => n1786, Q => 
                           REG_18_5_port);
   REG_reg_18_4_inst : DLH_X1 port map( G => n1962, D => n1792, Q => 
                           REG_18_4_port);
   REG_reg_18_3_inst : DLH_X1 port map( G => n1962, D => n1798, Q => 
                           REG_18_3_port);
   REG_reg_18_2_inst : DLH_X1 port map( G => n1962, D => n1804, Q => 
                           REG_18_2_port);
   REG_reg_18_1_inst : DLH_X1 port map( G => n1962, D => n1810, Q => 
                           REG_18_1_port);
   REG_reg_18_0_inst : DLH_X1 port map( G => n1962, D => n1816, Q => 
                           REG_18_0_port);
   REG_reg_19_31_inst : DLH_X1 port map( G => n1972, D => n1630, Q => 
                           REG_19_31_port);
   REG_reg_19_30_inst : DLH_X1 port map( G => n1972, D => n1636, Q => 
                           REG_19_30_port);
   REG_reg_19_29_inst : DLH_X1 port map( G => n1971, D => n1642, Q => 
                           REG_19_29_port);
   REG_reg_19_28_inst : DLH_X1 port map( G => n1971, D => n1648, Q => 
                           REG_19_28_port);
   REG_reg_19_27_inst : DLH_X1 port map( G => n1971, D => n1654, Q => 
                           REG_19_27_port);
   REG_reg_19_26_inst : DLH_X1 port map( G => n1971, D => n1660, Q => 
                           REG_19_26_port);
   REG_reg_19_25_inst : DLH_X1 port map( G => n1971, D => n1666, Q => 
                           REG_19_25_port);
   REG_reg_19_24_inst : DLH_X1 port map( G => n1971, D => n1672, Q => 
                           REG_19_24_port);
   REG_reg_19_23_inst : DLH_X1 port map( G => n1971, D => n1678, Q => 
                           REG_19_23_port);
   REG_reg_19_22_inst : DLH_X1 port map( G => n1971, D => n1684, Q => 
                           REG_19_22_port);
   REG_reg_19_21_inst : DLH_X1 port map( G => n1971, D => n1690, Q => 
                           REG_19_21_port);
   REG_reg_19_20_inst : DLH_X1 port map( G => n1971, D => n1696, Q => 
                           REG_19_20_port);
   REG_reg_19_19_inst : DLH_X1 port map( G => n1970, D => n1702, Q => 
                           REG_19_19_port);
   REG_reg_19_18_inst : DLH_X1 port map( G => n1970, D => n1708, Q => 
                           REG_19_18_port);
   REG_reg_19_17_inst : DLH_X1 port map( G => n1970, D => n1714, Q => 
                           REG_19_17_port);
   REG_reg_19_16_inst : DLH_X1 port map( G => n1970, D => n1720, Q => 
                           REG_19_16_port);
   REG_reg_19_15_inst : DLH_X1 port map( G => n1970, D => n1726, Q => 
                           REG_19_15_port);
   REG_reg_19_14_inst : DLH_X1 port map( G => n1970, D => n1732, Q => 
                           REG_19_14_port);
   REG_reg_19_13_inst : DLH_X1 port map( G => n1970, D => n1738, Q => 
                           REG_19_13_port);
   REG_reg_19_12_inst : DLH_X1 port map( G => n1970, D => n1744, Q => 
                           REG_19_12_port);
   REG_reg_19_11_inst : DLH_X1 port map( G => n1970, D => n1750, Q => 
                           REG_19_11_port);
   REG_reg_19_10_inst : DLH_X1 port map( G => n1970, D => n1756, Q => 
                           REG_19_10_port);
   REG_reg_19_9_inst : DLH_X1 port map( G => n1969, D => n1762, Q => 
                           REG_19_9_port);
   REG_reg_19_8_inst : DLH_X1 port map( G => n1969, D => n1768, Q => 
                           REG_19_8_port);
   REG_reg_19_7_inst : DLH_X1 port map( G => n1969, D => n1774, Q => 
                           REG_19_7_port);
   REG_reg_19_6_inst : DLH_X1 port map( G => n1969, D => n1780, Q => 
                           REG_19_6_port);
   REG_reg_19_5_inst : DLH_X1 port map( G => n1969, D => n1786, Q => 
                           REG_19_5_port);
   REG_reg_19_4_inst : DLH_X1 port map( G => n1969, D => n1792, Q => 
                           REG_19_4_port);
   REG_reg_19_3_inst : DLH_X1 port map( G => n1969, D => n1798, Q => 
                           REG_19_3_port);
   REG_reg_19_2_inst : DLH_X1 port map( G => n1969, D => n1804, Q => 
                           REG_19_2_port);
   REG_reg_19_1_inst : DLH_X1 port map( G => n1969, D => n1810, Q => 
                           REG_19_1_port);
   REG_reg_19_0_inst : DLH_X1 port map( G => n1969, D => n1816, Q => 
                           REG_19_0_port);
   REG_reg_20_31_inst : DLH_X1 port map( G => n1979, D => n1630, Q => 
                           REG_20_31_port);
   REG_reg_20_30_inst : DLH_X1 port map( G => n1979, D => n1636, Q => 
                           REG_20_30_port);
   REG_reg_20_29_inst : DLH_X1 port map( G => n1978, D => n1642, Q => 
                           REG_20_29_port);
   REG_reg_20_28_inst : DLH_X1 port map( G => n1978, D => n1648, Q => 
                           REG_20_28_port);
   REG_reg_20_27_inst : DLH_X1 port map( G => n1978, D => n1654, Q => 
                           REG_20_27_port);
   REG_reg_20_26_inst : DLH_X1 port map( G => n1978, D => n1660, Q => 
                           REG_20_26_port);
   REG_reg_20_25_inst : DLH_X1 port map( G => n1978, D => n1666, Q => 
                           REG_20_25_port);
   REG_reg_20_24_inst : DLH_X1 port map( G => n1978, D => n1672, Q => 
                           REG_20_24_port);
   REG_reg_20_23_inst : DLH_X1 port map( G => n1978, D => n1678, Q => 
                           REG_20_23_port);
   REG_reg_20_22_inst : DLH_X1 port map( G => n1978, D => n1684, Q => 
                           REG_20_22_port);
   REG_reg_20_21_inst : DLH_X1 port map( G => n1978, D => n1690, Q => 
                           REG_20_21_port);
   REG_reg_20_20_inst : DLH_X1 port map( G => n1978, D => n1696, Q => 
                           REG_20_20_port);
   REG_reg_20_19_inst : DLH_X1 port map( G => n1977, D => n1702, Q => 
                           REG_20_19_port);
   REG_reg_20_18_inst : DLH_X1 port map( G => n1977, D => n1708, Q => 
                           REG_20_18_port);
   REG_reg_20_17_inst : DLH_X1 port map( G => n1977, D => n1714, Q => 
                           REG_20_17_port);
   REG_reg_20_16_inst : DLH_X1 port map( G => n1977, D => n1720, Q => 
                           REG_20_16_port);
   REG_reg_20_15_inst : DLH_X1 port map( G => n1977, D => n1726, Q => 
                           REG_20_15_port);
   REG_reg_20_14_inst : DLH_X1 port map( G => n1977, D => n1732, Q => 
                           REG_20_14_port);
   REG_reg_20_13_inst : DLH_X1 port map( G => n1977, D => n1738, Q => 
                           REG_20_13_port);
   REG_reg_20_12_inst : DLH_X1 port map( G => n1977, D => n1744, Q => 
                           REG_20_12_port);
   REG_reg_20_11_inst : DLH_X1 port map( G => n1977, D => n1750, Q => 
                           REG_20_11_port);
   REG_reg_20_10_inst : DLH_X1 port map( G => n1977, D => n1756, Q => 
                           REG_20_10_port);
   REG_reg_20_9_inst : DLH_X1 port map( G => n1976, D => n1762, Q => 
                           REG_20_9_port);
   REG_reg_20_8_inst : DLH_X1 port map( G => n1976, D => n1768, Q => 
                           REG_20_8_port);
   REG_reg_20_7_inst : DLH_X1 port map( G => n1976, D => n1774, Q => 
                           REG_20_7_port);
   REG_reg_20_6_inst : DLH_X1 port map( G => n1976, D => n1780, Q => 
                           REG_20_6_port);
   REG_reg_20_5_inst : DLH_X1 port map( G => n1976, D => n1786, Q => 
                           REG_20_5_port);
   REG_reg_20_4_inst : DLH_X1 port map( G => n1976, D => n1792, Q => 
                           REG_20_4_port);
   REG_reg_20_3_inst : DLH_X1 port map( G => n1976, D => n1798, Q => 
                           REG_20_3_port);
   REG_reg_20_2_inst : DLH_X1 port map( G => n1976, D => n1804, Q => 
                           REG_20_2_port);
   REG_reg_20_1_inst : DLH_X1 port map( G => n1976, D => n1810, Q => 
                           REG_20_1_port);
   REG_reg_20_0_inst : DLH_X1 port map( G => n1976, D => n1816, Q => 
                           REG_20_0_port);
   REG_reg_21_31_inst : DLH_X1 port map( G => n1986, D => n1631, Q => 
                           REG_21_31_port);
   REG_reg_21_30_inst : DLH_X1 port map( G => n1986, D => n1637, Q => 
                           REG_21_30_port);
   REG_reg_21_29_inst : DLH_X1 port map( G => n1985, D => n1643, Q => 
                           REG_21_29_port);
   REG_reg_21_28_inst : DLH_X1 port map( G => n1985, D => n1649, Q => 
                           REG_21_28_port);
   REG_reg_21_27_inst : DLH_X1 port map( G => n1985, D => n1655, Q => 
                           REG_21_27_port);
   REG_reg_21_26_inst : DLH_X1 port map( G => n1985, D => n1661, Q => 
                           REG_21_26_port);
   REG_reg_21_25_inst : DLH_X1 port map( G => n1985, D => n1667, Q => 
                           REG_21_25_port);
   REG_reg_21_24_inst : DLH_X1 port map( G => n1985, D => n1673, Q => 
                           REG_21_24_port);
   REG_reg_21_23_inst : DLH_X1 port map( G => n1985, D => n1679, Q => 
                           REG_21_23_port);
   REG_reg_21_22_inst : DLH_X1 port map( G => n1985, D => n1685, Q => 
                           REG_21_22_port);
   REG_reg_21_21_inst : DLH_X1 port map( G => n1985, D => n1691, Q => 
                           REG_21_21_port);
   REG_reg_21_20_inst : DLH_X1 port map( G => n1985, D => n1697, Q => 
                           REG_21_20_port);
   REG_reg_21_19_inst : DLH_X1 port map( G => n1984, D => n1703, Q => 
                           REG_21_19_port);
   REG_reg_21_18_inst : DLH_X1 port map( G => n1984, D => n1709, Q => 
                           REG_21_18_port);
   REG_reg_21_17_inst : DLH_X1 port map( G => n1984, D => n1715, Q => 
                           REG_21_17_port);
   REG_reg_21_16_inst : DLH_X1 port map( G => n1984, D => n1721, Q => 
                           REG_21_16_port);
   REG_reg_21_15_inst : DLH_X1 port map( G => n1984, D => n1727, Q => 
                           REG_21_15_port);
   REG_reg_21_14_inst : DLH_X1 port map( G => n1984, D => n1733, Q => 
                           REG_21_14_port);
   REG_reg_21_13_inst : DLH_X1 port map( G => n1984, D => n1739, Q => 
                           REG_21_13_port);
   REG_reg_21_12_inst : DLH_X1 port map( G => n1984, D => n1745, Q => 
                           REG_21_12_port);
   REG_reg_21_11_inst : DLH_X1 port map( G => n1984, D => n1751, Q => 
                           REG_21_11_port);
   REG_reg_21_10_inst : DLH_X1 port map( G => n1984, D => n1757, Q => 
                           REG_21_10_port);
   REG_reg_21_9_inst : DLH_X1 port map( G => n1983, D => n1763, Q => 
                           REG_21_9_port);
   REG_reg_21_8_inst : DLH_X1 port map( G => n1983, D => n1769, Q => 
                           REG_21_8_port);
   REG_reg_21_7_inst : DLH_X1 port map( G => n1983, D => n1775, Q => 
                           REG_21_7_port);
   REG_reg_21_6_inst : DLH_X1 port map( G => n1983, D => n1781, Q => 
                           REG_21_6_port);
   REG_reg_21_5_inst : DLH_X1 port map( G => n1983, D => n1787, Q => 
                           REG_21_5_port);
   REG_reg_21_4_inst : DLH_X1 port map( G => n1983, D => n1793, Q => 
                           REG_21_4_port);
   REG_reg_21_3_inst : DLH_X1 port map( G => n1983, D => n1799, Q => 
                           REG_21_3_port);
   REG_reg_21_2_inst : DLH_X1 port map( G => n1983, D => n1805, Q => 
                           REG_21_2_port);
   REG_reg_21_1_inst : DLH_X1 port map( G => n1983, D => n1811, Q => 
                           REG_21_1_port);
   REG_reg_21_0_inst : DLH_X1 port map( G => n1983, D => n1817, Q => 
                           REG_21_0_port);
   REG_reg_22_31_inst : DLH_X1 port map( G => n1993, D => n1631, Q => 
                           REG_22_31_port);
   REG_reg_22_30_inst : DLH_X1 port map( G => n1993, D => n1637, Q => 
                           REG_22_30_port);
   REG_reg_22_29_inst : DLH_X1 port map( G => n1992, D => n1643, Q => 
                           REG_22_29_port);
   REG_reg_22_28_inst : DLH_X1 port map( G => n1992, D => n1649, Q => 
                           REG_22_28_port);
   REG_reg_22_27_inst : DLH_X1 port map( G => n1992, D => n1655, Q => 
                           REG_22_27_port);
   REG_reg_22_26_inst : DLH_X1 port map( G => n1992, D => n1661, Q => 
                           REG_22_26_port);
   REG_reg_22_25_inst : DLH_X1 port map( G => n1992, D => n1667, Q => 
                           REG_22_25_port);
   REG_reg_22_24_inst : DLH_X1 port map( G => n1992, D => n1673, Q => 
                           REG_22_24_port);
   REG_reg_22_23_inst : DLH_X1 port map( G => n1992, D => n1679, Q => 
                           REG_22_23_port);
   REG_reg_22_22_inst : DLH_X1 port map( G => n1992, D => n1685, Q => 
                           REG_22_22_port);
   REG_reg_22_21_inst : DLH_X1 port map( G => n1992, D => n1691, Q => 
                           REG_22_21_port);
   REG_reg_22_20_inst : DLH_X1 port map( G => n1992, D => n1697, Q => 
                           REG_22_20_port);
   REG_reg_22_19_inst : DLH_X1 port map( G => n1991, D => n1703, Q => 
                           REG_22_19_port);
   REG_reg_22_18_inst : DLH_X1 port map( G => n1991, D => n1709, Q => 
                           REG_22_18_port);
   REG_reg_22_17_inst : DLH_X1 port map( G => n1991, D => n1715, Q => 
                           REG_22_17_port);
   REG_reg_22_16_inst : DLH_X1 port map( G => n1991, D => n1721, Q => 
                           REG_22_16_port);
   REG_reg_22_15_inst : DLH_X1 port map( G => n1991, D => n1727, Q => 
                           REG_22_15_port);
   REG_reg_22_14_inst : DLH_X1 port map( G => n1991, D => n1733, Q => 
                           REG_22_14_port);
   REG_reg_22_13_inst : DLH_X1 port map( G => n1991, D => n1739, Q => 
                           REG_22_13_port);
   REG_reg_22_12_inst : DLH_X1 port map( G => n1991, D => n1745, Q => 
                           REG_22_12_port);
   REG_reg_22_11_inst : DLH_X1 port map( G => n1991, D => n1751, Q => 
                           REG_22_11_port);
   REG_reg_22_10_inst : DLH_X1 port map( G => n1991, D => n1757, Q => 
                           REG_22_10_port);
   REG_reg_22_9_inst : DLH_X1 port map( G => n1990, D => n1763, Q => 
                           REG_22_9_port);
   REG_reg_22_8_inst : DLH_X1 port map( G => n1990, D => n1769, Q => 
                           REG_22_8_port);
   REG_reg_22_7_inst : DLH_X1 port map( G => n1990, D => n1775, Q => 
                           REG_22_7_port);
   REG_reg_22_6_inst : DLH_X1 port map( G => n1990, D => n1781, Q => 
                           REG_22_6_port);
   REG_reg_22_5_inst : DLH_X1 port map( G => n1990, D => n1787, Q => 
                           REG_22_5_port);
   REG_reg_22_4_inst : DLH_X1 port map( G => n1990, D => n1793, Q => 
                           REG_22_4_port);
   REG_reg_22_3_inst : DLH_X1 port map( G => n1990, D => n1799, Q => 
                           REG_22_3_port);
   REG_reg_22_2_inst : DLH_X1 port map( G => n1990, D => n1805, Q => 
                           REG_22_2_port);
   REG_reg_22_1_inst : DLH_X1 port map( G => n1990, D => n1811, Q => 
                           REG_22_1_port);
   REG_reg_22_0_inst : DLH_X1 port map( G => n1990, D => n1817, Q => 
                           REG_22_0_port);
   REG_reg_23_31_inst : DLH_X1 port map( G => n2000, D => n1631, Q => 
                           REG_23_31_port);
   REG_reg_23_30_inst : DLH_X1 port map( G => n2000, D => n1637, Q => 
                           REG_23_30_port);
   REG_reg_23_29_inst : DLH_X1 port map( G => n1999, D => n1643, Q => 
                           REG_23_29_port);
   REG_reg_23_28_inst : DLH_X1 port map( G => n1999, D => n1649, Q => 
                           REG_23_28_port);
   REG_reg_23_27_inst : DLH_X1 port map( G => n1999, D => n1655, Q => 
                           REG_23_27_port);
   REG_reg_23_26_inst : DLH_X1 port map( G => n1999, D => n1661, Q => 
                           REG_23_26_port);
   REG_reg_23_25_inst : DLH_X1 port map( G => n1999, D => n1667, Q => 
                           REG_23_25_port);
   REG_reg_23_24_inst : DLH_X1 port map( G => n1999, D => n1673, Q => 
                           REG_23_24_port);
   REG_reg_23_23_inst : DLH_X1 port map( G => n1999, D => n1679, Q => 
                           REG_23_23_port);
   REG_reg_23_22_inst : DLH_X1 port map( G => n1999, D => n1685, Q => 
                           REG_23_22_port);
   REG_reg_23_21_inst : DLH_X1 port map( G => n1999, D => n1691, Q => 
                           REG_23_21_port);
   REG_reg_23_20_inst : DLH_X1 port map( G => n1999, D => n1697, Q => 
                           REG_23_20_port);
   REG_reg_23_19_inst : DLH_X1 port map( G => n1998, D => n1703, Q => 
                           REG_23_19_port);
   REG_reg_23_18_inst : DLH_X1 port map( G => n1998, D => n1709, Q => 
                           REG_23_18_port);
   REG_reg_23_17_inst : DLH_X1 port map( G => n1998, D => n1715, Q => 
                           REG_23_17_port);
   REG_reg_23_16_inst : DLH_X1 port map( G => n1998, D => n1721, Q => 
                           REG_23_16_port);
   REG_reg_23_15_inst : DLH_X1 port map( G => n1998, D => n1727, Q => 
                           REG_23_15_port);
   REG_reg_23_14_inst : DLH_X1 port map( G => n1998, D => n1733, Q => 
                           REG_23_14_port);
   REG_reg_23_13_inst : DLH_X1 port map( G => n1998, D => n1739, Q => 
                           REG_23_13_port);
   REG_reg_23_12_inst : DLH_X1 port map( G => n1998, D => n1745, Q => 
                           REG_23_12_port);
   REG_reg_23_11_inst : DLH_X1 port map( G => n1998, D => n1751, Q => 
                           REG_23_11_port);
   REG_reg_23_10_inst : DLH_X1 port map( G => n1998, D => n1757, Q => 
                           REG_23_10_port);
   REG_reg_23_9_inst : DLH_X1 port map( G => n1997, D => n1763, Q => 
                           REG_23_9_port);
   REG_reg_23_8_inst : DLH_X1 port map( G => n1997, D => n1769, Q => 
                           REG_23_8_port);
   REG_reg_23_7_inst : DLH_X1 port map( G => n1997, D => n1775, Q => 
                           REG_23_7_port);
   REG_reg_23_6_inst : DLH_X1 port map( G => n1997, D => n1781, Q => 
                           REG_23_6_port);
   REG_reg_23_5_inst : DLH_X1 port map( G => n1997, D => n1787, Q => 
                           REG_23_5_port);
   REG_reg_23_4_inst : DLH_X1 port map( G => n1997, D => n1793, Q => 
                           REG_23_4_port);
   REG_reg_23_3_inst : DLH_X1 port map( G => n1997, D => n1799, Q => 
                           REG_23_3_port);
   REG_reg_23_2_inst : DLH_X1 port map( G => n1997, D => n1805, Q => 
                           REG_23_2_port);
   REG_reg_23_1_inst : DLH_X1 port map( G => n1997, D => n1811, Q => 
                           REG_23_1_port);
   REG_reg_23_0_inst : DLH_X1 port map( G => n1997, D => n1817, Q => 
                           REG_23_0_port);
   REG_reg_24_31_inst : DLH_X1 port map( G => n2007, D => n1631, Q => 
                           REG_24_31_port);
   REG_reg_24_30_inst : DLH_X1 port map( G => n2007, D => n1637, Q => 
                           REG_24_30_port);
   REG_reg_24_29_inst : DLH_X1 port map( G => n2006, D => n1643, Q => 
                           REG_24_29_port);
   REG_reg_24_28_inst : DLH_X1 port map( G => n2006, D => n1649, Q => 
                           REG_24_28_port);
   REG_reg_24_27_inst : DLH_X1 port map( G => n2006, D => n1655, Q => 
                           REG_24_27_port);
   REG_reg_24_26_inst : DLH_X1 port map( G => n2006, D => n1661, Q => 
                           REG_24_26_port);
   REG_reg_24_25_inst : DLH_X1 port map( G => n2006, D => n1667, Q => 
                           REG_24_25_port);
   REG_reg_24_24_inst : DLH_X1 port map( G => n2006, D => n1673, Q => 
                           REG_24_24_port);
   REG_reg_24_23_inst : DLH_X1 port map( G => n2006, D => n1679, Q => 
                           REG_24_23_port);
   REG_reg_24_22_inst : DLH_X1 port map( G => n2006, D => n1685, Q => 
                           REG_24_22_port);
   REG_reg_24_21_inst : DLH_X1 port map( G => n2006, D => n1691, Q => 
                           REG_24_21_port);
   REG_reg_24_20_inst : DLH_X1 port map( G => n2006, D => n1697, Q => 
                           REG_24_20_port);
   REG_reg_24_19_inst : DLH_X1 port map( G => n2005, D => n1703, Q => 
                           REG_24_19_port);
   REG_reg_24_18_inst : DLH_X1 port map( G => n2005, D => n1709, Q => 
                           REG_24_18_port);
   REG_reg_24_17_inst : DLH_X1 port map( G => n2005, D => n1715, Q => 
                           REG_24_17_port);
   REG_reg_24_16_inst : DLH_X1 port map( G => n2005, D => n1721, Q => 
                           REG_24_16_port);
   REG_reg_24_15_inst : DLH_X1 port map( G => n2005, D => n1727, Q => 
                           REG_24_15_port);
   REG_reg_24_14_inst : DLH_X1 port map( G => n2005, D => n1733, Q => 
                           REG_24_14_port);
   REG_reg_24_13_inst : DLH_X1 port map( G => n2005, D => n1739, Q => 
                           REG_24_13_port);
   REG_reg_24_12_inst : DLH_X1 port map( G => n2005, D => n1745, Q => 
                           REG_24_12_port);
   REG_reg_24_11_inst : DLH_X1 port map( G => n2005, D => n1751, Q => 
                           REG_24_11_port);
   REG_reg_24_10_inst : DLH_X1 port map( G => n2005, D => n1757, Q => 
                           REG_24_10_port);
   REG_reg_24_9_inst : DLH_X1 port map( G => n2004, D => n1763, Q => 
                           REG_24_9_port);
   REG_reg_24_8_inst : DLH_X1 port map( G => n2004, D => n1769, Q => 
                           REG_24_8_port);
   REG_reg_24_7_inst : DLH_X1 port map( G => n2004, D => n1775, Q => 
                           REG_24_7_port);
   REG_reg_24_6_inst : DLH_X1 port map( G => n2004, D => n1781, Q => 
                           REG_24_6_port);
   REG_reg_24_5_inst : DLH_X1 port map( G => n2004, D => n1787, Q => 
                           REG_24_5_port);
   REG_reg_24_4_inst : DLH_X1 port map( G => n2004, D => n1793, Q => 
                           REG_24_4_port);
   REG_reg_24_3_inst : DLH_X1 port map( G => n2004, D => n1799, Q => 
                           REG_24_3_port);
   REG_reg_24_2_inst : DLH_X1 port map( G => n2004, D => n1805, Q => 
                           REG_24_2_port);
   REG_reg_24_1_inst : DLH_X1 port map( G => n2004, D => n1811, Q => 
                           REG_24_1_port);
   REG_reg_24_0_inst : DLH_X1 port map( G => n2004, D => n1817, Q => 
                           REG_24_0_port);
   REG_reg_25_31_inst : DLH_X1 port map( G => n2014, D => n1631, Q => 
                           REG_25_31_port);
   REG_reg_25_30_inst : DLH_X1 port map( G => n2014, D => n1637, Q => 
                           REG_25_30_port);
   REG_reg_25_29_inst : DLH_X1 port map( G => n2013, D => n1643, Q => 
                           REG_25_29_port);
   REG_reg_25_28_inst : DLH_X1 port map( G => n2013, D => n1649, Q => 
                           REG_25_28_port);
   REG_reg_25_27_inst : DLH_X1 port map( G => n2013, D => n1655, Q => 
                           REG_25_27_port);
   REG_reg_25_26_inst : DLH_X1 port map( G => n2013, D => n1661, Q => 
                           REG_25_26_port);
   REG_reg_25_25_inst : DLH_X1 port map( G => n2013, D => n1667, Q => 
                           REG_25_25_port);
   REG_reg_25_24_inst : DLH_X1 port map( G => n2013, D => n1673, Q => 
                           REG_25_24_port);
   REG_reg_25_23_inst : DLH_X1 port map( G => n2013, D => n1679, Q => 
                           REG_25_23_port);
   REG_reg_25_22_inst : DLH_X1 port map( G => n2013, D => n1685, Q => 
                           REG_25_22_port);
   REG_reg_25_21_inst : DLH_X1 port map( G => n2013, D => n1691, Q => 
                           REG_25_21_port);
   REG_reg_25_20_inst : DLH_X1 port map( G => n2013, D => n1697, Q => 
                           REG_25_20_port);
   REG_reg_25_19_inst : DLH_X1 port map( G => n2012, D => n1703, Q => 
                           REG_25_19_port);
   REG_reg_25_18_inst : DLH_X1 port map( G => n2012, D => n1709, Q => 
                           REG_25_18_port);
   REG_reg_25_17_inst : DLH_X1 port map( G => n2012, D => n1715, Q => 
                           REG_25_17_port);
   REG_reg_25_16_inst : DLH_X1 port map( G => n2012, D => n1721, Q => 
                           REG_25_16_port);
   REG_reg_25_15_inst : DLH_X1 port map( G => n2012, D => n1727, Q => 
                           REG_25_15_port);
   REG_reg_25_14_inst : DLH_X1 port map( G => n2012, D => n1733, Q => 
                           REG_25_14_port);
   REG_reg_25_13_inst : DLH_X1 port map( G => n2012, D => n1739, Q => 
                           REG_25_13_port);
   REG_reg_25_12_inst : DLH_X1 port map( G => n2012, D => n1745, Q => 
                           REG_25_12_port);
   REG_reg_25_11_inst : DLH_X1 port map( G => n2012, D => n1751, Q => 
                           REG_25_11_port);
   REG_reg_25_10_inst : DLH_X1 port map( G => n2012, D => n1757, Q => 
                           REG_25_10_port);
   REG_reg_25_9_inst : DLH_X1 port map( G => n2011, D => n1763, Q => 
                           REG_25_9_port);
   REG_reg_25_8_inst : DLH_X1 port map( G => n2011, D => n1769, Q => 
                           REG_25_8_port);
   REG_reg_25_7_inst : DLH_X1 port map( G => n2011, D => n1775, Q => 
                           REG_25_7_port);
   REG_reg_25_6_inst : DLH_X1 port map( G => n2011, D => n1781, Q => 
                           REG_25_6_port);
   REG_reg_25_5_inst : DLH_X1 port map( G => n2011, D => n1787, Q => 
                           REG_25_5_port);
   REG_reg_25_4_inst : DLH_X1 port map( G => n2011, D => n1793, Q => 
                           REG_25_4_port);
   REG_reg_25_3_inst : DLH_X1 port map( G => n2011, D => n1799, Q => 
                           REG_25_3_port);
   REG_reg_25_2_inst : DLH_X1 port map( G => n2011, D => n1805, Q => 
                           REG_25_2_port);
   REG_reg_25_1_inst : DLH_X1 port map( G => n2011, D => n1811, Q => 
                           REG_25_1_port);
   REG_reg_25_0_inst : DLH_X1 port map( G => n2011, D => n1817, Q => 
                           REG_25_0_port);
   REG_reg_26_31_inst : DLH_X1 port map( G => n2021, D => n1631, Q => 
                           REG_26_31_port);
   REG_reg_26_30_inst : DLH_X1 port map( G => n2021, D => n1637, Q => 
                           REG_26_30_port);
   REG_reg_26_29_inst : DLH_X1 port map( G => n2020, D => n1643, Q => 
                           REG_26_29_port);
   REG_reg_26_28_inst : DLH_X1 port map( G => n2020, D => n1649, Q => 
                           REG_26_28_port);
   REG_reg_26_27_inst : DLH_X1 port map( G => n2020, D => n1655, Q => 
                           REG_26_27_port);
   REG_reg_26_26_inst : DLH_X1 port map( G => n2020, D => n1661, Q => 
                           REG_26_26_port);
   REG_reg_26_25_inst : DLH_X1 port map( G => n2020, D => n1667, Q => 
                           REG_26_25_port);
   REG_reg_26_24_inst : DLH_X1 port map( G => n2020, D => n1673, Q => 
                           REG_26_24_port);
   REG_reg_26_23_inst : DLH_X1 port map( G => n2020, D => n1679, Q => 
                           REG_26_23_port);
   REG_reg_26_22_inst : DLH_X1 port map( G => n2020, D => n1685, Q => 
                           REG_26_22_port);
   REG_reg_26_21_inst : DLH_X1 port map( G => n2020, D => n1691, Q => 
                           REG_26_21_port);
   REG_reg_26_20_inst : DLH_X1 port map( G => n2020, D => n1697, Q => 
                           REG_26_20_port);
   REG_reg_26_19_inst : DLH_X1 port map( G => n2019, D => n1703, Q => 
                           REG_26_19_port);
   REG_reg_26_18_inst : DLH_X1 port map( G => n2019, D => n1709, Q => 
                           REG_26_18_port);
   REG_reg_26_17_inst : DLH_X1 port map( G => n2019, D => n1715, Q => 
                           REG_26_17_port);
   REG_reg_26_16_inst : DLH_X1 port map( G => n2019, D => n1721, Q => 
                           REG_26_16_port);
   REG_reg_26_15_inst : DLH_X1 port map( G => n2019, D => n1727, Q => 
                           REG_26_15_port);
   REG_reg_26_14_inst : DLH_X1 port map( G => n2019, D => n1733, Q => 
                           REG_26_14_port);
   REG_reg_26_13_inst : DLH_X1 port map( G => n2019, D => n1739, Q => 
                           REG_26_13_port);
   REG_reg_26_12_inst : DLH_X1 port map( G => n2019, D => n1745, Q => 
                           REG_26_12_port);
   REG_reg_26_11_inst : DLH_X1 port map( G => n2019, D => n1751, Q => 
                           REG_26_11_port);
   REG_reg_26_10_inst : DLH_X1 port map( G => n2019, D => n1757, Q => 
                           REG_26_10_port);
   REG_reg_26_9_inst : DLH_X1 port map( G => n2018, D => n1763, Q => 
                           REG_26_9_port);
   REG_reg_26_8_inst : DLH_X1 port map( G => n2018, D => n1769, Q => 
                           REG_26_8_port);
   REG_reg_26_7_inst : DLH_X1 port map( G => n2018, D => n1775, Q => 
                           REG_26_7_port);
   REG_reg_26_6_inst : DLH_X1 port map( G => n2018, D => n1781, Q => 
                           REG_26_6_port);
   REG_reg_26_5_inst : DLH_X1 port map( G => n2018, D => n1787, Q => 
                           REG_26_5_port);
   REG_reg_26_4_inst : DLH_X1 port map( G => n2018, D => n1793, Q => 
                           REG_26_4_port);
   REG_reg_26_3_inst : DLH_X1 port map( G => n2018, D => n1799, Q => 
                           REG_26_3_port);
   REG_reg_26_2_inst : DLH_X1 port map( G => n2018, D => n1805, Q => 
                           REG_26_2_port);
   REG_reg_26_1_inst : DLH_X1 port map( G => n2018, D => n1811, Q => 
                           REG_26_1_port);
   REG_reg_26_0_inst : DLH_X1 port map( G => n2018, D => n1817, Q => 
                           REG_26_0_port);
   REG_reg_27_31_inst : DLH_X1 port map( G => n2028, D => n1631, Q => 
                           REG_27_31_port);
   REG_reg_27_30_inst : DLH_X1 port map( G => n2028, D => n1637, Q => 
                           REG_27_30_port);
   REG_reg_27_29_inst : DLH_X1 port map( G => n2027, D => n1643, Q => 
                           REG_27_29_port);
   REG_reg_27_28_inst : DLH_X1 port map( G => n2027, D => n1649, Q => 
                           REG_27_28_port);
   REG_reg_27_27_inst : DLH_X1 port map( G => n2027, D => n1655, Q => 
                           REG_27_27_port);
   REG_reg_27_26_inst : DLH_X1 port map( G => n2027, D => n1661, Q => 
                           REG_27_26_port);
   REG_reg_27_25_inst : DLH_X1 port map( G => n2027, D => n1667, Q => 
                           REG_27_25_port);
   REG_reg_27_24_inst : DLH_X1 port map( G => n2027, D => n1673, Q => 
                           REG_27_24_port);
   REG_reg_27_23_inst : DLH_X1 port map( G => n2027, D => n1679, Q => 
                           REG_27_23_port);
   REG_reg_27_22_inst : DLH_X1 port map( G => n2027, D => n1685, Q => 
                           REG_27_22_port);
   REG_reg_27_21_inst : DLH_X1 port map( G => n2027, D => n1691, Q => 
                           REG_27_21_port);
   REG_reg_27_20_inst : DLH_X1 port map( G => n2027, D => n1697, Q => 
                           REG_27_20_port);
   REG_reg_27_19_inst : DLH_X1 port map( G => n2026, D => n1703, Q => 
                           REG_27_19_port);
   REG_reg_27_18_inst : DLH_X1 port map( G => n2026, D => n1709, Q => 
                           REG_27_18_port);
   REG_reg_27_17_inst : DLH_X1 port map( G => n2026, D => n1715, Q => 
                           REG_27_17_port);
   REG_reg_27_16_inst : DLH_X1 port map( G => n2026, D => n1721, Q => 
                           REG_27_16_port);
   REG_reg_27_15_inst : DLH_X1 port map( G => n2026, D => n1727, Q => 
                           REG_27_15_port);
   REG_reg_27_14_inst : DLH_X1 port map( G => n2026, D => n1733, Q => 
                           REG_27_14_port);
   REG_reg_27_13_inst : DLH_X1 port map( G => n2026, D => n1739, Q => 
                           REG_27_13_port);
   REG_reg_27_12_inst : DLH_X1 port map( G => n2026, D => n1745, Q => 
                           REG_27_12_port);
   REG_reg_27_11_inst : DLH_X1 port map( G => n2026, D => n1751, Q => 
                           REG_27_11_port);
   REG_reg_27_10_inst : DLH_X1 port map( G => n2026, D => n1757, Q => 
                           REG_27_10_port);
   REG_reg_27_9_inst : DLH_X1 port map( G => n2025, D => n1763, Q => 
                           REG_27_9_port);
   REG_reg_27_8_inst : DLH_X1 port map( G => n2025, D => n1769, Q => 
                           REG_27_8_port);
   REG_reg_27_7_inst : DLH_X1 port map( G => n2025, D => n1775, Q => 
                           REG_27_7_port);
   REG_reg_27_6_inst : DLH_X1 port map( G => n2025, D => n1781, Q => 
                           REG_27_6_port);
   REG_reg_27_5_inst : DLH_X1 port map( G => n2025, D => n1787, Q => 
                           REG_27_5_port);
   REG_reg_27_4_inst : DLH_X1 port map( G => n2025, D => n1793, Q => 
                           REG_27_4_port);
   REG_reg_27_3_inst : DLH_X1 port map( G => n2025, D => n1799, Q => 
                           REG_27_3_port);
   REG_reg_27_2_inst : DLH_X1 port map( G => n2025, D => n1805, Q => 
                           REG_27_2_port);
   REG_reg_27_1_inst : DLH_X1 port map( G => n2025, D => n1811, Q => 
                           REG_27_1_port);
   REG_reg_27_0_inst : DLH_X1 port map( G => n2025, D => n1817, Q => 
                           REG_27_0_port);
   REG_reg_28_31_inst : DLH_X1 port map( G => n2035, D => n1631, Q => 
                           REG_28_31_port);
   REG_reg_28_30_inst : DLH_X1 port map( G => n2035, D => n1637, Q => 
                           REG_28_30_port);
   REG_reg_28_29_inst : DLH_X1 port map( G => n2034, D => n1643, Q => 
                           REG_28_29_port);
   REG_reg_28_28_inst : DLH_X1 port map( G => n2034, D => n1649, Q => 
                           REG_28_28_port);
   REG_reg_28_27_inst : DLH_X1 port map( G => n2034, D => n1655, Q => 
                           REG_28_27_port);
   REG_reg_28_26_inst : DLH_X1 port map( G => n2034, D => n1661, Q => 
                           REG_28_26_port);
   REG_reg_28_25_inst : DLH_X1 port map( G => n2034, D => n1667, Q => 
                           REG_28_25_port);
   REG_reg_28_24_inst : DLH_X1 port map( G => n2034, D => n1673, Q => 
                           REG_28_24_port);
   REG_reg_28_23_inst : DLH_X1 port map( G => n2034, D => n1679, Q => 
                           REG_28_23_port);
   REG_reg_28_22_inst : DLH_X1 port map( G => n2034, D => n1685, Q => 
                           REG_28_22_port);
   REG_reg_28_21_inst : DLH_X1 port map( G => n2034, D => n1691, Q => 
                           REG_28_21_port);
   REG_reg_28_20_inst : DLH_X1 port map( G => n2034, D => n1697, Q => 
                           REG_28_20_port);
   REG_reg_28_19_inst : DLH_X1 port map( G => n2033, D => n1703, Q => 
                           REG_28_19_port);
   REG_reg_28_18_inst : DLH_X1 port map( G => n2033, D => n1709, Q => 
                           REG_28_18_port);
   REG_reg_28_17_inst : DLH_X1 port map( G => n2033, D => n1715, Q => 
                           REG_28_17_port);
   REG_reg_28_16_inst : DLH_X1 port map( G => n2033, D => n1721, Q => 
                           REG_28_16_port);
   REG_reg_28_15_inst : DLH_X1 port map( G => n2033, D => n1727, Q => 
                           REG_28_15_port);
   REG_reg_28_14_inst : DLH_X1 port map( G => n2033, D => n1733, Q => 
                           REG_28_14_port);
   REG_reg_28_13_inst : DLH_X1 port map( G => n2033, D => n1739, Q => 
                           REG_28_13_port);
   REG_reg_28_12_inst : DLH_X1 port map( G => n2033, D => n1745, Q => 
                           REG_28_12_port);
   REG_reg_28_11_inst : DLH_X1 port map( G => n2033, D => n1751, Q => 
                           REG_28_11_port);
   REG_reg_28_10_inst : DLH_X1 port map( G => n2033, D => n1757, Q => 
                           REG_28_10_port);
   REG_reg_28_9_inst : DLH_X1 port map( G => n2032, D => n1763, Q => 
                           REG_28_9_port);
   REG_reg_28_8_inst : DLH_X1 port map( G => n2032, D => n1769, Q => 
                           REG_28_8_port);
   REG_reg_28_7_inst : DLH_X1 port map( G => n2032, D => n1775, Q => 
                           REG_28_7_port);
   REG_reg_28_6_inst : DLH_X1 port map( G => n2032, D => n1781, Q => 
                           REG_28_6_port);
   REG_reg_28_5_inst : DLH_X1 port map( G => n2032, D => n1787, Q => 
                           REG_28_5_port);
   REG_reg_28_4_inst : DLH_X1 port map( G => n2032, D => n1793, Q => 
                           REG_28_4_port);
   REG_reg_28_3_inst : DLH_X1 port map( G => n2032, D => n1799, Q => 
                           REG_28_3_port);
   REG_reg_28_2_inst : DLH_X1 port map( G => n2032, D => n1805, Q => 
                           REG_28_2_port);
   REG_reg_28_1_inst : DLH_X1 port map( G => n2032, D => n1811, Q => 
                           REG_28_1_port);
   REG_reg_28_0_inst : DLH_X1 port map( G => n2032, D => n1817, Q => 
                           REG_28_0_port);
   REG_reg_29_31_inst : DLH_X1 port map( G => n2042, D => n1631, Q => 
                           REG_29_31_port);
   REG_reg_29_30_inst : DLH_X1 port map( G => n2042, D => n1637, Q => 
                           REG_29_30_port);
   REG_reg_29_29_inst : DLH_X1 port map( G => n2041, D => n1643, Q => 
                           REG_29_29_port);
   REG_reg_29_28_inst : DLH_X1 port map( G => n2041, D => n1649, Q => 
                           REG_29_28_port);
   REG_reg_29_27_inst : DLH_X1 port map( G => n2041, D => n1655, Q => 
                           REG_29_27_port);
   REG_reg_29_26_inst : DLH_X1 port map( G => n2041, D => n1661, Q => 
                           REG_29_26_port);
   REG_reg_29_25_inst : DLH_X1 port map( G => n2041, D => n1667, Q => 
                           REG_29_25_port);
   REG_reg_29_24_inst : DLH_X1 port map( G => n2041, D => n1673, Q => 
                           REG_29_24_port);
   REG_reg_29_23_inst : DLH_X1 port map( G => n2041, D => n1679, Q => 
                           REG_29_23_port);
   REG_reg_29_22_inst : DLH_X1 port map( G => n2041, D => n1685, Q => 
                           REG_29_22_port);
   REG_reg_29_21_inst : DLH_X1 port map( G => n2041, D => n1691, Q => 
                           REG_29_21_port);
   REG_reg_29_20_inst : DLH_X1 port map( G => n2041, D => n1697, Q => 
                           REG_29_20_port);
   REG_reg_29_19_inst : DLH_X1 port map( G => n2040, D => n1703, Q => 
                           REG_29_19_port);
   REG_reg_29_18_inst : DLH_X1 port map( G => n2040, D => n1709, Q => 
                           REG_29_18_port);
   REG_reg_29_17_inst : DLH_X1 port map( G => n2040, D => n1715, Q => 
                           REG_29_17_port);
   REG_reg_29_16_inst : DLH_X1 port map( G => n2040, D => n1721, Q => 
                           REG_29_16_port);
   REG_reg_29_15_inst : DLH_X1 port map( G => n2040, D => n1727, Q => 
                           REG_29_15_port);
   REG_reg_29_14_inst : DLH_X1 port map( G => n2040, D => n1733, Q => 
                           REG_29_14_port);
   REG_reg_29_13_inst : DLH_X1 port map( G => n2040, D => n1739, Q => 
                           REG_29_13_port);
   REG_reg_29_12_inst : DLH_X1 port map( G => n2040, D => n1745, Q => 
                           REG_29_12_port);
   REG_reg_29_11_inst : DLH_X1 port map( G => n2040, D => n1751, Q => 
                           REG_29_11_port);
   REG_reg_29_10_inst : DLH_X1 port map( G => n2040, D => n1757, Q => 
                           REG_29_10_port);
   REG_reg_29_9_inst : DLH_X1 port map( G => n2039, D => n1763, Q => 
                           REG_29_9_port);
   REG_reg_29_8_inst : DLH_X1 port map( G => n2039, D => n1769, Q => 
                           REG_29_8_port);
   REG_reg_29_7_inst : DLH_X1 port map( G => n2039, D => n1775, Q => 
                           REG_29_7_port);
   REG_reg_29_6_inst : DLH_X1 port map( G => n2039, D => n1781, Q => 
                           REG_29_6_port);
   REG_reg_29_5_inst : DLH_X1 port map( G => n2039, D => n1787, Q => 
                           REG_29_5_port);
   REG_reg_29_4_inst : DLH_X1 port map( G => n2039, D => n1793, Q => 
                           REG_29_4_port);
   REG_reg_29_3_inst : DLH_X1 port map( G => n2039, D => n1799, Q => 
                           REG_29_3_port);
   REG_reg_29_2_inst : DLH_X1 port map( G => n2039, D => n1805, Q => 
                           REG_29_2_port);
   REG_reg_29_1_inst : DLH_X1 port map( G => n2039, D => n1811, Q => 
                           REG_29_1_port);
   REG_reg_29_0_inst : DLH_X1 port map( G => n2039, D => n1817, Q => 
                           REG_29_0_port);
   REG_reg_30_31_inst : DLH_X1 port map( G => n2049, D => n1631, Q => 
                           REG_30_31_port);
   REG_reg_30_30_inst : DLH_X1 port map( G => n2049, D => n1637, Q => 
                           REG_30_30_port);
   REG_reg_30_29_inst : DLH_X1 port map( G => n2048, D => n1643, Q => 
                           REG_30_29_port);
   REG_reg_30_28_inst : DLH_X1 port map( G => n2048, D => n1649, Q => 
                           REG_30_28_port);
   REG_reg_30_27_inst : DLH_X1 port map( G => n2048, D => n1655, Q => 
                           REG_30_27_port);
   REG_reg_30_26_inst : DLH_X1 port map( G => n2048, D => n1661, Q => 
                           REG_30_26_port);
   REG_reg_30_25_inst : DLH_X1 port map( G => n2048, D => n1667, Q => 
                           REG_30_25_port);
   REG_reg_30_24_inst : DLH_X1 port map( G => n2048, D => n1673, Q => 
                           REG_30_24_port);
   REG_reg_30_23_inst : DLH_X1 port map( G => n2048, D => n1679, Q => 
                           REG_30_23_port);
   REG_reg_30_22_inst : DLH_X1 port map( G => n2048, D => n1685, Q => 
                           REG_30_22_port);
   REG_reg_30_21_inst : DLH_X1 port map( G => n2048, D => n1691, Q => 
                           REG_30_21_port);
   REG_reg_30_20_inst : DLH_X1 port map( G => n2048, D => n1697, Q => 
                           REG_30_20_port);
   REG_reg_30_19_inst : DLH_X1 port map( G => n2047, D => n1703, Q => 
                           REG_30_19_port);
   REG_reg_30_18_inst : DLH_X1 port map( G => n2047, D => n1709, Q => 
                           REG_30_18_port);
   REG_reg_30_17_inst : DLH_X1 port map( G => n2047, D => n1715, Q => 
                           REG_30_17_port);
   REG_reg_30_16_inst : DLH_X1 port map( G => n2047, D => n1721, Q => 
                           REG_30_16_port);
   REG_reg_30_15_inst : DLH_X1 port map( G => n2047, D => n1727, Q => 
                           REG_30_15_port);
   REG_reg_30_14_inst : DLH_X1 port map( G => n2047, D => n1733, Q => 
                           REG_30_14_port);
   REG_reg_30_13_inst : DLH_X1 port map( G => n2047, D => n1739, Q => 
                           REG_30_13_port);
   REG_reg_30_12_inst : DLH_X1 port map( G => n2047, D => n1745, Q => 
                           REG_30_12_port);
   REG_reg_30_11_inst : DLH_X1 port map( G => n2047, D => n1751, Q => 
                           REG_30_11_port);
   REG_reg_30_10_inst : DLH_X1 port map( G => n2047, D => n1757, Q => 
                           REG_30_10_port);
   REG_reg_30_9_inst : DLH_X1 port map( G => n2046, D => n1763, Q => 
                           REG_30_9_port);
   REG_reg_30_8_inst : DLH_X1 port map( G => n2046, D => n1769, Q => 
                           REG_30_8_port);
   REG_reg_30_7_inst : DLH_X1 port map( G => n2046, D => n1775, Q => 
                           REG_30_7_port);
   REG_reg_30_6_inst : DLH_X1 port map( G => n2046, D => n1781, Q => 
                           REG_30_6_port);
   REG_reg_30_5_inst : DLH_X1 port map( G => n2046, D => n1787, Q => 
                           REG_30_5_port);
   REG_reg_30_4_inst : DLH_X1 port map( G => n2046, D => n1793, Q => 
                           REG_30_4_port);
   REG_reg_30_3_inst : DLH_X1 port map( G => n2046, D => n1799, Q => 
                           REG_30_3_port);
   REG_reg_30_2_inst : DLH_X1 port map( G => n2046, D => n1805, Q => 
                           REG_30_2_port);
   REG_reg_30_1_inst : DLH_X1 port map( G => n2046, D => n1811, Q => 
                           REG_30_1_port);
   REG_reg_30_0_inst : DLH_X1 port map( G => n2046, D => n1817, Q => 
                           REG_30_0_port);
   REG_reg_31_31_inst : DLH_X1 port map( G => n2056, D => n2061, Q => 
                           REG_31_31_port);
   REG_reg_31_30_inst : DLH_X1 port map( G => n2056, D => n2062, Q => 
                           REG_31_30_port);
   REG_reg_31_29_inst : DLH_X1 port map( G => n2055, D => n2063, Q => 
                           REG_31_29_port);
   REG_reg_31_28_inst : DLH_X1 port map( G => n2055, D => n2064, Q => 
                           REG_31_28_port);
   REG_reg_31_27_inst : DLH_X1 port map( G => n2055, D => n2065, Q => 
                           REG_31_27_port);
   REG_reg_31_26_inst : DLH_X1 port map( G => n2055, D => n2066, Q => 
                           REG_31_26_port);
   REG_reg_31_25_inst : DLH_X1 port map( G => n2055, D => n2067, Q => 
                           REG_31_25_port);
   REG_reg_31_24_inst : DLH_X1 port map( G => n2055, D => n2068, Q => 
                           REG_31_24_port);
   REG_reg_31_23_inst : DLH_X1 port map( G => n2055, D => n2069, Q => 
                           REG_31_23_port);
   REG_reg_31_22_inst : DLH_X1 port map( G => n2055, D => n2070, Q => 
                           REG_31_22_port);
   REG_reg_31_21_inst : DLH_X1 port map( G => n2055, D => n2071, Q => 
                           REG_31_21_port);
   REG_reg_31_20_inst : DLH_X1 port map( G => n2055, D => n2072, Q => 
                           REG_31_20_port);
   REG_reg_31_19_inst : DLH_X1 port map( G => n2054, D => n2073, Q => 
                           REG_31_19_port);
   REG_reg_31_18_inst : DLH_X1 port map( G => n2054, D => n2074, Q => 
                           REG_31_18_port);
   REG_reg_31_17_inst : DLH_X1 port map( G => n2054, D => n2075, Q => 
                           REG_31_17_port);
   REG_reg_31_16_inst : DLH_X1 port map( G => n2054, D => n2076, Q => 
                           REG_31_16_port);
   REG_reg_31_15_inst : DLH_X1 port map( G => n2054, D => n2077, Q => 
                           REG_31_15_port);
   REG_reg_31_14_inst : DLH_X1 port map( G => n2054, D => n2078, Q => 
                           REG_31_14_port);
   REG_reg_31_13_inst : DLH_X1 port map( G => n2054, D => n2079, Q => 
                           REG_31_13_port);
   REG_reg_31_12_inst : DLH_X1 port map( G => n2054, D => n2080, Q => 
                           REG_31_12_port);
   REG_reg_31_11_inst : DLH_X1 port map( G => n2054, D => n2081, Q => 
                           REG_31_11_port);
   REG_reg_31_10_inst : DLH_X1 port map( G => n2054, D => n2082, Q => 
                           REG_31_10_port);
   REG_reg_31_9_inst : DLH_X1 port map( G => n2053, D => n2083, Q => 
                           REG_31_9_port);
   REG_reg_31_8_inst : DLH_X1 port map( G => n2053, D => n2084, Q => 
                           REG_31_8_port);
   REG_reg_31_7_inst : DLH_X1 port map( G => n2053, D => n2085, Q => 
                           REG_31_7_port);
   REG_reg_31_6_inst : DLH_X1 port map( G => n2053, D => n2086, Q => 
                           REG_31_6_port);
   REG_reg_31_5_inst : DLH_X1 port map( G => n2053, D => n2087, Q => 
                           REG_31_5_port);
   REG_reg_31_4_inst : DLH_X1 port map( G => n2053, D => n2088, Q => 
                           REG_31_4_port);
   REG_reg_31_3_inst : DLH_X1 port map( G => n2053, D => n2089, Q => 
                           REG_31_3_port);
   REG_reg_31_2_inst : DLH_X1 port map( G => n2053, D => n2090, Q => 
                           REG_31_2_port);
   REG_reg_31_1_inst : DLH_X1 port map( G => n2053, D => n2091, Q => 
                           REG_31_1_port);
   REG_reg_31_0_inst : DLH_X1 port map( G => n2053, D => n2092, Q => 
                           REG_31_0_port);
   OUT2_reg_31_inst : DLH_X1 port map( G => n1824, D => N284, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => n1824, D => N285, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => n1824, D => N286, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => n1824, D => N287, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => n1824, D => N288, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => n1824, D => N289, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => n1824, D => N290, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => n1824, D => N291, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => n1824, D => N292, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => n1824, D => N293, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => n1825, D => N294, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => n1825, D => N295, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => n1825, D => N296, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => n1825, D => N297, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => n1825, D => N298, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => n1825, D => N299, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => n1825, D => N300, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => n1825, D => N301, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => n1825, D => N302, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => n1825, D => N303, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => n1826, D => N304, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => n1826, D => N305, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => n1826, D => N306, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => n1826, D => N307, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => n1826, D => N308, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => n1826, D => N309, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => n1826, D => N310, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => n1826, D => N311, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => n1826, D => N312, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => n1826, D => N313, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => n1827, D => N314, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => n1827, D => N315, Q => OUT2(0));
   OUT1_reg_31_inst : DLH_X1 port map( G => n1830, D => N252, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => n1830, D => N253, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => n1830, D => N254, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => n1830, D => N255, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => n1830, D => N256, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => n1830, D => N257, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => n1830, D => N258, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => n1830, D => N259, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => n1830, D => N260, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => n1830, D => N261, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => n1831, D => N262, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => n1831, D => N263, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => n1831, D => N264, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => n1831, D => N265, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => n1831, D => N266, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => n1831, D => N267, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => n1831, D => N268, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => n1831, D => N269, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => n1831, D => N270, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => n1831, D => N271, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => n1832, D => N272, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => n1832, D => N273, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => n1832, D => N274, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => n1832, D => N275, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => n1832, D => N276, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => n1832, D => N277, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => n1832, D => N278, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => n1832, D => N279, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => n1832, D => N280, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => n1832, D => N281, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => n1833, D => N282, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => n1833, D => N283, Q => OUT1(0));
   U142 : NAND3_X1 port map( A1 => n2094, A2 => n2093, A3 => n2060, ZN => n75);
   U143 : NAND3_X1 port map( A1 => n2060, A2 => n2093, A3 => ADD_WR(3), ZN => 
                           n83);
   U144 : NAND3_X1 port map( A1 => n2060, A2 => n2094, A3 => ADD_WR(4), ZN => 
                           n84);
   U145 : NAND3_X1 port map( A1 => n2096, A2 => n2095, A3 => n2097, ZN => n74);
   U146 : NAND3_X1 port map( A1 => n2096, A2 => n2095, A3 => ADD_WR(0), ZN => 
                           n76);
   U147 : NAND3_X1 port map( A1 => n2097, A2 => n2095, A3 => ADD_WR(1), ZN => 
                           n77);
   U148 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2095, A3 => ADD_WR(1), ZN 
                           => n78);
   U149 : NAND3_X1 port map( A1 => n2097, A2 => n2096, A3 => ADD_WR(2), ZN => 
                           n79);
   U150 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2096, A3 => ADD_WR(2), ZN 
                           => n80);
   U151 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n2097, A3 => ADD_WR(2), ZN 
                           => n81);
   U152 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n2060, A3 => ADD_WR(4), ZN 
                           => n85);
   U153 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2),
                           ZN => n82);
   U3 : BUF_X2 port map( A => n8, Z => n1611);
   U4 : AND2_X4 port map( A1 => n912, A2 => n1592, ZN => n8);
   U5 : BUF_X2 port map( A => n5, Z => n1599);
   U6 : AND2_X4 port map( A1 => n912, A2 => ADD_RD2(0), ZN => n5);
   U7 : AND2_X2 port map( A1 => n911, A2 => n1592, ZN => n9);
   U8 : BUF_X2 port map( A => n6, Z => n1601);
   U9 : BUF_X2 port map( A => n6, Z => n1602);
   U10 : AND2_X2 port map( A1 => n911, A2 => ADD_RD2(0), ZN => n6);
   U11 : CLKBUF_X3 port map( A => n7, Z => n1610);
   U12 : AND2_X4 port map( A1 => n909, A2 => n1592, ZN => n7);
   U13 : CLKBUF_X3 port map( A => n4, Z => n1598);
   U14 : AND2_X4 port map( A1 => n909, A2 => ADD_RD2(0), ZN => n4);
   U15 : BUF_X2 port map( A => n3, Z => n1605);
   U16 : AND2_X2 port map( A1 => n910, A2 => n1592, ZN => n3);
   U17 : BUF_X2 port map( A => n2, Z => n1593);
   U18 : AND2_X2 port map( A1 => ADD_RD2(0), A2 => n910, ZN => n2);
   U19 : BUF_X2 port map( A => n1583, Z => n1619);
   U20 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n1585);
   U21 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => n1589, ZN => n1587);
   U22 : NOR2_X2 port map( A1 => n1589, A2 => ADD_RD2(4), ZN => n1581);
   U23 : OR3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(4), A3 => n74, ZN => n1
                           );
   U24 : AND2_X1 port map( A1 => n21, A2 => n748, ZN => n10);
   U25 : AND2_X1 port map( A1 => n20, A2 => n748, ZN => n11);
   U26 : AND2_X1 port map( A1 => n23, A2 => n748, ZN => n12);
   U27 : AND2_X1 port map( A1 => n22, A2 => n748, ZN => n13);
   U28 : AND2_X1 port map( A1 => EN_RD1, A2 => EN, ZN => n14);
   U29 : AND2_X1 port map( A1 => EN_RD2, A2 => EN, ZN => n15);
   U30 : BUF_X1 port map( A => n1620, Z => n1628);
   U31 : BUF_X1 port map( A => n1620, Z => n1627);
   U32 : BUF_X1 port map( A => n876, Z => n877);
   U33 : BUF_X1 port map( A => n858, Z => n859);
   U34 : BUF_X1 port map( A => n876, Z => n878);
   U35 : BUF_X1 port map( A => n858, Z => n860);
   U36 : BUF_X1 port map( A => n876, Z => n879);
   U37 : BUF_X1 port map( A => n858, Z => n861);
   U38 : BUF_X1 port map( A => n840, Z => n841);
   U39 : BUF_X1 port map( A => n822, Z => n823);
   U40 : BUF_X1 port map( A => n840, Z => n842);
   U41 : BUF_X1 port map( A => n822, Z => n824);
   U42 : BUF_X1 port map( A => n840, Z => n843);
   U43 : BUF_X1 port map( A => n822, Z => n825);
   U44 : BUF_X1 port map( A => n13, Z => n876);
   U45 : BUF_X1 port map( A => n12, Z => n858);
   U46 : BUF_X1 port map( A => n11, Z => n840);
   U47 : BUF_X1 port map( A => n10, Z => n822);
   U48 : BUF_X1 port map( A => n804, Z => n805);
   U49 : BUF_X1 port map( A => n786, Z => n787);
   U50 : BUF_X1 port map( A => n768, Z => n769);
   U51 : BUF_X1 port map( A => n750, Z => n751);
   U52 : BUF_X1 port map( A => n804, Z => n806);
   U53 : BUF_X1 port map( A => n786, Z => n788);
   U54 : BUF_X1 port map( A => n768, Z => n770);
   U55 : BUF_X1 port map( A => n750, Z => n752);
   U56 : BUF_X1 port map( A => n804, Z => n807);
   U57 : BUF_X1 port map( A => n786, Z => n789);
   U58 : BUF_X1 port map( A => n768, Z => n771);
   U59 : BUF_X1 port map( A => n750, Z => n753);
   U60 : BUF_X1 port map( A => n1820, Z => n1818);
   U61 : BUF_X1 port map( A => n1814, Z => n1812);
   U62 : BUF_X1 port map( A => n1808, Z => n1806);
   U63 : BUF_X1 port map( A => n1802, Z => n1800);
   U64 : BUF_X1 port map( A => n1796, Z => n1794);
   U65 : BUF_X1 port map( A => n1790, Z => n1788);
   U66 : BUF_X1 port map( A => n1784, Z => n1782);
   U67 : BUF_X1 port map( A => n1778, Z => n1776);
   U68 : BUF_X1 port map( A => n1772, Z => n1770);
   U69 : BUF_X1 port map( A => n1766, Z => n1764);
   U70 : BUF_X1 port map( A => n1760, Z => n1758);
   U71 : BUF_X1 port map( A => n1754, Z => n1752);
   U72 : BUF_X1 port map( A => n1748, Z => n1746);
   U73 : BUF_X1 port map( A => n1742, Z => n1740);
   U74 : BUF_X1 port map( A => n1736, Z => n1734);
   U75 : BUF_X1 port map( A => n1730, Z => n1728);
   U76 : BUF_X1 port map( A => n1724, Z => n1722);
   U77 : BUF_X1 port map( A => n1718, Z => n1716);
   U78 : BUF_X1 port map( A => n1712, Z => n1710);
   U79 : BUF_X1 port map( A => n1706, Z => n1704);
   U80 : BUF_X1 port map( A => n1700, Z => n1698);
   U81 : BUF_X1 port map( A => n1694, Z => n1692);
   U82 : BUF_X1 port map( A => n1688, Z => n1686);
   U83 : BUF_X1 port map( A => n1682, Z => n1680);
   U84 : BUF_X1 port map( A => n1676, Z => n1674);
   U85 : BUF_X1 port map( A => n1670, Z => n1668);
   U86 : BUF_X1 port map( A => n1664, Z => n1662);
   U87 : BUF_X1 port map( A => n1658, Z => n1656);
   U88 : BUF_X1 port map( A => n1652, Z => n1650);
   U89 : BUF_X1 port map( A => n1646, Z => n1644);
   U90 : BUF_X1 port map( A => n1640, Z => n1638);
   U91 : BUF_X1 port map( A => n1634, Z => n1632);
   U92 : BUF_X1 port map( A => n875, Z => n880);
   U93 : BUF_X1 port map( A => n857, Z => n862);
   U94 : BUF_X1 port map( A => n839, Z => n844);
   U95 : BUF_X1 port map( A => n821, Z => n826);
   U96 : BUF_X1 port map( A => n16, Z => n804);
   U97 : BUF_X1 port map( A => n17, Z => n786);
   U98 : BUF_X1 port map( A => n18, Z => n768);
   U99 : BUF_X1 port map( A => n19, Z => n750);
   U100 : BUF_X1 port map( A => n2059, Z => n2057);
   U101 : BUF_X1 port map( A => n2052, Z => n2050);
   U102 : BUF_X1 port map( A => n2045, Z => n2043);
   U103 : BUF_X1 port map( A => n2038, Z => n2036);
   U104 : BUF_X1 port map( A => n2031, Z => n2029);
   U105 : BUF_X1 port map( A => n2024, Z => n2022);
   U106 : BUF_X1 port map( A => n2017, Z => n2015);
   U107 : BUF_X1 port map( A => n2010, Z => n2008);
   U108 : BUF_X1 port map( A => n2003, Z => n2001);
   U109 : BUF_X1 port map( A => n1996, Z => n1994);
   U110 : BUF_X1 port map( A => n1989, Z => n1987);
   U111 : BUF_X1 port map( A => n1982, Z => n1980);
   U112 : BUF_X1 port map( A => n1975, Z => n1973);
   U113 : BUF_X1 port map( A => n1968, Z => n1966);
   U114 : BUF_X1 port map( A => n1961, Z => n1959);
   U115 : BUF_X1 port map( A => n1954, Z => n1952);
   U116 : BUF_X1 port map( A => n1947, Z => n1945);
   U117 : BUF_X1 port map( A => n1940, Z => n1938);
   U118 : BUF_X1 port map( A => n1933, Z => n1931);
   U119 : BUF_X1 port map( A => n1926, Z => n1924);
   U120 : BUF_X1 port map( A => n1919, Z => n1917);
   U121 : BUF_X1 port map( A => n1912, Z => n1910);
   U122 : BUF_X1 port map( A => n1905, Z => n1903);
   U123 : BUF_X1 port map( A => n1898, Z => n1896);
   U124 : BUF_X1 port map( A => n1891, Z => n1889);
   U125 : BUF_X1 port map( A => n1884, Z => n1882);
   U126 : BUF_X1 port map( A => n1877, Z => n1875);
   U127 : BUF_X1 port map( A => n1870, Z => n1868);
   U128 : BUF_X1 port map( A => n1863, Z => n1861);
   U129 : BUF_X1 port map( A => n1856, Z => n1854);
   U130 : BUF_X1 port map( A => n1849, Z => n1847);
   U131 : BUF_X1 port map( A => n1842, Z => n1840);
   U132 : BUF_X1 port map( A => n803, Z => n808);
   U133 : BUF_X1 port map( A => n785, Z => n790);
   U134 : BUF_X1 port map( A => n767, Z => n772);
   U135 : BUF_X1 port map( A => n749, Z => n754);
   U136 : BUF_X1 port map( A => n739, Z => n897);
   U137 : BUF_X1 port map( A => n737, Z => n893);
   U138 : BUF_X1 port map( A => n741, Z => n901);
   U139 : BUF_X1 port map( A => n743, Z => n905);
   U140 : AND2_X1 port map( A1 => n22, A2 => ADD_RD1(0), ZN => n16);
   U141 : AND2_X1 port map( A1 => n23, A2 => ADD_RD1(0), ZN => n17);
   U154 : AND2_X1 port map( A1 => n20, A2 => ADD_RD1(0), ZN => n18);
   U155 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n21, ZN => n19);
   U156 : BUF_X1 port map( A => n1, Z => n1823);
   U157 : BUF_X1 port map( A => n14, Z => n1834);
   U158 : BUF_X1 port map( A => n15, Z => n1828);
   U159 : BUF_X1 port map( A => n9, Z => n1617);
   U160 : BUF_X1 port map( A => n9, Z => n1615);
   U161 : BUF_X1 port map( A => n9, Z => n1614);
   U162 : BUF_X1 port map( A => n9, Z => n1616);
   U163 : BUF_X1 port map( A => n3, Z => n1609);
   U164 : BUF_X1 port map( A => n6, Z => n1604);
   U165 : BUF_X1 port map( A => n6, Z => n1603);
   U166 : BUF_X1 port map( A => n5, Z => n1600);
   U167 : BUF_X1 port map( A => n2, Z => n1597);
   U168 : BUF_X1 port map( A => n2, Z => n1596);
   U169 : BUF_X1 port map( A => n3, Z => n1608);
   U170 : BUF_X1 port map( A => n3, Z => n1607);
   U171 : BUF_X1 port map( A => n1612, Z => n1613);
   U172 : BUF_X1 port map( A => n3, Z => n1606);
   U173 : BUF_X1 port map( A => n9, Z => n1612);
   U174 : BUF_X1 port map( A => n1628, Z => n1621);
   U175 : BUF_X1 port map( A => n1628, Z => n1622);
   U176 : BUF_X1 port map( A => n1628, Z => n1623);
   U177 : BUF_X1 port map( A => n1627, Z => n1624);
   U178 : BUF_X1 port map( A => n1627, Z => n1625);
   U179 : BUF_X1 port map( A => n877, Z => n892);
   U180 : BUF_X1 port map( A => n878, Z => n889);
   U181 : BUF_X1 port map( A => n878, Z => n888);
   U182 : BUF_X1 port map( A => n879, Z => n885);
   U183 : BUF_X1 port map( A => n879, Z => n884);
   U184 : BUF_X1 port map( A => n841, Z => n856);
   U185 : BUF_X1 port map( A => n877, Z => n891);
   U186 : BUF_X1 port map( A => n841, Z => n855);
   U187 : BUF_X1 port map( A => n877, Z => n890);
   U188 : BUF_X1 port map( A => n841, Z => n854);
   U189 : BUF_X1 port map( A => n842, Z => n853);
   U190 : BUF_X1 port map( A => n842, Z => n852);
   U191 : BUF_X1 port map( A => n878, Z => n887);
   U192 : BUF_X1 port map( A => n842, Z => n851);
   U193 : BUF_X1 port map( A => n879, Z => n886);
   U194 : BUF_X1 port map( A => n843, Z => n850);
   U195 : BUF_X1 port map( A => n843, Z => n849);
   U196 : BUF_X1 port map( A => n843, Z => n848);
   U197 : BUF_X1 port map( A => n859, Z => n874);
   U198 : BUF_X1 port map( A => n860, Z => n871);
   U199 : BUF_X1 port map( A => n860, Z => n870);
   U200 : BUF_X1 port map( A => n861, Z => n867);
   U201 : BUF_X1 port map( A => n861, Z => n866);
   U202 : BUF_X1 port map( A => n823, Z => n838);
   U203 : BUF_X1 port map( A => n859, Z => n873);
   U204 : BUF_X1 port map( A => n823, Z => n837);
   U205 : BUF_X1 port map( A => n859, Z => n872);
   U206 : BUF_X1 port map( A => n823, Z => n836);
   U207 : BUF_X1 port map( A => n824, Z => n835);
   U208 : BUF_X1 port map( A => n824, Z => n834);
   U209 : BUF_X1 port map( A => n860, Z => n869);
   U210 : BUF_X1 port map( A => n824, Z => n833);
   U211 : BUF_X1 port map( A => n861, Z => n868);
   U212 : BUF_X1 port map( A => n825, Z => n832);
   U213 : BUF_X1 port map( A => n825, Z => n831);
   U214 : BUF_X1 port map( A => n825, Z => n830);
   U215 : BUF_X1 port map( A => n2, Z => n1595);
   U216 : BUF_X1 port map( A => n2, Z => n1594);
   U217 : BUF_X1 port map( A => n1627, Z => n1626);
   U218 : BUF_X1 port map( A => n1581, Z => n1618);
   U219 : BUF_X1 port map( A => n805, Z => n820);
   U220 : BUF_X1 port map( A => n769, Z => n784);
   U221 : BUF_X1 port map( A => n805, Z => n819);
   U222 : BUF_X1 port map( A => n769, Z => n783);
   U223 : BUF_X1 port map( A => n805, Z => n818);
   U224 : BUF_X1 port map( A => n769, Z => n782);
   U225 : BUF_X1 port map( A => n806, Z => n817);
   U226 : BUF_X1 port map( A => n770, Z => n781);
   U227 : BUF_X1 port map( A => n806, Z => n816);
   U228 : BUF_X1 port map( A => n770, Z => n780);
   U229 : BUF_X1 port map( A => n806, Z => n815);
   U230 : BUF_X1 port map( A => n770, Z => n779);
   U231 : BUF_X1 port map( A => n807, Z => n814);
   U232 : BUF_X1 port map( A => n771, Z => n778);
   U233 : BUF_X1 port map( A => n807, Z => n813);
   U234 : BUF_X1 port map( A => n771, Z => n777);
   U235 : BUF_X1 port map( A => n807, Z => n812);
   U236 : BUF_X1 port map( A => n771, Z => n776);
   U237 : BUF_X1 port map( A => n880, Z => n883);
   U238 : BUF_X1 port map( A => n844, Z => n847);
   U239 : BUF_X1 port map( A => n880, Z => n882);
   U240 : BUF_X1 port map( A => n844, Z => n846);
   U241 : BUF_X1 port map( A => n787, Z => n802);
   U242 : BUF_X1 port map( A => n751, Z => n766);
   U243 : BUF_X1 port map( A => n787, Z => n801);
   U244 : BUF_X1 port map( A => n751, Z => n765);
   U245 : BUF_X1 port map( A => n787, Z => n800);
   U246 : BUF_X1 port map( A => n751, Z => n764);
   U247 : BUF_X1 port map( A => n788, Z => n799);
   U248 : BUF_X1 port map( A => n752, Z => n763);
   U249 : BUF_X1 port map( A => n788, Z => n798);
   U250 : BUF_X1 port map( A => n752, Z => n762);
   U251 : BUF_X1 port map( A => n788, Z => n797);
   U252 : BUF_X1 port map( A => n752, Z => n761);
   U253 : BUF_X1 port map( A => n789, Z => n796);
   U254 : BUF_X1 port map( A => n753, Z => n760);
   U255 : BUF_X1 port map( A => n789, Z => n795);
   U256 : BUF_X1 port map( A => n753, Z => n759);
   U257 : BUF_X1 port map( A => n789, Z => n794);
   U258 : BUF_X1 port map( A => n753, Z => n758);
   U259 : BUF_X1 port map( A => n862, Z => n865);
   U260 : BUF_X1 port map( A => n826, Z => n829);
   U261 : BUF_X1 port map( A => n862, Z => n864);
   U262 : BUF_X1 port map( A => n826, Z => n828);
   U263 : BUF_X1 port map( A => n880, Z => n881);
   U264 : BUF_X1 port map( A => n844, Z => n845);
   U265 : BUF_X1 port map( A => n1818, Z => n1817);
   U266 : BUF_X1 port map( A => n1812, Z => n1811);
   U267 : BUF_X1 port map( A => n1806, Z => n1805);
   U268 : BUF_X1 port map( A => n1800, Z => n1799);
   U269 : BUF_X1 port map( A => n1794, Z => n1793);
   U270 : BUF_X1 port map( A => n1788, Z => n1787);
   U271 : BUF_X1 port map( A => n1782, Z => n1781);
   U272 : BUF_X1 port map( A => n1776, Z => n1775);
   U273 : BUF_X1 port map( A => n1770, Z => n1769);
   U274 : BUF_X1 port map( A => n1764, Z => n1763);
   U275 : BUF_X1 port map( A => n1758, Z => n1757);
   U276 : BUF_X1 port map( A => n1752, Z => n1751);
   U277 : BUF_X1 port map( A => n1746, Z => n1745);
   U278 : BUF_X1 port map( A => n1740, Z => n1739);
   U279 : BUF_X1 port map( A => n1734, Z => n1733);
   U280 : BUF_X1 port map( A => n1728, Z => n1727);
   U281 : BUF_X1 port map( A => n1722, Z => n1721);
   U282 : BUF_X1 port map( A => n1716, Z => n1715);
   U283 : BUF_X1 port map( A => n1710, Z => n1709);
   U284 : BUF_X1 port map( A => n1704, Z => n1703);
   U285 : BUF_X1 port map( A => n1698, Z => n1697);
   U286 : BUF_X1 port map( A => n1692, Z => n1691);
   U287 : BUF_X1 port map( A => n1686, Z => n1685);
   U288 : BUF_X1 port map( A => n1680, Z => n1679);
   U289 : BUF_X1 port map( A => n1674, Z => n1673);
   U290 : BUF_X1 port map( A => n1668, Z => n1667);
   U291 : BUF_X1 port map( A => n1662, Z => n1661);
   U292 : BUF_X1 port map( A => n1656, Z => n1655);
   U293 : BUF_X1 port map( A => n1650, Z => n1649);
   U294 : BUF_X1 port map( A => n1644, Z => n1643);
   U295 : BUF_X1 port map( A => n1638, Z => n1637);
   U296 : BUF_X1 port map( A => n1632, Z => n1631);
   U297 : BUF_X1 port map( A => n1818, Z => n1816);
   U298 : BUF_X1 port map( A => n1812, Z => n1810);
   U299 : BUF_X1 port map( A => n1806, Z => n1804);
   U300 : BUF_X1 port map( A => n1800, Z => n1798);
   U301 : BUF_X1 port map( A => n1794, Z => n1792);
   U302 : BUF_X1 port map( A => n1788, Z => n1786);
   U303 : BUF_X1 port map( A => n1782, Z => n1780);
   U304 : BUF_X1 port map( A => n1776, Z => n1774);
   U305 : BUF_X1 port map( A => n1770, Z => n1768);
   U306 : BUF_X1 port map( A => n1764, Z => n1762);
   U307 : BUF_X1 port map( A => n1758, Z => n1756);
   U308 : BUF_X1 port map( A => n1752, Z => n1750);
   U309 : BUF_X1 port map( A => n1746, Z => n1744);
   U310 : BUF_X1 port map( A => n1740, Z => n1738);
   U311 : BUF_X1 port map( A => n1734, Z => n1732);
   U312 : BUF_X1 port map( A => n1728, Z => n1726);
   U313 : BUF_X1 port map( A => n1722, Z => n1720);
   U314 : BUF_X1 port map( A => n1716, Z => n1714);
   U315 : BUF_X1 port map( A => n1710, Z => n1708);
   U316 : BUF_X1 port map( A => n1704, Z => n1702);
   U317 : BUF_X1 port map( A => n1698, Z => n1696);
   U318 : BUF_X1 port map( A => n1692, Z => n1690);
   U319 : BUF_X1 port map( A => n1686, Z => n1684);
   U320 : BUF_X1 port map( A => n1680, Z => n1678);
   U321 : BUF_X1 port map( A => n1674, Z => n1672);
   U322 : BUF_X1 port map( A => n1668, Z => n1666);
   U323 : BUF_X1 port map( A => n1662, Z => n1660);
   U324 : BUF_X1 port map( A => n1656, Z => n1654);
   U325 : BUF_X1 port map( A => n1650, Z => n1648);
   U326 : BUF_X1 port map( A => n1644, Z => n1642);
   U327 : BUF_X1 port map( A => n1638, Z => n1636);
   U328 : BUF_X1 port map( A => n1632, Z => n1630);
   U329 : BUF_X1 port map( A => n862, Z => n863);
   U330 : BUF_X1 port map( A => n826, Z => n827);
   U331 : INV_X1 port map( A => ADD_RD2(0), ZN => n1592);
   U332 : INV_X1 port map( A => ADD_RD2(2), ZN => n1590);
   U333 : INV_X1 port map( A => ADD_RD2(1), ZN => n1591);
   U334 : INV_X1 port map( A => ADD_RD2(3), ZN => n1589);
   U335 : BUF_X1 port map( A => n13, Z => n875);
   U336 : BUF_X1 port map( A => n12, Z => n857);
   U337 : BUF_X1 port map( A => n11, Z => n839);
   U338 : BUF_X1 port map( A => n10, Z => n821);
   U339 : BUF_X1 port map( A => RST, Z => n1620);
   U340 : BUF_X1 port map( A => n808, Z => n811);
   U341 : BUF_X1 port map( A => n772, Z => n775);
   U342 : BUF_X1 port map( A => n808, Z => n810);
   U343 : BUF_X1 port map( A => n772, Z => n774);
   U344 : BUF_X1 port map( A => n790, Z => n793);
   U345 : BUF_X1 port map( A => n754, Z => n757);
   U346 : BUF_X1 port map( A => n790, Z => n792);
   U347 : BUF_X1 port map( A => n754, Z => n756);
   U348 : BUF_X1 port map( A => n2057, Z => n2054);
   U349 : BUF_X1 port map( A => n2057, Z => n2055);
   U350 : BUF_X1 port map( A => n2050, Z => n2047);
   U351 : BUF_X1 port map( A => n2050, Z => n2048);
   U352 : BUF_X1 port map( A => n2043, Z => n2040);
   U353 : BUF_X1 port map( A => n2043, Z => n2041);
   U354 : BUF_X1 port map( A => n2036, Z => n2033);
   U355 : BUF_X1 port map( A => n2036, Z => n2034);
   U356 : BUF_X1 port map( A => n2029, Z => n2026);
   U357 : BUF_X1 port map( A => n2029, Z => n2027);
   U358 : BUF_X1 port map( A => n2022, Z => n2019);
   U359 : BUF_X1 port map( A => n2022, Z => n2020);
   U360 : BUF_X1 port map( A => n2015, Z => n2012);
   U361 : BUF_X1 port map( A => n2015, Z => n2013);
   U362 : BUF_X1 port map( A => n2008, Z => n2005);
   U363 : BUF_X1 port map( A => n2008, Z => n2006);
   U364 : BUF_X1 port map( A => n2001, Z => n1998);
   U365 : BUF_X1 port map( A => n2001, Z => n1999);
   U366 : BUF_X1 port map( A => n1994, Z => n1991);
   U367 : BUF_X1 port map( A => n1994, Z => n1992);
   U368 : BUF_X1 port map( A => n1987, Z => n1984);
   U369 : BUF_X1 port map( A => n1987, Z => n1985);
   U370 : BUF_X1 port map( A => n1980, Z => n1977);
   U371 : BUF_X1 port map( A => n1980, Z => n1978);
   U372 : BUF_X1 port map( A => n1973, Z => n1970);
   U373 : BUF_X1 port map( A => n1973, Z => n1971);
   U374 : BUF_X1 port map( A => n1966, Z => n1963);
   U375 : BUF_X1 port map( A => n1966, Z => n1964);
   U376 : BUF_X1 port map( A => n1959, Z => n1956);
   U377 : BUF_X1 port map( A => n1959, Z => n1957);
   U378 : BUF_X1 port map( A => n1952, Z => n1949);
   U379 : BUF_X1 port map( A => n1952, Z => n1950);
   U380 : BUF_X1 port map( A => n1945, Z => n1942);
   U381 : BUF_X1 port map( A => n1945, Z => n1943);
   U382 : BUF_X1 port map( A => n1938, Z => n1935);
   U383 : BUF_X1 port map( A => n1938, Z => n1936);
   U384 : BUF_X1 port map( A => n1931, Z => n1928);
   U385 : BUF_X1 port map( A => n1931, Z => n1929);
   U386 : BUF_X1 port map( A => n1924, Z => n1921);
   U387 : BUF_X1 port map( A => n1924, Z => n1922);
   U388 : BUF_X1 port map( A => n1917, Z => n1914);
   U389 : BUF_X1 port map( A => n1917, Z => n1915);
   U390 : BUF_X1 port map( A => n1910, Z => n1907);
   U391 : BUF_X1 port map( A => n1910, Z => n1908);
   U392 : BUF_X1 port map( A => n1903, Z => n1900);
   U393 : BUF_X1 port map( A => n1903, Z => n1901);
   U394 : BUF_X1 port map( A => n1896, Z => n1893);
   U395 : BUF_X1 port map( A => n1896, Z => n1894);
   U396 : BUF_X1 port map( A => n1889, Z => n1886);
   U397 : BUF_X1 port map( A => n1889, Z => n1887);
   U398 : BUF_X1 port map( A => n1882, Z => n1879);
   U399 : BUF_X1 port map( A => n1882, Z => n1880);
   U400 : BUF_X1 port map( A => n1875, Z => n1872);
   U401 : BUF_X1 port map( A => n1875, Z => n1873);
   U402 : BUF_X1 port map( A => n1868, Z => n1865);
   U403 : BUF_X1 port map( A => n1868, Z => n1866);
   U404 : BUF_X1 port map( A => n1861, Z => n1858);
   U405 : BUF_X1 port map( A => n1861, Z => n1859);
   U406 : BUF_X1 port map( A => n1854, Z => n1851);
   U407 : BUF_X1 port map( A => n1854, Z => n1852);
   U408 : BUF_X1 port map( A => n1847, Z => n1844);
   U409 : BUF_X1 port map( A => n1847, Z => n1845);
   U410 : BUF_X1 port map( A => n1840, Z => n1837);
   U411 : BUF_X1 port map( A => n1840, Z => n1838);
   U412 : BUF_X1 port map( A => n808, Z => n809);
   U413 : BUF_X1 port map( A => n772, Z => n773);
   U414 : BUF_X1 port map( A => n790, Z => n791);
   U415 : BUF_X1 port map( A => n754, Z => n755);
   U416 : BUF_X1 port map( A => n1819, Z => n1815);
   U417 : BUF_X1 port map( A => n1820, Z => n1819);
   U418 : BUF_X1 port map( A => n1813, Z => n1809);
   U419 : BUF_X1 port map( A => n1814, Z => n1813);
   U420 : BUF_X1 port map( A => n1807, Z => n1803);
   U421 : BUF_X1 port map( A => n1808, Z => n1807);
   U422 : BUF_X1 port map( A => n1801, Z => n1797);
   U423 : BUF_X1 port map( A => n1802, Z => n1801);
   U424 : BUF_X1 port map( A => n1795, Z => n1791);
   U425 : BUF_X1 port map( A => n1796, Z => n1795);
   U426 : BUF_X1 port map( A => n1789, Z => n1785);
   U427 : BUF_X1 port map( A => n1790, Z => n1789);
   U428 : BUF_X1 port map( A => n1783, Z => n1779);
   U429 : BUF_X1 port map( A => n1784, Z => n1783);
   U430 : BUF_X1 port map( A => n1777, Z => n1773);
   U431 : BUF_X1 port map( A => n1778, Z => n1777);
   U432 : BUF_X1 port map( A => n1771, Z => n1767);
   U433 : BUF_X1 port map( A => n1772, Z => n1771);
   U434 : BUF_X1 port map( A => n1765, Z => n1761);
   U435 : BUF_X1 port map( A => n1766, Z => n1765);
   U436 : BUF_X1 port map( A => n1759, Z => n1755);
   U437 : BUF_X1 port map( A => n1760, Z => n1759);
   U438 : BUF_X1 port map( A => n1753, Z => n1749);
   U439 : BUF_X1 port map( A => n1754, Z => n1753);
   U440 : BUF_X1 port map( A => n1747, Z => n1743);
   U441 : BUF_X1 port map( A => n1748, Z => n1747);
   U442 : BUF_X1 port map( A => n1741, Z => n1737);
   U443 : BUF_X1 port map( A => n1742, Z => n1741);
   U444 : BUF_X1 port map( A => n1735, Z => n1731);
   U445 : BUF_X1 port map( A => n1736, Z => n1735);
   U446 : BUF_X1 port map( A => n1729, Z => n1725);
   U447 : BUF_X1 port map( A => n1730, Z => n1729);
   U448 : BUF_X1 port map( A => n1723, Z => n1719);
   U449 : BUF_X1 port map( A => n1724, Z => n1723);
   U450 : BUF_X1 port map( A => n1717, Z => n1713);
   U451 : BUF_X1 port map( A => n1718, Z => n1717);
   U452 : BUF_X1 port map( A => n1711, Z => n1707);
   U453 : BUF_X1 port map( A => n1712, Z => n1711);
   U454 : BUF_X1 port map( A => n1705, Z => n1701);
   U455 : BUF_X1 port map( A => n1706, Z => n1705);
   U456 : BUF_X1 port map( A => n1699, Z => n1695);
   U457 : BUF_X1 port map( A => n1700, Z => n1699);
   U458 : BUF_X1 port map( A => n1693, Z => n1689);
   U459 : BUF_X1 port map( A => n1694, Z => n1693);
   U460 : BUF_X1 port map( A => n1687, Z => n1683);
   U461 : BUF_X1 port map( A => n1688, Z => n1687);
   U462 : BUF_X1 port map( A => n1681, Z => n1677);
   U463 : BUF_X1 port map( A => n1682, Z => n1681);
   U464 : BUF_X1 port map( A => n1675, Z => n1671);
   U465 : BUF_X1 port map( A => n1676, Z => n1675);
   U466 : BUF_X1 port map( A => n1669, Z => n1665);
   U467 : BUF_X1 port map( A => n1670, Z => n1669);
   U468 : BUF_X1 port map( A => n1663, Z => n1659);
   U469 : BUF_X1 port map( A => n1664, Z => n1663);
   U470 : BUF_X1 port map( A => n1657, Z => n1653);
   U471 : BUF_X1 port map( A => n1658, Z => n1657);
   U472 : BUF_X1 port map( A => n1651, Z => n1647);
   U473 : BUF_X1 port map( A => n1652, Z => n1651);
   U474 : BUF_X1 port map( A => n1645, Z => n1641);
   U475 : BUF_X1 port map( A => n1646, Z => n1645);
   U476 : BUF_X1 port map( A => n1639, Z => n1635);
   U477 : BUF_X1 port map( A => n1640, Z => n1639);
   U478 : BUF_X1 port map( A => n1633, Z => n1629);
   U479 : BUF_X1 port map( A => n1634, Z => n1633);
   U480 : BUF_X1 port map( A => n2057, Z => n2056);
   U481 : BUF_X1 port map( A => n2050, Z => n2049);
   U482 : BUF_X1 port map( A => n2043, Z => n2042);
   U483 : BUF_X1 port map( A => n2036, Z => n2035);
   U484 : BUF_X1 port map( A => n2029, Z => n2028);
   U485 : BUF_X1 port map( A => n2022, Z => n2021);
   U486 : BUF_X1 port map( A => n2015, Z => n2014);
   U487 : BUF_X1 port map( A => n2008, Z => n2007);
   U488 : BUF_X1 port map( A => n2001, Z => n2000);
   U489 : BUF_X1 port map( A => n1994, Z => n1993);
   U490 : BUF_X1 port map( A => n1987, Z => n1986);
   U491 : BUF_X1 port map( A => n1980, Z => n1979);
   U492 : BUF_X1 port map( A => n1973, Z => n1972);
   U493 : BUF_X1 port map( A => n1966, Z => n1965);
   U494 : BUF_X1 port map( A => n1959, Z => n1958);
   U495 : BUF_X1 port map( A => n1952, Z => n1951);
   U496 : BUF_X1 port map( A => n1945, Z => n1944);
   U497 : BUF_X1 port map( A => n1938, Z => n1937);
   U498 : BUF_X1 port map( A => n1931, Z => n1930);
   U499 : BUF_X1 port map( A => n1924, Z => n1923);
   U500 : BUF_X1 port map( A => n1917, Z => n1916);
   U501 : BUF_X1 port map( A => n1910, Z => n1909);
   U502 : BUF_X1 port map( A => n1903, Z => n1902);
   U503 : BUF_X1 port map( A => n1896, Z => n1895);
   U504 : BUF_X1 port map( A => n1889, Z => n1888);
   U505 : BUF_X1 port map( A => n1882, Z => n1881);
   U506 : BUF_X1 port map( A => n1875, Z => n1874);
   U507 : BUF_X1 port map( A => n1868, Z => n1867);
   U508 : BUF_X1 port map( A => n1861, Z => n1860);
   U509 : BUF_X1 port map( A => n1854, Z => n1853);
   U510 : BUF_X1 port map( A => n1847, Z => n1846);
   U511 : BUF_X1 port map( A => n1840, Z => n1839);
   U512 : NOR2_X1 port map( A1 => n1821, A2 => n72, ZN => N219);
   U513 : NOR2_X1 port map( A1 => n1821, A2 => n71, ZN => N220);
   U514 : NOR2_X1 port map( A1 => n1821, A2 => n70, ZN => N221);
   U515 : NOR2_X1 port map( A1 => n1821, A2 => n69, ZN => N222);
   U516 : NOR2_X1 port map( A1 => n1821, A2 => n68, ZN => N223);
   U517 : NOR2_X1 port map( A1 => n1821, A2 => n67, ZN => N224);
   U518 : NOR2_X1 port map( A1 => n1821, A2 => n66, ZN => N225);
   U519 : NOR2_X1 port map( A1 => n1821, A2 => n65, ZN => N226);
   U520 : NOR2_X1 port map( A1 => n1821, A2 => n64, ZN => N227);
   U521 : NOR2_X1 port map( A1 => n1821, A2 => n63, ZN => N228);
   U522 : NOR2_X1 port map( A1 => n1821, A2 => n62, ZN => N229);
   U523 : NOR2_X1 port map( A1 => n1822, A2 => n61, ZN => N230);
   U524 : NOR2_X1 port map( A1 => n1822, A2 => n60, ZN => N231);
   U525 : NOR2_X1 port map( A1 => n1822, A2 => n59, ZN => N232);
   U526 : NOR2_X1 port map( A1 => n1822, A2 => n58, ZN => N233);
   U527 : NOR2_X1 port map( A1 => n1822, A2 => n57, ZN => N234);
   U528 : NOR2_X1 port map( A1 => n1822, A2 => n56, ZN => N235);
   U529 : NOR2_X1 port map( A1 => n1822, A2 => n55, ZN => N236);
   U530 : NOR2_X1 port map( A1 => n1822, A2 => n54, ZN => N237);
   U531 : NOR2_X1 port map( A1 => n1822, A2 => n53, ZN => N238);
   U532 : NOR2_X1 port map( A1 => n1822, A2 => n52, ZN => N239);
   U533 : NOR2_X1 port map( A1 => n1822, A2 => n51, ZN => N240);
   U534 : NOR2_X1 port map( A1 => n1821, A2 => n50, ZN => N241);
   U535 : NOR2_X1 port map( A1 => n1822, A2 => n49, ZN => N242);
   U536 : NOR2_X1 port map( A1 => n1821, A2 => n48, ZN => N243);
   U537 : NOR2_X1 port map( A1 => n1822, A2 => n47, ZN => N244);
   U538 : NOR2_X1 port map( A1 => n1821, A2 => n46, ZN => N245);
   U539 : NOR2_X1 port map( A1 => n1822, A2 => n45, ZN => N246);
   U540 : NOR2_X1 port map( A1 => n1821, A2 => n44, ZN => N247);
   U541 : NOR2_X1 port map( A1 => n1822, A2 => n43, ZN => N248);
   U542 : NOR2_X1 port map( A1 => n1821, A2 => n42, ZN => N249);
   U543 : NOR2_X1 port map( A1 => n1822, A2 => n41, ZN => N250);
   U544 : BUF_X1 port map( A => n16, Z => n803);
   U545 : BUF_X1 port map( A => n17, Z => n785);
   U546 : BUF_X1 port map( A => n18, Z => n767);
   U547 : BUF_X1 port map( A => n19, Z => n749);
   U548 : BUF_X1 port map( A => n2092, Z => n1820);
   U549 : INV_X1 port map( A => n72, ZN => n2092);
   U550 : BUF_X1 port map( A => n2091, Z => n1814);
   U551 : INV_X1 port map( A => n71, ZN => n2091);
   U552 : BUF_X1 port map( A => n2090, Z => n1808);
   U553 : INV_X1 port map( A => n70, ZN => n2090);
   U554 : BUF_X1 port map( A => n2089, Z => n1802);
   U555 : INV_X1 port map( A => n69, ZN => n2089);
   U556 : BUF_X1 port map( A => n2088, Z => n1796);
   U557 : INV_X1 port map( A => n68, ZN => n2088);
   U558 : BUF_X1 port map( A => n2087, Z => n1790);
   U559 : INV_X1 port map( A => n67, ZN => n2087);
   U560 : BUF_X1 port map( A => n2086, Z => n1784);
   U561 : INV_X1 port map( A => n66, ZN => n2086);
   U562 : BUF_X1 port map( A => n2085, Z => n1778);
   U563 : INV_X1 port map( A => n65, ZN => n2085);
   U564 : BUF_X1 port map( A => n2084, Z => n1772);
   U565 : INV_X1 port map( A => n64, ZN => n2084);
   U566 : BUF_X1 port map( A => n2083, Z => n1766);
   U567 : INV_X1 port map( A => n63, ZN => n2083);
   U568 : BUF_X1 port map( A => n2082, Z => n1760);
   U569 : INV_X1 port map( A => n62, ZN => n2082);
   U570 : BUF_X1 port map( A => n2081, Z => n1754);
   U571 : INV_X1 port map( A => n61, ZN => n2081);
   U572 : BUF_X1 port map( A => n2080, Z => n1748);
   U573 : INV_X1 port map( A => n60, ZN => n2080);
   U574 : BUF_X1 port map( A => n2079, Z => n1742);
   U575 : INV_X1 port map( A => n59, ZN => n2079);
   U576 : BUF_X1 port map( A => n2078, Z => n1736);
   U577 : INV_X1 port map( A => n58, ZN => n2078);
   U578 : BUF_X1 port map( A => n2077, Z => n1730);
   U579 : INV_X1 port map( A => n57, ZN => n2077);
   U580 : BUF_X1 port map( A => n2076, Z => n1724);
   U581 : INV_X1 port map( A => n56, ZN => n2076);
   U582 : BUF_X1 port map( A => n2075, Z => n1718);
   U583 : INV_X1 port map( A => n55, ZN => n2075);
   U584 : BUF_X1 port map( A => n2074, Z => n1712);
   U585 : INV_X1 port map( A => n54, ZN => n2074);
   U586 : BUF_X1 port map( A => n2073, Z => n1706);
   U587 : INV_X1 port map( A => n53, ZN => n2073);
   U588 : BUF_X1 port map( A => n2072, Z => n1700);
   U589 : INV_X1 port map( A => n52, ZN => n2072);
   U590 : BUF_X1 port map( A => n2071, Z => n1694);
   U591 : INV_X1 port map( A => n51, ZN => n2071);
   U592 : BUF_X1 port map( A => n2070, Z => n1688);
   U593 : INV_X1 port map( A => n50, ZN => n2070);
   U594 : BUF_X1 port map( A => n2069, Z => n1682);
   U595 : INV_X1 port map( A => n49, ZN => n2069);
   U596 : BUF_X1 port map( A => n2068, Z => n1676);
   U597 : INV_X1 port map( A => n48, ZN => n2068);
   U598 : BUF_X1 port map( A => n2067, Z => n1670);
   U599 : INV_X1 port map( A => n47, ZN => n2067);
   U600 : BUF_X1 port map( A => n2066, Z => n1664);
   U601 : INV_X1 port map( A => n46, ZN => n2066);
   U602 : BUF_X1 port map( A => n2065, Z => n1658);
   U603 : INV_X1 port map( A => n45, ZN => n2065);
   U604 : BUF_X1 port map( A => n2064, Z => n1652);
   U605 : INV_X1 port map( A => n44, ZN => n2064);
   U606 : BUF_X1 port map( A => n2063, Z => n1646);
   U607 : INV_X1 port map( A => n43, ZN => n2063);
   U608 : BUF_X1 port map( A => n2062, Z => n1640);
   U609 : INV_X1 port map( A => n42, ZN => n2062);
   U610 : BUF_X1 port map( A => n2061, Z => n1634);
   U611 : INV_X1 port map( A => n41, ZN => n2061);
   U612 : INV_X1 port map( A => n1823, ZN => n1821);
   U613 : INV_X1 port map( A => n1823, ZN => n1822);
   U614 : BUF_X1 port map( A => n897, Z => n900);
   U615 : BUF_X1 port map( A => n897, Z => n899);
   U616 : BUF_X1 port map( A => n893, Z => n896);
   U617 : BUF_X1 port map( A => n893, Z => n895);
   U618 : BUF_X1 port map( A => n905, Z => n908);
   U619 : BUF_X1 port map( A => n905, Z => n907);
   U620 : BUF_X1 port map( A => n901, Z => n904);
   U621 : BUF_X1 port map( A => n901, Z => n903);
   U622 : BUF_X1 port map( A => n897, Z => n898);
   U623 : BUF_X1 port map( A => n893, Z => n894);
   U624 : BUF_X1 port map( A => n905, Z => n906);
   U625 : BUF_X1 port map( A => n901, Z => n902);
   U626 : BUF_X1 port map( A => n1834, Z => n1832);
   U627 : BUF_X1 port map( A => n1834, Z => n1831);
   U628 : BUF_X1 port map( A => n1828, Z => n1826);
   U629 : BUF_X1 port map( A => n1828, Z => n1825);
   U630 : BUF_X1 port map( A => n2058, Z => n2053);
   U631 : BUF_X1 port map( A => n2059, Z => n2058);
   U632 : BUF_X1 port map( A => n2051, Z => n2046);
   U633 : BUF_X1 port map( A => n2052, Z => n2051);
   U634 : BUF_X1 port map( A => n2044, Z => n2039);
   U635 : BUF_X1 port map( A => n2045, Z => n2044);
   U636 : BUF_X1 port map( A => n2037, Z => n2032);
   U637 : BUF_X1 port map( A => n2038, Z => n2037);
   U638 : BUF_X1 port map( A => n2030, Z => n2025);
   U639 : BUF_X1 port map( A => n2031, Z => n2030);
   U640 : BUF_X1 port map( A => n2023, Z => n2018);
   U641 : BUF_X1 port map( A => n2024, Z => n2023);
   U642 : BUF_X1 port map( A => n2016, Z => n2011);
   U643 : BUF_X1 port map( A => n2017, Z => n2016);
   U644 : BUF_X1 port map( A => n2009, Z => n2004);
   U645 : BUF_X1 port map( A => n2010, Z => n2009);
   U646 : BUF_X1 port map( A => n2002, Z => n1997);
   U647 : BUF_X1 port map( A => n2003, Z => n2002);
   U648 : BUF_X1 port map( A => n1995, Z => n1990);
   U649 : BUF_X1 port map( A => n1996, Z => n1995);
   U650 : BUF_X1 port map( A => n1988, Z => n1983);
   U651 : BUF_X1 port map( A => n1989, Z => n1988);
   U652 : BUF_X1 port map( A => n1981, Z => n1976);
   U653 : BUF_X1 port map( A => n1982, Z => n1981);
   U654 : BUF_X1 port map( A => n1974, Z => n1969);
   U655 : BUF_X1 port map( A => n1975, Z => n1974);
   U656 : BUF_X1 port map( A => n1967, Z => n1962);
   U657 : BUF_X1 port map( A => n1968, Z => n1967);
   U658 : BUF_X1 port map( A => n1960, Z => n1955);
   U659 : BUF_X1 port map( A => n1961, Z => n1960);
   U660 : BUF_X1 port map( A => n1953, Z => n1948);
   U661 : BUF_X1 port map( A => n1954, Z => n1953);
   U662 : BUF_X1 port map( A => n1946, Z => n1941);
   U663 : BUF_X1 port map( A => n1947, Z => n1946);
   U664 : BUF_X1 port map( A => n1939, Z => n1934);
   U665 : BUF_X1 port map( A => n1940, Z => n1939);
   U666 : BUF_X1 port map( A => n1932, Z => n1927);
   U667 : BUF_X1 port map( A => n1933, Z => n1932);
   U668 : BUF_X1 port map( A => n1925, Z => n1920);
   U669 : BUF_X1 port map( A => n1926, Z => n1925);
   U670 : BUF_X1 port map( A => n1918, Z => n1913);
   U671 : BUF_X1 port map( A => n1919, Z => n1918);
   U672 : BUF_X1 port map( A => n1911, Z => n1906);
   U673 : BUF_X1 port map( A => n1912, Z => n1911);
   U674 : BUF_X1 port map( A => n1904, Z => n1899);
   U675 : BUF_X1 port map( A => n1905, Z => n1904);
   U676 : BUF_X1 port map( A => n1897, Z => n1892);
   U677 : BUF_X1 port map( A => n1898, Z => n1897);
   U678 : BUF_X1 port map( A => n1890, Z => n1885);
   U679 : BUF_X1 port map( A => n1891, Z => n1890);
   U680 : BUF_X1 port map( A => n1883, Z => n1878);
   U681 : BUF_X1 port map( A => n1884, Z => n1883);
   U682 : BUF_X1 port map( A => n1876, Z => n1871);
   U683 : BUF_X1 port map( A => n1877, Z => n1876);
   U684 : BUF_X1 port map( A => n1869, Z => n1864);
   U685 : BUF_X1 port map( A => n1870, Z => n1869);
   U686 : BUF_X1 port map( A => n1862, Z => n1857);
   U687 : BUF_X1 port map( A => n1863, Z => n1862);
   U688 : BUF_X1 port map( A => n1855, Z => n1850);
   U689 : BUF_X1 port map( A => n1856, Z => n1855);
   U690 : BUF_X1 port map( A => n1848, Z => n1843);
   U691 : BUF_X1 port map( A => n1849, Z => n1848);
   U692 : BUF_X1 port map( A => n1841, Z => n1836);
   U693 : BUF_X1 port map( A => n1842, Z => n1841);
   U694 : BUF_X1 port map( A => n1834, Z => n1833);
   U695 : BUF_X1 port map( A => n1828, Z => n1827);
   U696 : NAND2_X1 port map( A1 => n1626, A2 => DATAIN(31), ZN => n41);
   U697 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n1621, ZN => n72);
   U698 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n1621, ZN => n71);
   U699 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n1621, ZN => n70);
   U700 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n1621, ZN => n69);
   U701 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n1621, ZN => n68);
   U702 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n1621, ZN => n67);
   U703 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n1621, ZN => n66);
   U704 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n1622, ZN => n65);
   U705 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n1622, ZN => n64);
   U706 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n1622, ZN => n63);
   U707 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n1622, ZN => n62);
   U708 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n1622, ZN => n61);
   U709 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n1622, ZN => n60);
   U710 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n1622, ZN => n59);
   U711 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n1621, ZN => n58);
   U712 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n1621, ZN => n57);
   U713 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n1621, ZN => n56);
   U714 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n1621, ZN => n55);
   U715 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n1621, ZN => n54);
   U716 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n1622, ZN => n53);
   U717 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n1623, ZN => n52);
   U718 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n1623, ZN => n51);
   U719 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n1623, ZN => n50);
   U720 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n1623, ZN => n49);
   U721 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n1623, ZN => n48);
   U722 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n1623, ZN => n47);
   U723 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n1623, ZN => n46);
   U724 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n1622, ZN => n45);
   U725 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n1622, ZN => n44);
   U726 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n1622, ZN => n43);
   U727 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n1622, ZN => n42);
   U728 : INV_X1 port map( A => n73, ZN => n2060);
   U729 : INV_X1 port map( A => ADD_RD1(0), ZN => n748);
   U730 : BUF_X1 port map( A => N155, Z => n2059);
   U731 : OAI21_X1 port map( B1 => n82, B2 => n85, A => n1626, ZN => N155);
   U732 : BUF_X1 port map( A => N188, Z => n2052);
   U733 : OAI21_X1 port map( B1 => n81, B2 => n85, A => n1623, ZN => N188);
   U734 : BUF_X1 port map( A => N189, Z => n2045);
   U735 : OAI21_X1 port map( B1 => n80, B2 => n85, A => n1623, ZN => N189);
   U736 : BUF_X1 port map( A => N190, Z => n2038);
   U737 : OAI21_X1 port map( B1 => n79, B2 => n85, A => n1623, ZN => N190);
   U738 : BUF_X1 port map( A => N191, Z => n2031);
   U739 : OAI21_X1 port map( B1 => n78, B2 => n85, A => n1623, ZN => N191);
   U740 : BUF_X1 port map( A => N192, Z => n2024);
   U741 : OAI21_X1 port map( B1 => n77, B2 => n85, A => n1624, ZN => N192);
   U742 : BUF_X1 port map( A => N193, Z => n2017);
   U743 : OAI21_X1 port map( B1 => n76, B2 => n85, A => n1624, ZN => N193);
   U744 : BUF_X1 port map( A => N194, Z => n2010);
   U745 : OAI21_X1 port map( B1 => n74, B2 => n85, A => n1624, ZN => N194);
   U746 : BUF_X1 port map( A => N195, Z => n2003);
   U747 : OAI21_X1 port map( B1 => n82, B2 => n84, A => n1624, ZN => N195);
   U748 : BUF_X1 port map( A => N196, Z => n1996);
   U749 : OAI21_X1 port map( B1 => n81, B2 => n84, A => n1624, ZN => N196);
   U750 : BUF_X1 port map( A => N197, Z => n1989);
   U751 : OAI21_X1 port map( B1 => n80, B2 => n84, A => n1624, ZN => N197);
   U752 : BUF_X1 port map( A => N198, Z => n1982);
   U753 : OAI21_X1 port map( B1 => n79, B2 => n84, A => n1624, ZN => N198);
   U754 : BUF_X1 port map( A => N199, Z => n1975);
   U755 : OAI21_X1 port map( B1 => n78, B2 => n84, A => n1624, ZN => N199);
   U756 : BUF_X1 port map( A => N200, Z => n1968);
   U757 : OAI21_X1 port map( B1 => n77, B2 => n84, A => n1624, ZN => N200);
   U758 : BUF_X1 port map( A => N201, Z => n1961);
   U759 : OAI21_X1 port map( B1 => n76, B2 => n84, A => n1624, ZN => N201);
   U760 : BUF_X1 port map( A => N202, Z => n1954);
   U761 : OAI21_X1 port map( B1 => n74, B2 => n84, A => n1624, ZN => N202);
   U762 : BUF_X1 port map( A => N203, Z => n1947);
   U763 : OAI21_X1 port map( B1 => n82, B2 => n83, A => n1624, ZN => N203);
   U764 : BUF_X1 port map( A => N204, Z => n1940);
   U765 : OAI21_X1 port map( B1 => n81, B2 => n83, A => n1625, ZN => N204);
   U766 : BUF_X1 port map( A => N205, Z => n1933);
   U767 : OAI21_X1 port map( B1 => n80, B2 => n83, A => n1625, ZN => N205);
   U768 : BUF_X1 port map( A => N206, Z => n1926);
   U769 : OAI21_X1 port map( B1 => n79, B2 => n83, A => n1625, ZN => N206);
   U770 : BUF_X1 port map( A => N207, Z => n1919);
   U771 : OAI21_X1 port map( B1 => n78, B2 => n83, A => n1625, ZN => N207);
   U772 : BUF_X1 port map( A => N208, Z => n1912);
   U773 : OAI21_X1 port map( B1 => n77, B2 => n83, A => n1625, ZN => N208);
   U774 : BUF_X1 port map( A => N209, Z => n1905);
   U775 : OAI21_X1 port map( B1 => n76, B2 => n83, A => n1625, ZN => N209);
   U776 : BUF_X1 port map( A => N210, Z => n1898);
   U777 : OAI21_X1 port map( B1 => n74, B2 => n83, A => n1625, ZN => N210);
   U778 : BUF_X1 port map( A => N211, Z => n1891);
   U779 : OAI21_X1 port map( B1 => n75, B2 => n82, A => n1625, ZN => N211);
   U780 : BUF_X1 port map( A => N212, Z => n1884);
   U781 : OAI21_X1 port map( B1 => n75, B2 => n81, A => n1625, ZN => N212);
   U782 : BUF_X1 port map( A => N213, Z => n1877);
   U783 : OAI21_X1 port map( B1 => n75, B2 => n80, A => n1625, ZN => N213);
   U784 : BUF_X1 port map( A => N214, Z => n1870);
   U785 : OAI21_X1 port map( B1 => n75, B2 => n79, A => n1625, ZN => N214);
   U786 : BUF_X1 port map( A => N215, Z => n1863);
   U787 : OAI21_X1 port map( B1 => n75, B2 => n78, A => n1625, ZN => N215);
   U788 : BUF_X1 port map( A => N216, Z => n1856);
   U789 : OAI21_X1 port map( B1 => n75, B2 => n77, A => n1626, ZN => N216);
   U790 : BUF_X1 port map( A => N217, Z => n1849);
   U791 : OAI21_X1 port map( B1 => n75, B2 => n76, A => n1626, ZN => N217);
   U792 : BUF_X1 port map( A => N218, Z => n1842);
   U793 : OAI21_X1 port map( B1 => n1, B2 => n73, A => n1623, ZN => N218);
   U794 : INV_X1 port map( A => ADD_RD1(2), ZN => n746);
   U795 : INV_X1 port map( A => ADD_RD1(3), ZN => n745);
   U796 : INV_X1 port map( A => ADD_RD1(1), ZN => n747);
   U797 : BUF_X1 port map( A => n1835, Z => n1830);
   U798 : BUF_X1 port map( A => n14, Z => n1835);
   U799 : BUF_X1 port map( A => n1829, Z => n1824);
   U800 : BUF_X1 port map( A => n15, Z => n1829);
   U801 : INV_X1 port map( A => ADD_WR(2), ZN => n2095);
   U802 : INV_X1 port map( A => ADD_WR(1), ZN => n2096);
   U803 : INV_X1 port map( A => ADD_WR(0), ZN => n2097);
   U804 : NAND2_X1 port map( A1 => EN_WR, A2 => EN, ZN => n73);
   U805 : INV_X1 port map( A => ADD_WR(4), ZN => n2093);
   U806 : INV_X1 port map( A => ADD_WR(3), ZN => n2094);
   U807 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n745, ZN => n743);
   U808 : NOR2_X1 port map( A1 => n746, A2 => ADD_RD1(1), ZN => n20);
   U809 : NOR2_X1 port map( A1 => n746, A2 => n747, ZN => n21);
   U810 : AOI22_X1 port map( A1 => REG_21_0_port, A2 => n784, B1 => 
                           REG_23_0_port, B2 => n766, ZN => n27);
   U811 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n22);
   U812 : NOR2_X1 port map( A1 => n747, A2 => ADD_RD1(2), ZN => n23);
   U813 : AOI22_X1 port map( A1 => REG_17_0_port, A2 => n820, B1 => 
                           REG_19_0_port, B2 => n802, ZN => n26);
   U814 : AOI22_X1 port map( A1 => REG_20_0_port, A2 => n856, B1 => 
                           REG_22_0_port, B2 => n838, ZN => n25);
   U815 : AOI22_X1 port map( A1 => REG_16_0_port, A2 => n892, B1 => 
                           REG_18_0_port, B2 => n874, ZN => n24);
   U816 : AND4_X1 port map( A1 => n27, A2 => n26, A3 => n25, A4 => n24, ZN => 
                           n89);
   U817 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n741);
   U818 : AOI22_X1 port map( A1 => REG_29_0_port, A2 => n784, B1 => 
                           REG_31_0_port, B2 => n766, ZN => n31);
   U819 : AOI22_X1 port map( A1 => REG_25_0_port, A2 => n820, B1 => 
                           REG_27_0_port, B2 => n802, ZN => n30);
   U820 : AOI22_X1 port map( A1 => REG_28_0_port, A2 => n856, B1 => 
                           REG_30_0_port, B2 => n838, ZN => n29);
   U821 : AOI22_X1 port map( A1 => REG_24_0_port, A2 => n892, B1 => 
                           REG_26_0_port, B2 => n874, ZN => n28);
   U822 : AND4_X1 port map( A1 => n31, A2 => n30, A3 => n29, A4 => n28, ZN => 
                           n88);
   U823 : AOI22_X1 port map( A1 => REG_5_0_port, A2 => n784, B1 => REG_7_0_port
                           , B2 => n766, ZN => n35);
   U824 : AOI22_X1 port map( A1 => REG_1_0_port, A2 => n820, B1 => REG_3_0_port
                           , B2 => n802, ZN => n34);
   U825 : AOI22_X1 port map( A1 => REG_4_0_port, A2 => n856, B1 => REG_6_0_port
                           , B2 => n838, ZN => n33);
   U826 : AOI22_X1 port map( A1 => REG_0_0_port, A2 => n892, B1 => REG_2_0_port
                           , B2 => n874, ZN => n32);
   U827 : NAND4_X1 port map( A1 => n35, A2 => n34, A3 => n33, A4 => n32, ZN => 
                           n86);
   U828 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n739);
   U829 : AOI22_X1 port map( A1 => REG_13_0_port, A2 => n784, B1 => 
                           REG_15_0_port, B2 => n766, ZN => n39);
   U830 : AOI22_X1 port map( A1 => REG_9_0_port, A2 => n820, B1 => 
                           REG_11_0_port, B2 => n802, ZN => n38);
   U831 : AOI22_X1 port map( A1 => REG_12_0_port, A2 => n856, B1 => 
                           REG_14_0_port, B2 => n838, ZN => n37);
   U832 : AOI22_X1 port map( A1 => REG_8_0_port, A2 => n892, B1 => 
                           REG_10_0_port, B2 => n874, ZN => n36);
   U833 : NAND4_X1 port map( A1 => n39, A2 => n38, A3 => n37, A4 => n36, ZN => 
                           n40);
   U834 : NOR2_X1 port map( A1 => n745, A2 => ADD_RD1(4), ZN => n737);
   U835 : AOI22_X1 port map( A1 => n86, A2 => n900, B1 => n40, B2 => n896, ZN 
                           => n87);
   U836 : OAI221_X1 port map( B1 => n908, B2 => n89, C1 => n902, C2 => n88, A 
                           => n87, ZN => N283);
   U837 : AOI22_X1 port map( A1 => REG_21_1_port, A2 => n784, B1 => 
                           REG_23_1_port, B2 => n766, ZN => n93);
   U838 : AOI22_X1 port map( A1 => REG_17_1_port, A2 => n820, B1 => 
                           REG_19_1_port, B2 => n802, ZN => n92);
   U839 : AOI22_X1 port map( A1 => REG_20_1_port, A2 => n856, B1 => 
                           REG_22_1_port, B2 => n838, ZN => n91);
   U840 : AOI22_X1 port map( A1 => REG_16_1_port, A2 => n892, B1 => 
                           REG_18_1_port, B2 => n874, ZN => n90);
   U841 : AND4_X1 port map( A1 => n93, A2 => n92, A3 => n91, A4 => n90, ZN => 
                           n110);
   U842 : AOI22_X1 port map( A1 => REG_29_1_port, A2 => n784, B1 => 
                           REG_31_1_port, B2 => n766, ZN => n97);
   U843 : AOI22_X1 port map( A1 => REG_25_1_port, A2 => n820, B1 => 
                           REG_27_1_port, B2 => n802, ZN => n96);
   U844 : AOI22_X1 port map( A1 => REG_28_1_port, A2 => n856, B1 => 
                           REG_30_1_port, B2 => n838, ZN => n95);
   U845 : AOI22_X1 port map( A1 => REG_24_1_port, A2 => n892, B1 => 
                           REG_26_1_port, B2 => n874, ZN => n94);
   U846 : AND4_X1 port map( A1 => n97, A2 => n96, A3 => n95, A4 => n94, ZN => 
                           n109);
   U847 : AOI22_X1 port map( A1 => REG_5_1_port, A2 => n784, B1 => REG_7_1_port
                           , B2 => n766, ZN => n101);
   U848 : AOI22_X1 port map( A1 => REG_1_1_port, A2 => n820, B1 => REG_3_1_port
                           , B2 => n802, ZN => n100);
   U849 : AOI22_X1 port map( A1 => REG_4_1_port, A2 => n856, B1 => REG_6_1_port
                           , B2 => n838, ZN => n99);
   U850 : AOI22_X1 port map( A1 => REG_0_1_port, A2 => n892, B1 => REG_2_1_port
                           , B2 => n874, ZN => n98);
   U851 : NAND4_X1 port map( A1 => n101, A2 => n100, A3 => n99, A4 => n98, ZN 
                           => n107);
   U852 : AOI22_X1 port map( A1 => REG_13_1_port, A2 => n784, B1 => 
                           REG_15_1_port, B2 => n766, ZN => n105);
   U853 : AOI22_X1 port map( A1 => REG_9_1_port, A2 => n820, B1 => 
                           REG_11_1_port, B2 => n802, ZN => n104);
   U854 : AOI22_X1 port map( A1 => REG_12_1_port, A2 => n856, B1 => 
                           REG_14_1_port, B2 => n838, ZN => n103);
   U855 : AOI22_X1 port map( A1 => REG_8_1_port, A2 => n892, B1 => 
                           REG_10_1_port, B2 => n874, ZN => n102);
   U856 : NAND4_X1 port map( A1 => n105, A2 => n104, A3 => n103, A4 => n102, ZN
                           => n106);
   U857 : AOI22_X1 port map( A1 => n107, A2 => n900, B1 => n106, B2 => n896, ZN
                           => n108);
   U858 : OAI221_X1 port map( B1 => n908, B2 => n110, C1 => n902, C2 => n109, A
                           => n108, ZN => N282);
   U859 : AOI22_X1 port map( A1 => REG_21_2_port, A2 => n784, B1 => 
                           REG_23_2_port, B2 => n766, ZN => n114);
   U860 : AOI22_X1 port map( A1 => REG_17_2_port, A2 => n820, B1 => 
                           REG_19_2_port, B2 => n802, ZN => n113);
   U861 : AOI22_X1 port map( A1 => REG_20_2_port, A2 => n856, B1 => 
                           REG_22_2_port, B2 => n838, ZN => n112);
   U862 : AOI22_X1 port map( A1 => REG_16_2_port, A2 => n892, B1 => 
                           REG_18_2_port, B2 => n874, ZN => n111);
   U863 : AND4_X1 port map( A1 => n114, A2 => n113, A3 => n112, A4 => n111, ZN 
                           => n131);
   U864 : AOI22_X1 port map( A1 => REG_29_2_port, A2 => n784, B1 => 
                           REG_31_2_port, B2 => n766, ZN => n118);
   U865 : AOI22_X1 port map( A1 => REG_25_2_port, A2 => n820, B1 => 
                           REG_27_2_port, B2 => n802, ZN => n117);
   U866 : AOI22_X1 port map( A1 => REG_28_2_port, A2 => n856, B1 => 
                           REG_30_2_port, B2 => n838, ZN => n116);
   U867 : AOI22_X1 port map( A1 => REG_24_2_port, A2 => n892, B1 => 
                           REG_26_2_port, B2 => n874, ZN => n115);
   U868 : AND4_X1 port map( A1 => n118, A2 => n117, A3 => n116, A4 => n115, ZN 
                           => n130);
   U869 : AOI22_X1 port map( A1 => REG_5_2_port, A2 => n784, B1 => REG_7_2_port
                           , B2 => n766, ZN => n122);
   U870 : AOI22_X1 port map( A1 => REG_1_2_port, A2 => n820, B1 => REG_3_2_port
                           , B2 => n802, ZN => n121);
   U871 : AOI22_X1 port map( A1 => REG_4_2_port, A2 => n856, B1 => REG_6_2_port
                           , B2 => n838, ZN => n120);
   U872 : AOI22_X1 port map( A1 => REG_0_2_port, A2 => n892, B1 => REG_2_2_port
                           , B2 => n874, ZN => n119);
   U873 : NAND4_X1 port map( A1 => n122, A2 => n121, A3 => n120, A4 => n119, ZN
                           => n128);
   U874 : AOI22_X1 port map( A1 => REG_13_2_port, A2 => n783, B1 => 
                           REG_15_2_port, B2 => n765, ZN => n126);
   U875 : AOI22_X1 port map( A1 => REG_9_2_port, A2 => n819, B1 => 
                           REG_11_2_port, B2 => n801, ZN => n125);
   U876 : AOI22_X1 port map( A1 => REG_12_2_port, A2 => n855, B1 => 
                           REG_14_2_port, B2 => n837, ZN => n124);
   U877 : AOI22_X1 port map( A1 => REG_8_2_port, A2 => n891, B1 => 
                           REG_10_2_port, B2 => n873, ZN => n123);
   U878 : NAND4_X1 port map( A1 => n126, A2 => n125, A3 => n124, A4 => n123, ZN
                           => n127);
   U879 : AOI22_X1 port map( A1 => n128, A2 => n900, B1 => n127, B2 => n896, ZN
                           => n129);
   U880 : OAI221_X1 port map( B1 => n908, B2 => n131, C1 => n902, C2 => n130, A
                           => n129, ZN => N281);
   U881 : AOI22_X1 port map( A1 => REG_21_3_port, A2 => n783, B1 => 
                           REG_23_3_port, B2 => n765, ZN => n135);
   U882 : AOI22_X1 port map( A1 => REG_17_3_port, A2 => n819, B1 => 
                           REG_19_3_port, B2 => n801, ZN => n134);
   U883 : AOI22_X1 port map( A1 => REG_20_3_port, A2 => n855, B1 => 
                           REG_22_3_port, B2 => n837, ZN => n133);
   U884 : AOI22_X1 port map( A1 => REG_16_3_port, A2 => n891, B1 => 
                           REG_18_3_port, B2 => n873, ZN => n132);
   U885 : AND4_X1 port map( A1 => n135, A2 => n134, A3 => n133, A4 => n132, ZN 
                           => n152);
   U886 : AOI22_X1 port map( A1 => REG_29_3_port, A2 => n783, B1 => 
                           REG_31_3_port, B2 => n765, ZN => n139);
   U887 : AOI22_X1 port map( A1 => REG_25_3_port, A2 => n819, B1 => 
                           REG_27_3_port, B2 => n801, ZN => n138);
   U888 : AOI22_X1 port map( A1 => REG_28_3_port, A2 => n855, B1 => 
                           REG_30_3_port, B2 => n837, ZN => n137);
   U889 : AOI22_X1 port map( A1 => REG_24_3_port, A2 => n891, B1 => 
                           REG_26_3_port, B2 => n873, ZN => n136);
   U890 : AND4_X1 port map( A1 => n139, A2 => n138, A3 => n137, A4 => n136, ZN 
                           => n151);
   U891 : AOI22_X1 port map( A1 => REG_5_3_port, A2 => n783, B1 => REG_7_3_port
                           , B2 => n765, ZN => n143);
   U892 : AOI22_X1 port map( A1 => REG_1_3_port, A2 => n819, B1 => REG_3_3_port
                           , B2 => n801, ZN => n142);
   U893 : AOI22_X1 port map( A1 => REG_4_3_port, A2 => n855, B1 => REG_6_3_port
                           , B2 => n837, ZN => n141);
   U894 : AOI22_X1 port map( A1 => REG_0_3_port, A2 => n891, B1 => REG_2_3_port
                           , B2 => n873, ZN => n140);
   U895 : NAND4_X1 port map( A1 => n143, A2 => n142, A3 => n141, A4 => n140, ZN
                           => n149);
   U896 : AOI22_X1 port map( A1 => REG_13_3_port, A2 => n783, B1 => 
                           REG_15_3_port, B2 => n765, ZN => n147);
   U897 : AOI22_X1 port map( A1 => REG_9_3_port, A2 => n819, B1 => 
                           REG_11_3_port, B2 => n801, ZN => n146);
   U898 : AOI22_X1 port map( A1 => REG_12_3_port, A2 => n855, B1 => 
                           REG_14_3_port, B2 => n837, ZN => n145);
   U899 : AOI22_X1 port map( A1 => REG_8_3_port, A2 => n891, B1 => 
                           REG_10_3_port, B2 => n873, ZN => n144);
   U900 : NAND4_X1 port map( A1 => n147, A2 => n146, A3 => n145, A4 => n144, ZN
                           => n148);
   U901 : AOI22_X1 port map( A1 => n149, A2 => n900, B1 => n148, B2 => n896, ZN
                           => n150);
   U902 : OAI221_X1 port map( B1 => n908, B2 => n152, C1 => n902, C2 => n151, A
                           => n150, ZN => N280);
   U903 : AOI22_X1 port map( A1 => REG_21_4_port, A2 => n783, B1 => 
                           REG_23_4_port, B2 => n765, ZN => n156);
   U904 : AOI22_X1 port map( A1 => REG_17_4_port, A2 => n819, B1 => 
                           REG_19_4_port, B2 => n801, ZN => n155_port);
   U905 : AOI22_X1 port map( A1 => REG_20_4_port, A2 => n855, B1 => 
                           REG_22_4_port, B2 => n837, ZN => n154);
   U906 : AOI22_X1 port map( A1 => REG_16_4_port, A2 => n891, B1 => 
                           REG_18_4_port, B2 => n873, ZN => n153);
   U907 : AND4_X1 port map( A1 => n156, A2 => n155_port, A3 => n154, A4 => n153
                           , ZN => n173);
   U908 : AOI22_X1 port map( A1 => REG_29_4_port, A2 => n783, B1 => 
                           REG_31_4_port, B2 => n765, ZN => n160);
   U909 : AOI22_X1 port map( A1 => REG_25_4_port, A2 => n819, B1 => 
                           REG_27_4_port, B2 => n801, ZN => n159);
   U910 : AOI22_X1 port map( A1 => REG_28_4_port, A2 => n855, B1 => 
                           REG_30_4_port, B2 => n837, ZN => n158);
   U911 : AOI22_X1 port map( A1 => REG_24_4_port, A2 => n891, B1 => 
                           REG_26_4_port, B2 => n873, ZN => n157);
   U912 : AND4_X1 port map( A1 => n160, A2 => n159, A3 => n158, A4 => n157, ZN 
                           => n172);
   U913 : AOI22_X1 port map( A1 => REG_5_4_port, A2 => n783, B1 => REG_7_4_port
                           , B2 => n765, ZN => n164);
   U914 : AOI22_X1 port map( A1 => REG_1_4_port, A2 => n819, B1 => REG_3_4_port
                           , B2 => n801, ZN => n163);
   U915 : AOI22_X1 port map( A1 => REG_4_4_port, A2 => n855, B1 => REG_6_4_port
                           , B2 => n837, ZN => n162);
   U916 : AOI22_X1 port map( A1 => REG_0_4_port, A2 => n891, B1 => REG_2_4_port
                           , B2 => n873, ZN => n161);
   U917 : NAND4_X1 port map( A1 => n164, A2 => n163, A3 => n162, A4 => n161, ZN
                           => n170);
   U918 : AOI22_X1 port map( A1 => REG_13_4_port, A2 => n783, B1 => 
                           REG_15_4_port, B2 => n765, ZN => n168);
   U919 : AOI22_X1 port map( A1 => REG_9_4_port, A2 => n819, B1 => 
                           REG_11_4_port, B2 => n801, ZN => n167);
   U920 : AOI22_X1 port map( A1 => REG_12_4_port, A2 => n855, B1 => 
                           REG_14_4_port, B2 => n837, ZN => n166);
   U921 : AOI22_X1 port map( A1 => REG_8_4_port, A2 => n891, B1 => 
                           REG_10_4_port, B2 => n873, ZN => n165);
   U922 : NAND4_X1 port map( A1 => n168, A2 => n167, A3 => n166, A4 => n165, ZN
                           => n169);
   U923 : AOI22_X1 port map( A1 => n170, A2 => n900, B1 => n169, B2 => n896, ZN
                           => n171);
   U924 : OAI221_X1 port map( B1 => n908, B2 => n173, C1 => n902, C2 => n172, A
                           => n171, ZN => N279);
   U925 : AOI22_X1 port map( A1 => REG_21_5_port, A2 => n783, B1 => 
                           REG_23_5_port, B2 => n765, ZN => n177);
   U926 : AOI22_X1 port map( A1 => REG_17_5_port, A2 => n819, B1 => 
                           REG_19_5_port, B2 => n801, ZN => n176);
   U927 : AOI22_X1 port map( A1 => REG_20_5_port, A2 => n855, B1 => 
                           REG_22_5_port, B2 => n837, ZN => n175);
   U928 : AOI22_X1 port map( A1 => REG_16_5_port, A2 => n891, B1 => 
                           REG_18_5_port, B2 => n873, ZN => n174);
   U929 : AND4_X1 port map( A1 => n177, A2 => n176, A3 => n175, A4 => n174, ZN 
                           => n194_port);
   U930 : AOI22_X1 port map( A1 => REG_29_5_port, A2 => n783, B1 => 
                           REG_31_5_port, B2 => n765, ZN => n181);
   U931 : AOI22_X1 port map( A1 => REG_25_5_port, A2 => n819, B1 => 
                           REG_27_5_port, B2 => n801, ZN => n180);
   U932 : AOI22_X1 port map( A1 => REG_28_5_port, A2 => n855, B1 => 
                           REG_30_5_port, B2 => n837, ZN => n179);
   U933 : AOI22_X1 port map( A1 => REG_24_5_port, A2 => n891, B1 => 
                           REG_26_5_port, B2 => n873, ZN => n178);
   U934 : AND4_X1 port map( A1 => n181, A2 => n180, A3 => n179, A4 => n178, ZN 
                           => n193_port);
   U935 : AOI22_X1 port map( A1 => REG_5_5_port, A2 => n782, B1 => REG_7_5_port
                           , B2 => n764, ZN => n185);
   U936 : AOI22_X1 port map( A1 => REG_1_5_port, A2 => n818, B1 => REG_3_5_port
                           , B2 => n800, ZN => n184);
   U937 : AOI22_X1 port map( A1 => REG_4_5_port, A2 => n854, B1 => REG_6_5_port
                           , B2 => n836, ZN => n183);
   U938 : AOI22_X1 port map( A1 => REG_0_5_port, A2 => n890, B1 => REG_2_5_port
                           , B2 => n872, ZN => n182);
   U939 : NAND4_X1 port map( A1 => n185, A2 => n184, A3 => n183, A4 => n182, ZN
                           => n191_port);
   U940 : AOI22_X1 port map( A1 => REG_13_5_port, A2 => n782, B1 => 
                           REG_15_5_port, B2 => n764, ZN => n189_port);
   U941 : AOI22_X1 port map( A1 => REG_9_5_port, A2 => n818, B1 => 
                           REG_11_5_port, B2 => n800, ZN => n188_port);
   U942 : AOI22_X1 port map( A1 => REG_12_5_port, A2 => n854, B1 => 
                           REG_14_5_port, B2 => n836, ZN => n187);
   U943 : AOI22_X1 port map( A1 => REG_8_5_port, A2 => n890, B1 => 
                           REG_10_5_port, B2 => n872, ZN => n186);
   U944 : NAND4_X1 port map( A1 => n189_port, A2 => n188_port, A3 => n187, A4 
                           => n186, ZN => n190_port);
   U945 : AOI22_X1 port map( A1 => n191_port, A2 => n900, B1 => n190_port, B2 
                           => n896, ZN => n192_port);
   U946 : OAI221_X1 port map( B1 => n908, B2 => n194_port, C1 => n902, C2 => 
                           n193_port, A => n192_port, ZN => N278);
   U947 : AOI22_X1 port map( A1 => REG_21_6_port, A2 => n782, B1 => 
                           REG_23_6_port, B2 => n764, ZN => n198_port);
   U948 : AOI22_X1 port map( A1 => REG_17_6_port, A2 => n818, B1 => 
                           REG_19_6_port, B2 => n800, ZN => n197_port);
   U949 : AOI22_X1 port map( A1 => REG_20_6_port, A2 => n854, B1 => 
                           REG_22_6_port, B2 => n836, ZN => n196_port);
   U950 : AOI22_X1 port map( A1 => REG_16_6_port, A2 => n890, B1 => 
                           REG_18_6_port, B2 => n872, ZN => n195_port);
   U951 : AND4_X1 port map( A1 => n198_port, A2 => n197_port, A3 => n196_port, 
                           A4 => n195_port, ZN => n215_port);
   U952 : AOI22_X1 port map( A1 => REG_29_6_port, A2 => n782, B1 => 
                           REG_31_6_port, B2 => n764, ZN => n202_port);
   U953 : AOI22_X1 port map( A1 => REG_25_6_port, A2 => n818, B1 => 
                           REG_27_6_port, B2 => n800, ZN => n201_port);
   U954 : AOI22_X1 port map( A1 => REG_28_6_port, A2 => n854, B1 => 
                           REG_30_6_port, B2 => n836, ZN => n200_port);
   U955 : AOI22_X1 port map( A1 => REG_24_6_port, A2 => n890, B1 => 
                           REG_26_6_port, B2 => n872, ZN => n199_port);
   U956 : AND4_X1 port map( A1 => n202_port, A2 => n201_port, A3 => n200_port, 
                           A4 => n199_port, ZN => n214_port);
   U957 : AOI22_X1 port map( A1 => REG_5_6_port, A2 => n782, B1 => REG_7_6_port
                           , B2 => n764, ZN => n206_port);
   U958 : AOI22_X1 port map( A1 => REG_1_6_port, A2 => n818, B1 => REG_3_6_port
                           , B2 => n800, ZN => n205_port);
   U959 : AOI22_X1 port map( A1 => REG_4_6_port, A2 => n854, B1 => REG_6_6_port
                           , B2 => n836, ZN => n204_port);
   U960 : AOI22_X1 port map( A1 => REG_0_6_port, A2 => n890, B1 => REG_2_6_port
                           , B2 => n872, ZN => n203_port);
   U961 : NAND4_X1 port map( A1 => n206_port, A2 => n205_port, A3 => n204_port,
                           A4 => n203_port, ZN => n212_port);
   U962 : AOI22_X1 port map( A1 => REG_13_6_port, A2 => n782, B1 => 
                           REG_15_6_port, B2 => n764, ZN => n210_port);
   U963 : AOI22_X1 port map( A1 => REG_9_6_port, A2 => n818, B1 => 
                           REG_11_6_port, B2 => n800, ZN => n209_port);
   U964 : AOI22_X1 port map( A1 => REG_12_6_port, A2 => n854, B1 => 
                           REG_14_6_port, B2 => n836, ZN => n208_port);
   U965 : AOI22_X1 port map( A1 => REG_8_6_port, A2 => n890, B1 => 
                           REG_10_6_port, B2 => n872, ZN => n207_port);
   U966 : NAND4_X1 port map( A1 => n210_port, A2 => n209_port, A3 => n208_port,
                           A4 => n207_port, ZN => n211_port);
   U967 : AOI22_X1 port map( A1 => n212_port, A2 => n900, B1 => n211_port, B2 
                           => n896, ZN => n213_port);
   U968 : OAI221_X1 port map( B1 => n908, B2 => n215_port, C1 => n902, C2 => 
                           n214_port, A => n213_port, ZN => N277);
   U969 : AOI22_X1 port map( A1 => REG_21_7_port, A2 => n782, B1 => 
                           REG_23_7_port, B2 => n764, ZN => n219_port);
   U970 : AOI22_X1 port map( A1 => REG_17_7_port, A2 => n818, B1 => 
                           REG_19_7_port, B2 => n800, ZN => n218_port);
   U971 : AOI22_X1 port map( A1 => REG_20_7_port, A2 => n854, B1 => 
                           REG_22_7_port, B2 => n836, ZN => n217_port);
   U972 : AOI22_X1 port map( A1 => REG_16_7_port, A2 => n890, B1 => 
                           REG_18_7_port, B2 => n872, ZN => n216_port);
   U973 : AND4_X1 port map( A1 => n219_port, A2 => n218_port, A3 => n217_port, 
                           A4 => n216_port, ZN => n236_port);
   U974 : AOI22_X1 port map( A1 => REG_29_7_port, A2 => n782, B1 => 
                           REG_31_7_port, B2 => n764, ZN => n223_port);
   U975 : AOI22_X1 port map( A1 => REG_25_7_port, A2 => n818, B1 => 
                           REG_27_7_port, B2 => n800, ZN => n222_port);
   U976 : AOI22_X1 port map( A1 => REG_28_7_port, A2 => n854, B1 => 
                           REG_30_7_port, B2 => n836, ZN => n221_port);
   U977 : AOI22_X1 port map( A1 => REG_24_7_port, A2 => n890, B1 => 
                           REG_26_7_port, B2 => n872, ZN => n220_port);
   U978 : AND4_X1 port map( A1 => n223_port, A2 => n222_port, A3 => n221_port, 
                           A4 => n220_port, ZN => n235_port);
   U979 : AOI22_X1 port map( A1 => REG_5_7_port, A2 => n782, B1 => REG_7_7_port
                           , B2 => n764, ZN => n227_port);
   U980 : AOI22_X1 port map( A1 => REG_1_7_port, A2 => n818, B1 => REG_3_7_port
                           , B2 => n800, ZN => n226_port);
   U981 : AOI22_X1 port map( A1 => REG_4_7_port, A2 => n854, B1 => REG_6_7_port
                           , B2 => n836, ZN => n225_port);
   U982 : AOI22_X1 port map( A1 => REG_0_7_port, A2 => n890, B1 => REG_2_7_port
                           , B2 => n872, ZN => n224_port);
   U983 : NAND4_X1 port map( A1 => n227_port, A2 => n226_port, A3 => n225_port,
                           A4 => n224_port, ZN => n233_port);
   U984 : AOI22_X1 port map( A1 => REG_13_7_port, A2 => n782, B1 => 
                           REG_15_7_port, B2 => n764, ZN => n231_port);
   U985 : AOI22_X1 port map( A1 => REG_9_7_port, A2 => n818, B1 => 
                           REG_11_7_port, B2 => n800, ZN => n230_port);
   U986 : AOI22_X1 port map( A1 => REG_12_7_port, A2 => n854, B1 => 
                           REG_14_7_port, B2 => n836, ZN => n229_port);
   U987 : AOI22_X1 port map( A1 => REG_8_7_port, A2 => n890, B1 => 
                           REG_10_7_port, B2 => n872, ZN => n228_port);
   U988 : NAND4_X1 port map( A1 => n231_port, A2 => n230_port, A3 => n229_port,
                           A4 => n228_port, ZN => n232_port);
   U989 : AOI22_X1 port map( A1 => n233_port, A2 => n900, B1 => n232_port, B2 
                           => n896, ZN => n234_port);
   U990 : OAI221_X1 port map( B1 => n908, B2 => n236_port, C1 => n902, C2 => 
                           n235_port, A => n234_port, ZN => N276);
   U991 : AOI22_X1 port map( A1 => REG_21_8_port, A2 => n782, B1 => 
                           REG_23_8_port, B2 => n764, ZN => n240_port);
   U992 : AOI22_X1 port map( A1 => REG_17_8_port, A2 => n818, B1 => 
                           REG_19_8_port, B2 => n800, ZN => n239_port);
   U993 : AOI22_X1 port map( A1 => REG_20_8_port, A2 => n854, B1 => 
                           REG_22_8_port, B2 => n836, ZN => n238_port);
   U994 : AOI22_X1 port map( A1 => REG_16_8_port, A2 => n890, B1 => 
                           REG_18_8_port, B2 => n872, ZN => n237_port);
   U995 : AND4_X1 port map( A1 => n240_port, A2 => n239_port, A3 => n238_port, 
                           A4 => n237_port, ZN => n257_port);
   U996 : AOI22_X1 port map( A1 => REG_29_8_port, A2 => n781, B1 => 
                           REG_31_8_port, B2 => n763, ZN => n244_port);
   U997 : AOI22_X1 port map( A1 => REG_25_8_port, A2 => n817, B1 => 
                           REG_27_8_port, B2 => n799, ZN => n243_port);
   U998 : AOI22_X1 port map( A1 => REG_28_8_port, A2 => n853, B1 => 
                           REG_30_8_port, B2 => n835, ZN => n242_port);
   U999 : AOI22_X1 port map( A1 => REG_24_8_port, A2 => n889, B1 => 
                           REG_26_8_port, B2 => n871, ZN => n241_port);
   U1000 : AND4_X1 port map( A1 => n244_port, A2 => n243_port, A3 => n242_port,
                           A4 => n241_port, ZN => n256_port);
   U1001 : AOI22_X1 port map( A1 => REG_5_8_port, A2 => n781, B1 => 
                           REG_7_8_port, B2 => n763, ZN => n248_port);
   U1002 : AOI22_X1 port map( A1 => REG_1_8_port, A2 => n817, B1 => 
                           REG_3_8_port, B2 => n799, ZN => n247_port);
   U1003 : AOI22_X1 port map( A1 => REG_4_8_port, A2 => n853, B1 => 
                           REG_6_8_port, B2 => n835, ZN => n246_port);
   U1004 : AOI22_X1 port map( A1 => REG_0_8_port, A2 => n889, B1 => 
                           REG_2_8_port, B2 => n871, ZN => n245_port);
   U1005 : NAND4_X1 port map( A1 => n248_port, A2 => n247_port, A3 => n246_port
                           , A4 => n245_port, ZN => n254_port);
   U1006 : AOI22_X1 port map( A1 => REG_13_8_port, A2 => n781, B1 => 
                           REG_15_8_port, B2 => n763, ZN => n252_port);
   U1007 : AOI22_X1 port map( A1 => REG_9_8_port, A2 => n817, B1 => 
                           REG_11_8_port, B2 => n799, ZN => n251);
   U1008 : AOI22_X1 port map( A1 => REG_12_8_port, A2 => n853, B1 => 
                           REG_14_8_port, B2 => n835, ZN => n250_port);
   U1009 : AOI22_X1 port map( A1 => REG_8_8_port, A2 => n889, B1 => 
                           REG_10_8_port, B2 => n871, ZN => n249_port);
   U1010 : NAND4_X1 port map( A1 => n252_port, A2 => n251, A3 => n250_port, A4 
                           => n249_port, ZN => n253_port);
   U1011 : AOI22_X1 port map( A1 => n254_port, A2 => n900, B1 => n253_port, B2 
                           => n896, ZN => n255_port);
   U1012 : OAI221_X1 port map( B1 => n908, B2 => n257_port, C1 => n902, C2 => 
                           n256_port, A => n255_port, ZN => N275);
   U1013 : AOI22_X1 port map( A1 => REG_21_9_port, A2 => n781, B1 => 
                           REG_23_9_port, B2 => n763, ZN => n261_port);
   U1014 : AOI22_X1 port map( A1 => REG_17_9_port, A2 => n817, B1 => 
                           REG_19_9_port, B2 => n799, ZN => n260_port);
   U1015 : AOI22_X1 port map( A1 => REG_20_9_port, A2 => n853, B1 => 
                           REG_22_9_port, B2 => n835, ZN => n259_port);
   U1016 : AOI22_X1 port map( A1 => REG_16_9_port, A2 => n889, B1 => 
                           REG_18_9_port, B2 => n871, ZN => n258_port);
   U1017 : AND4_X1 port map( A1 => n261_port, A2 => n260_port, A3 => n259_port,
                           A4 => n258_port, ZN => n278_port);
   U1018 : AOI22_X1 port map( A1 => REG_29_9_port, A2 => n781, B1 => 
                           REG_31_9_port, B2 => n763, ZN => n265_port);
   U1019 : AOI22_X1 port map( A1 => REG_25_9_port, A2 => n817, B1 => 
                           REG_27_9_port, B2 => n799, ZN => n264_port);
   U1020 : AOI22_X1 port map( A1 => REG_28_9_port, A2 => n853, B1 => 
                           REG_30_9_port, B2 => n835, ZN => n263_port);
   U1021 : AOI22_X1 port map( A1 => REG_24_9_port, A2 => n889, B1 => 
                           REG_26_9_port, B2 => n871, ZN => n262_port);
   U1022 : AND4_X1 port map( A1 => n265_port, A2 => n264_port, A3 => n263_port,
                           A4 => n262_port, ZN => n277_port);
   U1023 : AOI22_X1 port map( A1 => REG_5_9_port, A2 => n781, B1 => 
                           REG_7_9_port, B2 => n763, ZN => n269_port);
   U1024 : AOI22_X1 port map( A1 => REG_1_9_port, A2 => n817, B1 => 
                           REG_3_9_port, B2 => n799, ZN => n268_port);
   U1025 : AOI22_X1 port map( A1 => REG_4_9_port, A2 => n853, B1 => 
                           REG_6_9_port, B2 => n835, ZN => n267_port);
   U1026 : AOI22_X1 port map( A1 => REG_0_9_port, A2 => n889, B1 => 
                           REG_2_9_port, B2 => n871, ZN => n266_port);
   U1027 : NAND4_X1 port map( A1 => n269_port, A2 => n268_port, A3 => n267_port
                           , A4 => n266_port, ZN => n275_port);
   U1028 : AOI22_X1 port map( A1 => REG_13_9_port, A2 => n781, B1 => 
                           REG_15_9_port, B2 => n763, ZN => n273_port);
   U1029 : AOI22_X1 port map( A1 => REG_9_9_port, A2 => n817, B1 => 
                           REG_11_9_port, B2 => n799, ZN => n272_port);
   U1030 : AOI22_X1 port map( A1 => REG_12_9_port, A2 => n853, B1 => 
                           REG_14_9_port, B2 => n835, ZN => n271_port);
   U1031 : AOI22_X1 port map( A1 => REG_8_9_port, A2 => n889, B1 => 
                           REG_10_9_port, B2 => n871, ZN => n270_port);
   U1032 : NAND4_X1 port map( A1 => n273_port, A2 => n272_port, A3 => n271_port
                           , A4 => n270_port, ZN => n274_port);
   U1033 : AOI22_X1 port map( A1 => n275_port, A2 => n900, B1 => n274_port, B2 
                           => n896, ZN => n276_port);
   U1034 : OAI221_X1 port map( B1 => n908, B2 => n278_port, C1 => n902, C2 => 
                           n277_port, A => n276_port, ZN => N274);
   U1035 : AOI22_X1 port map( A1 => REG_21_10_port, A2 => n781, B1 => 
                           REG_23_10_port, B2 => n763, ZN => n282_port);
   U1036 : AOI22_X1 port map( A1 => REG_17_10_port, A2 => n817, B1 => 
                           REG_19_10_port, B2 => n799, ZN => n281_port);
   U1037 : AOI22_X1 port map( A1 => REG_20_10_port, A2 => n853, B1 => 
                           REG_22_10_port, B2 => n835, ZN => n280_port);
   U1038 : AOI22_X1 port map( A1 => REG_16_10_port, A2 => n889, B1 => 
                           REG_18_10_port, B2 => n871, ZN => n279_port);
   U1039 : AND4_X1 port map( A1 => n282_port, A2 => n281_port, A3 => n280_port,
                           A4 => n279_port, ZN => n299_port);
   U1040 : AOI22_X1 port map( A1 => REG_29_10_port, A2 => n781, B1 => 
                           REG_31_10_port, B2 => n763, ZN => n286_port);
   U1041 : AOI22_X1 port map( A1 => REG_25_10_port, A2 => n817, B1 => 
                           REG_27_10_port, B2 => n799, ZN => n285_port);
   U1042 : AOI22_X1 port map( A1 => REG_28_10_port, A2 => n853, B1 => 
                           REG_30_10_port, B2 => n835, ZN => n284_port);
   U1043 : AOI22_X1 port map( A1 => REG_24_10_port, A2 => n889, B1 => 
                           REG_26_10_port, B2 => n871, ZN => n283_port);
   U1044 : AND4_X1 port map( A1 => n286_port, A2 => n285_port, A3 => n284_port,
                           A4 => n283_port, ZN => n298_port);
   U1045 : AOI22_X1 port map( A1 => REG_5_10_port, A2 => n781, B1 => 
                           REG_7_10_port, B2 => n763, ZN => n290_port);
   U1046 : AOI22_X1 port map( A1 => REG_1_10_port, A2 => n817, B1 => 
                           REG_3_10_port, B2 => n799, ZN => n289_port);
   U1047 : AOI22_X1 port map( A1 => REG_4_10_port, A2 => n853, B1 => 
                           REG_6_10_port, B2 => n835, ZN => n288_port);
   U1048 : AOI22_X1 port map( A1 => REG_0_10_port, A2 => n889, B1 => 
                           REG_2_10_port, B2 => n871, ZN => n287_port);
   U1049 : NAND4_X1 port map( A1 => n290_port, A2 => n289_port, A3 => n288_port
                           , A4 => n287_port, ZN => n296_port);
   U1050 : AOI22_X1 port map( A1 => REG_13_10_port, A2 => n781, B1 => 
                           REG_15_10_port, B2 => n763, ZN => n294_port);
   U1051 : AOI22_X1 port map( A1 => REG_9_10_port, A2 => n817, B1 => 
                           REG_11_10_port, B2 => n799, ZN => n293_port);
   U1052 : AOI22_X1 port map( A1 => REG_12_10_port, A2 => n853, B1 => 
                           REG_14_10_port, B2 => n835, ZN => n292_port);
   U1053 : AOI22_X1 port map( A1 => REG_8_10_port, A2 => n889, B1 => 
                           REG_10_10_port, B2 => n871, ZN => n291_port);
   U1054 : NAND4_X1 port map( A1 => n294_port, A2 => n293_port, A3 => n292_port
                           , A4 => n291_port, ZN => n295_port);
   U1055 : AOI22_X1 port map( A1 => n296_port, A2 => n900, B1 => n295_port, B2 
                           => n896, ZN => n297_port);
   U1056 : OAI221_X1 port map( B1 => n908, B2 => n299_port, C1 => n903, C2 => 
                           n298_port, A => n297_port, ZN => N273);
   U1057 : AOI22_X1 port map( A1 => REG_21_11_port, A2 => n780, B1 => 
                           REG_23_11_port, B2 => n762, ZN => n303_port);
   U1058 : AOI22_X1 port map( A1 => REG_17_11_port, A2 => n816, B1 => 
                           REG_19_11_port, B2 => n798, ZN => n302_port);
   U1059 : AOI22_X1 port map( A1 => REG_20_11_port, A2 => n852, B1 => 
                           REG_22_11_port, B2 => n834, ZN => n301_port);
   U1060 : AOI22_X1 port map( A1 => REG_16_11_port, A2 => n888, B1 => 
                           REG_18_11_port, B2 => n870, ZN => n300_port);
   U1061 : AND4_X1 port map( A1 => n303_port, A2 => n302_port, A3 => n301_port,
                           A4 => n300_port, ZN => n320);
   U1062 : AOI22_X1 port map( A1 => REG_29_11_port, A2 => n780, B1 => 
                           REG_31_11_port, B2 => n762, ZN => n307_port);
   U1063 : AOI22_X1 port map( A1 => REG_25_11_port, A2 => n816, B1 => 
                           REG_27_11_port, B2 => n798, ZN => n306_port);
   U1064 : AOI22_X1 port map( A1 => REG_28_11_port, A2 => n852, B1 => 
                           REG_30_11_port, B2 => n834, ZN => n305_port);
   U1065 : AOI22_X1 port map( A1 => REG_24_11_port, A2 => n888, B1 => 
                           REG_26_11_port, B2 => n870, ZN => n304_port);
   U1066 : AND4_X1 port map( A1 => n307_port, A2 => n306_port, A3 => n305_port,
                           A4 => n304_port, ZN => n319);
   U1067 : AOI22_X1 port map( A1 => REG_5_11_port, A2 => n780, B1 => 
                           REG_7_11_port, B2 => n762, ZN => n311_port);
   U1068 : AOI22_X1 port map( A1 => REG_1_11_port, A2 => n816, B1 => 
                           REG_3_11_port, B2 => n798, ZN => n310_port);
   U1069 : AOI22_X1 port map( A1 => REG_4_11_port, A2 => n852, B1 => 
                           REG_6_11_port, B2 => n834, ZN => n309_port);
   U1070 : AOI22_X1 port map( A1 => REG_0_11_port, A2 => n888, B1 => 
                           REG_2_11_port, B2 => n870, ZN => n308_port);
   U1071 : NAND4_X1 port map( A1 => n311_port, A2 => n310_port, A3 => n309_port
                           , A4 => n308_port, ZN => n317);
   U1072 : AOI22_X1 port map( A1 => REG_13_11_port, A2 => n780, B1 => 
                           REG_15_11_port, B2 => n762, ZN => n315_port);
   U1073 : AOI22_X1 port map( A1 => REG_9_11_port, A2 => n816, B1 => 
                           REG_11_11_port, B2 => n798, ZN => n314_port);
   U1074 : AOI22_X1 port map( A1 => REG_12_11_port, A2 => n852, B1 => 
                           REG_14_11_port, B2 => n834, ZN => n313_port);
   U1075 : AOI22_X1 port map( A1 => REG_8_11_port, A2 => n888, B1 => 
                           REG_10_11_port, B2 => n870, ZN => n312_port);
   U1076 : NAND4_X1 port map( A1 => n315_port, A2 => n314_port, A3 => n313_port
                           , A4 => n312_port, ZN => n316);
   U1077 : AOI22_X1 port map( A1 => n317, A2 => n899, B1 => n316, B2 => n895, 
                           ZN => n318);
   U1078 : OAI221_X1 port map( B1 => n907, B2 => n320, C1 => n903, C2 => n319, 
                           A => n318, ZN => N272);
   U1079 : AOI22_X1 port map( A1 => REG_21_12_port, A2 => n780, B1 => 
                           REG_23_12_port, B2 => n762, ZN => n324);
   U1080 : AOI22_X1 port map( A1 => REG_17_12_port, A2 => n816, B1 => 
                           REG_19_12_port, B2 => n798, ZN => n323);
   U1081 : AOI22_X1 port map( A1 => REG_20_12_port, A2 => n852, B1 => 
                           REG_22_12_port, B2 => n834, ZN => n322);
   U1082 : AOI22_X1 port map( A1 => REG_16_12_port, A2 => n888, B1 => 
                           REG_18_12_port, B2 => n870, ZN => n321);
   U1083 : AND4_X1 port map( A1 => n324, A2 => n323, A3 => n322, A4 => n321, ZN
                           => n341);
   U1084 : AOI22_X1 port map( A1 => REG_29_12_port, A2 => n780, B1 => 
                           REG_31_12_port, B2 => n762, ZN => n328);
   U1085 : AOI22_X1 port map( A1 => REG_25_12_port, A2 => n816, B1 => 
                           REG_27_12_port, B2 => n798, ZN => n327);
   U1086 : AOI22_X1 port map( A1 => REG_28_12_port, A2 => n852, B1 => 
                           REG_30_12_port, B2 => n834, ZN => n326);
   U1087 : AOI22_X1 port map( A1 => REG_24_12_port, A2 => n888, B1 => 
                           REG_26_12_port, B2 => n870, ZN => n325);
   U1088 : AND4_X1 port map( A1 => n328, A2 => n327, A3 => n326, A4 => n325, ZN
                           => n340);
   U1089 : AOI22_X1 port map( A1 => REG_5_12_port, A2 => n780, B1 => 
                           REG_7_12_port, B2 => n762, ZN => n332);
   U1090 : AOI22_X1 port map( A1 => REG_1_12_port, A2 => n816, B1 => 
                           REG_3_12_port, B2 => n798, ZN => n331);
   U1091 : AOI22_X1 port map( A1 => REG_4_12_port, A2 => n852, B1 => 
                           REG_6_12_port, B2 => n834, ZN => n330);
   U1092 : AOI22_X1 port map( A1 => REG_0_12_port, A2 => n888, B1 => 
                           REG_2_12_port, B2 => n870, ZN => n329);
   U1093 : NAND4_X1 port map( A1 => n332, A2 => n331, A3 => n330, A4 => n329, 
                           ZN => n338);
   U1094 : AOI22_X1 port map( A1 => REG_13_12_port, A2 => n780, B1 => 
                           REG_15_12_port, B2 => n762, ZN => n336);
   U1095 : AOI22_X1 port map( A1 => REG_9_12_port, A2 => n816, B1 => 
                           REG_11_12_port, B2 => n798, ZN => n335);
   U1096 : AOI22_X1 port map( A1 => REG_12_12_port, A2 => n852, B1 => 
                           REG_14_12_port, B2 => n834, ZN => n334);
   U1097 : AOI22_X1 port map( A1 => REG_8_12_port, A2 => n888, B1 => 
                           REG_10_12_port, B2 => n870, ZN => n333);
   U1098 : NAND4_X1 port map( A1 => n336, A2 => n335, A3 => n334, A4 => n333, 
                           ZN => n337);
   U1099 : AOI22_X1 port map( A1 => n338, A2 => n899, B1 => n337, B2 => n895, 
                           ZN => n339);
   U1100 : OAI221_X1 port map( B1 => n907, B2 => n341, C1 => n903, C2 => n340, 
                           A => n339, ZN => N271);
   U1101 : AOI22_X1 port map( A1 => REG_21_13_port, A2 => n780, B1 => 
                           REG_23_13_port, B2 => n762, ZN => n345);
   U1102 : AOI22_X1 port map( A1 => REG_17_13_port, A2 => n816, B1 => 
                           REG_19_13_port, B2 => n798, ZN => n344);
   U1103 : AOI22_X1 port map( A1 => REG_20_13_port, A2 => n852, B1 => 
                           REG_22_13_port, B2 => n834, ZN => n343);
   U1104 : AOI22_X1 port map( A1 => REG_16_13_port, A2 => n888, B1 => 
                           REG_18_13_port, B2 => n870, ZN => n342);
   U1105 : AND4_X1 port map( A1 => n345, A2 => n344, A3 => n343, A4 => n342, ZN
                           => n362);
   U1106 : AOI22_X1 port map( A1 => REG_29_13_port, A2 => n780, B1 => 
                           REG_31_13_port, B2 => n762, ZN => n349);
   U1107 : AOI22_X1 port map( A1 => REG_25_13_port, A2 => n816, B1 => 
                           REG_27_13_port, B2 => n798, ZN => n348);
   U1108 : AOI22_X1 port map( A1 => REG_28_13_port, A2 => n852, B1 => 
                           REG_30_13_port, B2 => n834, ZN => n347);
   U1109 : AOI22_X1 port map( A1 => REG_24_13_port, A2 => n888, B1 => 
                           REG_26_13_port, B2 => n870, ZN => n346);
   U1110 : AND4_X1 port map( A1 => n349, A2 => n348, A3 => n347, A4 => n346, ZN
                           => n361);
   U1111 : AOI22_X1 port map( A1 => REG_5_13_port, A2 => n780, B1 => 
                           REG_7_13_port, B2 => n762, ZN => n353);
   U1112 : AOI22_X1 port map( A1 => REG_1_13_port, A2 => n816, B1 => 
                           REG_3_13_port, B2 => n798, ZN => n352);
   U1113 : AOI22_X1 port map( A1 => REG_4_13_port, A2 => n852, B1 => 
                           REG_6_13_port, B2 => n834, ZN => n351);
   U1114 : AOI22_X1 port map( A1 => REG_0_13_port, A2 => n888, B1 => 
                           REG_2_13_port, B2 => n870, ZN => n350);
   U1115 : NAND4_X1 port map( A1 => n353, A2 => n352, A3 => n351, A4 => n350, 
                           ZN => n359);
   U1116 : AOI22_X1 port map( A1 => REG_13_13_port, A2 => n779, B1 => 
                           REG_15_13_port, B2 => n761, ZN => n357);
   U1117 : AOI22_X1 port map( A1 => REG_9_13_port, A2 => n815, B1 => 
                           REG_11_13_port, B2 => n797, ZN => n356);
   U1118 : AOI22_X1 port map( A1 => REG_12_13_port, A2 => n851, B1 => 
                           REG_14_13_port, B2 => n833, ZN => n355);
   U1119 : AOI22_X1 port map( A1 => REG_8_13_port, A2 => n887, B1 => 
                           REG_10_13_port, B2 => n869, ZN => n354);
   U1120 : NAND4_X1 port map( A1 => n357, A2 => n356, A3 => n355, A4 => n354, 
                           ZN => n358);
   U1121 : AOI22_X1 port map( A1 => n359, A2 => n899, B1 => n358, B2 => n895, 
                           ZN => n360);
   U1122 : OAI221_X1 port map( B1 => n907, B2 => n362, C1 => n903, C2 => n361, 
                           A => n360, ZN => N270);
   U1123 : AOI22_X1 port map( A1 => REG_21_14_port, A2 => n779, B1 => 
                           REG_23_14_port, B2 => n761, ZN => n366);
   U1124 : AOI22_X1 port map( A1 => REG_17_14_port, A2 => n815, B1 => 
                           REG_19_14_port, B2 => n797, ZN => n365);
   U1125 : AOI22_X1 port map( A1 => REG_20_14_port, A2 => n851, B1 => 
                           REG_22_14_port, B2 => n833, ZN => n364);
   U1126 : AOI22_X1 port map( A1 => REG_16_14_port, A2 => n887, B1 => 
                           REG_18_14_port, B2 => n869, ZN => n363);
   U1127 : AND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => n383);
   U1128 : AOI22_X1 port map( A1 => REG_29_14_port, A2 => n779, B1 => 
                           REG_31_14_port, B2 => n761, ZN => n370);
   U1129 : AOI22_X1 port map( A1 => REG_25_14_port, A2 => n815, B1 => 
                           REG_27_14_port, B2 => n797, ZN => n369);
   U1130 : AOI22_X1 port map( A1 => REG_28_14_port, A2 => n851, B1 => 
                           REG_30_14_port, B2 => n833, ZN => n368);
   U1131 : AOI22_X1 port map( A1 => REG_24_14_port, A2 => n887, B1 => 
                           REG_26_14_port, B2 => n869, ZN => n367);
   U1132 : AND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => n382);
   U1133 : AOI22_X1 port map( A1 => REG_5_14_port, A2 => n779, B1 => 
                           REG_7_14_port, B2 => n761, ZN => n374);
   U1134 : AOI22_X1 port map( A1 => REG_1_14_port, A2 => n815, B1 => 
                           REG_3_14_port, B2 => n797, ZN => n373);
   U1135 : AOI22_X1 port map( A1 => REG_4_14_port, A2 => n851, B1 => 
                           REG_6_14_port, B2 => n833, ZN => n372);
   U1136 : AOI22_X1 port map( A1 => REG_0_14_port, A2 => n887, B1 => 
                           REG_2_14_port, B2 => n869, ZN => n371);
   U1137 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, 
                           ZN => n380);
   U1138 : AOI22_X1 port map( A1 => REG_13_14_port, A2 => n779, B1 => 
                           REG_15_14_port, B2 => n761, ZN => n378);
   U1139 : AOI22_X1 port map( A1 => REG_9_14_port, A2 => n815, B1 => 
                           REG_11_14_port, B2 => n797, ZN => n377);
   U1140 : AOI22_X1 port map( A1 => REG_12_14_port, A2 => n851, B1 => 
                           REG_14_14_port, B2 => n833, ZN => n376);
   U1141 : AOI22_X1 port map( A1 => REG_8_14_port, A2 => n887, B1 => 
                           REG_10_14_port, B2 => n869, ZN => n375);
   U1142 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, 
                           ZN => n379);
   U1143 : AOI22_X1 port map( A1 => n380, A2 => n899, B1 => n379, B2 => n895, 
                           ZN => n381);
   U1144 : OAI221_X1 port map( B1 => n907, B2 => n383, C1 => n903, C2 => n382, 
                           A => n381, ZN => N269);
   U1145 : AOI22_X1 port map( A1 => REG_21_15_port, A2 => n779, B1 => 
                           REG_23_15_port, B2 => n761, ZN => n387);
   U1146 : AOI22_X1 port map( A1 => REG_17_15_port, A2 => n815, B1 => 
                           REG_19_15_port, B2 => n797, ZN => n386);
   U1147 : AOI22_X1 port map( A1 => REG_20_15_port, A2 => n851, B1 => 
                           REG_22_15_port, B2 => n833, ZN => n385);
   U1148 : AOI22_X1 port map( A1 => REG_16_15_port, A2 => n887, B1 => 
                           REG_18_15_port, B2 => n869, ZN => n384);
   U1149 : AND4_X1 port map( A1 => n387, A2 => n386, A3 => n385, A4 => n384, ZN
                           => n404);
   U1150 : AOI22_X1 port map( A1 => REG_29_15_port, A2 => n779, B1 => 
                           REG_31_15_port, B2 => n761, ZN => n391);
   U1151 : AOI22_X1 port map( A1 => REG_25_15_port, A2 => n815, B1 => 
                           REG_27_15_port, B2 => n797, ZN => n390);
   U1152 : AOI22_X1 port map( A1 => REG_28_15_port, A2 => n851, B1 => 
                           REG_30_15_port, B2 => n833, ZN => n389);
   U1153 : AOI22_X1 port map( A1 => REG_24_15_port, A2 => n887, B1 => 
                           REG_26_15_port, B2 => n869, ZN => n388);
   U1154 : AND4_X1 port map( A1 => n391, A2 => n390, A3 => n389, A4 => n388, ZN
                           => n403);
   U1155 : AOI22_X1 port map( A1 => REG_5_15_port, A2 => n779, B1 => 
                           REG_7_15_port, B2 => n761, ZN => n395);
   U1156 : AOI22_X1 port map( A1 => REG_1_15_port, A2 => n815, B1 => 
                           REG_3_15_port, B2 => n797, ZN => n394);
   U1157 : AOI22_X1 port map( A1 => REG_4_15_port, A2 => n851, B1 => 
                           REG_6_15_port, B2 => n833, ZN => n393);
   U1158 : AOI22_X1 port map( A1 => REG_0_15_port, A2 => n887, B1 => 
                           REG_2_15_port, B2 => n869, ZN => n392);
   U1159 : NAND4_X1 port map( A1 => n395, A2 => n394, A3 => n393, A4 => n392, 
                           ZN => n401);
   U1160 : AOI22_X1 port map( A1 => REG_13_15_port, A2 => n779, B1 => 
                           REG_15_15_port, B2 => n761, ZN => n399);
   U1161 : AOI22_X1 port map( A1 => REG_9_15_port, A2 => n815, B1 => 
                           REG_11_15_port, B2 => n797, ZN => n398);
   U1162 : AOI22_X1 port map( A1 => REG_12_15_port, A2 => n851, B1 => 
                           REG_14_15_port, B2 => n833, ZN => n397);
   U1163 : AOI22_X1 port map( A1 => REG_8_15_port, A2 => n887, B1 => 
                           REG_10_15_port, B2 => n869, ZN => n396);
   U1164 : NAND4_X1 port map( A1 => n399, A2 => n398, A3 => n397, A4 => n396, 
                           ZN => n400);
   U1165 : AOI22_X1 port map( A1 => n401, A2 => n899, B1 => n400, B2 => n895, 
                           ZN => n402);
   U1166 : OAI221_X1 port map( B1 => n907, B2 => n404, C1 => n903, C2 => n403, 
                           A => n402, ZN => N268);
   U1167 : AOI22_X1 port map( A1 => REG_21_16_port, A2 => n779, B1 => 
                           REG_23_16_port, B2 => n761, ZN => n408);
   U1168 : AOI22_X1 port map( A1 => REG_17_16_port, A2 => n815, B1 => 
                           REG_19_16_port, B2 => n797, ZN => n407);
   U1169 : AOI22_X1 port map( A1 => REG_20_16_port, A2 => n851, B1 => 
                           REG_22_16_port, B2 => n833, ZN => n406);
   U1170 : AOI22_X1 port map( A1 => REG_16_16_port, A2 => n887, B1 => 
                           REG_18_16_port, B2 => n869, ZN => n405);
   U1171 : AND4_X1 port map( A1 => n408, A2 => n407, A3 => n406, A4 => n405, ZN
                           => n425);
   U1172 : AOI22_X1 port map( A1 => REG_29_16_port, A2 => n779, B1 => 
                           REG_31_16_port, B2 => n761, ZN => n412);
   U1173 : AOI22_X1 port map( A1 => REG_25_16_port, A2 => n815, B1 => 
                           REG_27_16_port, B2 => n797, ZN => n411);
   U1174 : AOI22_X1 port map( A1 => REG_28_16_port, A2 => n851, B1 => 
                           REG_30_16_port, B2 => n833, ZN => n410);
   U1175 : AOI22_X1 port map( A1 => REG_24_16_port, A2 => n887, B1 => 
                           REG_26_16_port, B2 => n869, ZN => n409);
   U1176 : AND4_X1 port map( A1 => n412, A2 => n411, A3 => n410, A4 => n409, ZN
                           => n424);
   U1177 : AOI22_X1 port map( A1 => REG_5_16_port, A2 => n778, B1 => 
                           REG_7_16_port, B2 => n760, ZN => n416);
   U1178 : AOI22_X1 port map( A1 => REG_1_16_port, A2 => n814, B1 => 
                           REG_3_16_port, B2 => n796, ZN => n415);
   U1179 : AOI22_X1 port map( A1 => REG_4_16_port, A2 => n850, B1 => 
                           REG_6_16_port, B2 => n832, ZN => n414);
   U1180 : AOI22_X1 port map( A1 => REG_0_16_port, A2 => n886, B1 => 
                           REG_2_16_port, B2 => n868, ZN => n413);
   U1181 : NAND4_X1 port map( A1 => n416, A2 => n415, A3 => n414, A4 => n413, 
                           ZN => n422);
   U1182 : AOI22_X1 port map( A1 => REG_13_16_port, A2 => n778, B1 => 
                           REG_15_16_port, B2 => n760, ZN => n420);
   U1183 : AOI22_X1 port map( A1 => REG_9_16_port, A2 => n814, B1 => 
                           REG_11_16_port, B2 => n796, ZN => n419);
   U1184 : AOI22_X1 port map( A1 => REG_12_16_port, A2 => n850, B1 => 
                           REG_14_16_port, B2 => n832, ZN => n418);
   U1185 : AOI22_X1 port map( A1 => REG_8_16_port, A2 => n886, B1 => 
                           REG_10_16_port, B2 => n868, ZN => n417);
   U1186 : NAND4_X1 port map( A1 => n420, A2 => n419, A3 => n418, A4 => n417, 
                           ZN => n421);
   U1187 : AOI22_X1 port map( A1 => n422, A2 => n899, B1 => n421, B2 => n895, 
                           ZN => n423);
   U1188 : OAI221_X1 port map( B1 => n907, B2 => n425, C1 => n903, C2 => n424, 
                           A => n423, ZN => N267);
   U1189 : AOI22_X1 port map( A1 => REG_21_17_port, A2 => n778, B1 => 
                           REG_23_17_port, B2 => n760, ZN => n429);
   U1190 : AOI22_X1 port map( A1 => REG_17_17_port, A2 => n814, B1 => 
                           REG_19_17_port, B2 => n796, ZN => n428);
   U1191 : AOI22_X1 port map( A1 => REG_20_17_port, A2 => n850, B1 => 
                           REG_22_17_port, B2 => n832, ZN => n427);
   U1192 : AOI22_X1 port map( A1 => REG_16_17_port, A2 => n886, B1 => 
                           REG_18_17_port, B2 => n868, ZN => n426);
   U1193 : AND4_X1 port map( A1 => n429, A2 => n428, A3 => n427, A4 => n426, ZN
                           => n446);
   U1194 : AOI22_X1 port map( A1 => REG_29_17_port, A2 => n778, B1 => 
                           REG_31_17_port, B2 => n760, ZN => n433);
   U1195 : AOI22_X1 port map( A1 => REG_25_17_port, A2 => n814, B1 => 
                           REG_27_17_port, B2 => n796, ZN => n432);
   U1196 : AOI22_X1 port map( A1 => REG_28_17_port, A2 => n850, B1 => 
                           REG_30_17_port, B2 => n832, ZN => n431);
   U1197 : AOI22_X1 port map( A1 => REG_24_17_port, A2 => n886, B1 => 
                           REG_26_17_port, B2 => n868, ZN => n430);
   U1198 : AND4_X1 port map( A1 => n433, A2 => n432, A3 => n431, A4 => n430, ZN
                           => n445);
   U1199 : AOI22_X1 port map( A1 => REG_5_17_port, A2 => n778, B1 => 
                           REG_7_17_port, B2 => n760, ZN => n437);
   U1200 : AOI22_X1 port map( A1 => REG_1_17_port, A2 => n814, B1 => 
                           REG_3_17_port, B2 => n796, ZN => n436);
   U1201 : AOI22_X1 port map( A1 => REG_4_17_port, A2 => n850, B1 => 
                           REG_6_17_port, B2 => n832, ZN => n435);
   U1202 : AOI22_X1 port map( A1 => REG_0_17_port, A2 => n886, B1 => 
                           REG_2_17_port, B2 => n868, ZN => n434);
   U1203 : NAND4_X1 port map( A1 => n437, A2 => n436, A3 => n435, A4 => n434, 
                           ZN => n443);
   U1204 : AOI22_X1 port map( A1 => REG_13_17_port, A2 => n778, B1 => 
                           REG_15_17_port, B2 => n760, ZN => n441);
   U1205 : AOI22_X1 port map( A1 => REG_9_17_port, A2 => n814, B1 => 
                           REG_11_17_port, B2 => n796, ZN => n440);
   U1206 : AOI22_X1 port map( A1 => REG_12_17_port, A2 => n850, B1 => 
                           REG_14_17_port, B2 => n832, ZN => n439);
   U1207 : AOI22_X1 port map( A1 => REG_8_17_port, A2 => n886, B1 => 
                           REG_10_17_port, B2 => n868, ZN => n438);
   U1208 : NAND4_X1 port map( A1 => n441, A2 => n440, A3 => n439, A4 => n438, 
                           ZN => n442);
   U1209 : AOI22_X1 port map( A1 => n443, A2 => n899, B1 => n442, B2 => n895, 
                           ZN => n444);
   U1210 : OAI221_X1 port map( B1 => n907, B2 => n446, C1 => n903, C2 => n445, 
                           A => n444, ZN => N266);
   U1211 : AOI22_X1 port map( A1 => REG_21_18_port, A2 => n778, B1 => 
                           REG_23_18_port, B2 => n760, ZN => n450);
   U1212 : AOI22_X1 port map( A1 => REG_17_18_port, A2 => n814, B1 => 
                           REG_19_18_port, B2 => n796, ZN => n449);
   U1213 : AOI22_X1 port map( A1 => REG_20_18_port, A2 => n850, B1 => 
                           REG_22_18_port, B2 => n832, ZN => n448);
   U1214 : AOI22_X1 port map( A1 => REG_16_18_port, A2 => n886, B1 => 
                           REG_18_18_port, B2 => n868, ZN => n447);
   U1215 : AND4_X1 port map( A1 => n450, A2 => n449, A3 => n448, A4 => n447, ZN
                           => n467);
   U1216 : AOI22_X1 port map( A1 => REG_29_18_port, A2 => n778, B1 => 
                           REG_31_18_port, B2 => n760, ZN => n454);
   U1217 : AOI22_X1 port map( A1 => REG_25_18_port, A2 => n814, B1 => 
                           REG_27_18_port, B2 => n796, ZN => n453);
   U1218 : AOI22_X1 port map( A1 => REG_28_18_port, A2 => n850, B1 => 
                           REG_30_18_port, B2 => n832, ZN => n452);
   U1219 : AOI22_X1 port map( A1 => REG_24_18_port, A2 => n886, B1 => 
                           REG_26_18_port, B2 => n868, ZN => n451);
   U1220 : AND4_X1 port map( A1 => n454, A2 => n453, A3 => n452, A4 => n451, ZN
                           => n466);
   U1221 : AOI22_X1 port map( A1 => REG_5_18_port, A2 => n778, B1 => 
                           REG_7_18_port, B2 => n760, ZN => n458);
   U1222 : AOI22_X1 port map( A1 => REG_1_18_port, A2 => n814, B1 => 
                           REG_3_18_port, B2 => n796, ZN => n457);
   U1223 : AOI22_X1 port map( A1 => REG_4_18_port, A2 => n850, B1 => 
                           REG_6_18_port, B2 => n832, ZN => n456);
   U1224 : AOI22_X1 port map( A1 => REG_0_18_port, A2 => n886, B1 => 
                           REG_2_18_port, B2 => n868, ZN => n455);
   U1225 : NAND4_X1 port map( A1 => n458, A2 => n457, A3 => n456, A4 => n455, 
                           ZN => n464);
   U1226 : AOI22_X1 port map( A1 => REG_13_18_port, A2 => n778, B1 => 
                           REG_15_18_port, B2 => n760, ZN => n462);
   U1227 : AOI22_X1 port map( A1 => REG_9_18_port, A2 => n814, B1 => 
                           REG_11_18_port, B2 => n796, ZN => n461);
   U1228 : AOI22_X1 port map( A1 => REG_12_18_port, A2 => n850, B1 => 
                           REG_14_18_port, B2 => n832, ZN => n460);
   U1229 : AOI22_X1 port map( A1 => REG_8_18_port, A2 => n886, B1 => 
                           REG_10_18_port, B2 => n868, ZN => n459);
   U1230 : NAND4_X1 port map( A1 => n462, A2 => n461, A3 => n460, A4 => n459, 
                           ZN => n463);
   U1231 : AOI22_X1 port map( A1 => n464, A2 => n899, B1 => n463, B2 => n895, 
                           ZN => n465);
   U1232 : OAI221_X1 port map( B1 => n907, B2 => n467, C1 => n903, C2 => n466, 
                           A => n465, ZN => N265);
   U1233 : AOI22_X1 port map( A1 => REG_21_19_port, A2 => n778, B1 => 
                           REG_23_19_port, B2 => n760, ZN => n471);
   U1234 : AOI22_X1 port map( A1 => REG_17_19_port, A2 => n814, B1 => 
                           REG_19_19_port, B2 => n796, ZN => n470);
   U1235 : AOI22_X1 port map( A1 => REG_20_19_port, A2 => n850, B1 => 
                           REG_22_19_port, B2 => n832, ZN => n469);
   U1236 : AOI22_X1 port map( A1 => REG_16_19_port, A2 => n886, B1 => 
                           REG_18_19_port, B2 => n868, ZN => n468);
   U1237 : AND4_X1 port map( A1 => n471, A2 => n470, A3 => n469, A4 => n468, ZN
                           => n488);
   U1238 : AOI22_X1 port map( A1 => REG_29_19_port, A2 => n777, B1 => 
                           REG_31_19_port, B2 => n759, ZN => n475);
   U1239 : AOI22_X1 port map( A1 => REG_25_19_port, A2 => n813, B1 => 
                           REG_27_19_port, B2 => n795, ZN => n474);
   U1240 : AOI22_X1 port map( A1 => REG_28_19_port, A2 => n849, B1 => 
                           REG_30_19_port, B2 => n831, ZN => n473);
   U1241 : AOI22_X1 port map( A1 => REG_24_19_port, A2 => n885, B1 => 
                           REG_26_19_port, B2 => n867, ZN => n472);
   U1242 : AND4_X1 port map( A1 => n475, A2 => n474, A3 => n473, A4 => n472, ZN
                           => n487);
   U1243 : AOI22_X1 port map( A1 => REG_5_19_port, A2 => n777, B1 => 
                           REG_7_19_port, B2 => n759, ZN => n479);
   U1244 : AOI22_X1 port map( A1 => REG_1_19_port, A2 => n813, B1 => 
                           REG_3_19_port, B2 => n795, ZN => n478);
   U1245 : AOI22_X1 port map( A1 => REG_4_19_port, A2 => n849, B1 => 
                           REG_6_19_port, B2 => n831, ZN => n477);
   U1246 : AOI22_X1 port map( A1 => REG_0_19_port, A2 => n885, B1 => 
                           REG_2_19_port, B2 => n867, ZN => n476);
   U1247 : NAND4_X1 port map( A1 => n479, A2 => n478, A3 => n477, A4 => n476, 
                           ZN => n485);
   U1248 : AOI22_X1 port map( A1 => REG_13_19_port, A2 => n777, B1 => 
                           REG_15_19_port, B2 => n759, ZN => n483);
   U1249 : AOI22_X1 port map( A1 => REG_9_19_port, A2 => n813, B1 => 
                           REG_11_19_port, B2 => n795, ZN => n482);
   U1250 : AOI22_X1 port map( A1 => REG_12_19_port, A2 => n849, B1 => 
                           REG_14_19_port, B2 => n831, ZN => n481);
   U1251 : AOI22_X1 port map( A1 => REG_8_19_port, A2 => n885, B1 => 
                           REG_10_19_port, B2 => n867, ZN => n480);
   U1252 : NAND4_X1 port map( A1 => n483, A2 => n482, A3 => n481, A4 => n480, 
                           ZN => n484);
   U1253 : AOI22_X1 port map( A1 => n485, A2 => n899, B1 => n484, B2 => n895, 
                           ZN => n486);
   U1254 : OAI221_X1 port map( B1 => n907, B2 => n488, C1 => n903, C2 => n487, 
                           A => n486, ZN => N264);
   U1255 : AOI22_X1 port map( A1 => REG_21_20_port, A2 => n777, B1 => 
                           REG_23_20_port, B2 => n759, ZN => n492);
   U1256 : AOI22_X1 port map( A1 => REG_17_20_port, A2 => n813, B1 => 
                           REG_19_20_port, B2 => n795, ZN => n491);
   U1257 : AOI22_X1 port map( A1 => REG_20_20_port, A2 => n849, B1 => 
                           REG_22_20_port, B2 => n831, ZN => n490);
   U1258 : AOI22_X1 port map( A1 => REG_16_20_port, A2 => n885, B1 => 
                           REG_18_20_port, B2 => n867, ZN => n489);
   U1259 : AND4_X1 port map( A1 => n492, A2 => n491, A3 => n490, A4 => n489, ZN
                           => n509);
   U1260 : AOI22_X1 port map( A1 => REG_29_20_port, A2 => n777, B1 => 
                           REG_31_20_port, B2 => n759, ZN => n496);
   U1261 : AOI22_X1 port map( A1 => REG_25_20_port, A2 => n813, B1 => 
                           REG_27_20_port, B2 => n795, ZN => n495);
   U1262 : AOI22_X1 port map( A1 => REG_28_20_port, A2 => n849, B1 => 
                           REG_30_20_port, B2 => n831, ZN => n494);
   U1263 : AOI22_X1 port map( A1 => REG_24_20_port, A2 => n885, B1 => 
                           REG_26_20_port, B2 => n867, ZN => n493);
   U1264 : AND4_X1 port map( A1 => n496, A2 => n495, A3 => n494, A4 => n493, ZN
                           => n508);
   U1265 : AOI22_X1 port map( A1 => REG_5_20_port, A2 => n777, B1 => 
                           REG_7_20_port, B2 => n759, ZN => n500);
   U1266 : AOI22_X1 port map( A1 => REG_1_20_port, A2 => n813, B1 => 
                           REG_3_20_port, B2 => n795, ZN => n499);
   U1267 : AOI22_X1 port map( A1 => REG_4_20_port, A2 => n849, B1 => 
                           REG_6_20_port, B2 => n831, ZN => n498);
   U1268 : AOI22_X1 port map( A1 => REG_0_20_port, A2 => n885, B1 => 
                           REG_2_20_port, B2 => n867, ZN => n497);
   U1269 : NAND4_X1 port map( A1 => n500, A2 => n499, A3 => n498, A4 => n497, 
                           ZN => n506);
   U1270 : AOI22_X1 port map( A1 => REG_13_20_port, A2 => n777, B1 => 
                           REG_15_20_port, B2 => n759, ZN => n504);
   U1271 : AOI22_X1 port map( A1 => REG_9_20_port, A2 => n813, B1 => 
                           REG_11_20_port, B2 => n795, ZN => n503);
   U1272 : AOI22_X1 port map( A1 => REG_12_20_port, A2 => n849, B1 => 
                           REG_14_20_port, B2 => n831, ZN => n502);
   U1273 : AOI22_X1 port map( A1 => REG_8_20_port, A2 => n885, B1 => 
                           REG_10_20_port, B2 => n867, ZN => n501);
   U1274 : NAND4_X1 port map( A1 => n504, A2 => n503, A3 => n502, A4 => n501, 
                           ZN => n505);
   U1275 : AOI22_X1 port map( A1 => n506, A2 => n899, B1 => n505, B2 => n895, 
                           ZN => n507);
   U1276 : OAI221_X1 port map( B1 => n907, B2 => n509, C1 => n903, C2 => n508, 
                           A => n507, ZN => N263);
   U1277 : AOI22_X1 port map( A1 => REG_21_21_port, A2 => n777, B1 => 
                           REG_23_21_port, B2 => n759, ZN => n513);
   U1278 : AOI22_X1 port map( A1 => REG_17_21_port, A2 => n813, B1 => 
                           REG_19_21_port, B2 => n795, ZN => n512);
   U1279 : AOI22_X1 port map( A1 => REG_20_21_port, A2 => n849, B1 => 
                           REG_22_21_port, B2 => n831, ZN => n511);
   U1280 : AOI22_X1 port map( A1 => REG_16_21_port, A2 => n885, B1 => 
                           REG_18_21_port, B2 => n867, ZN => n510);
   U1281 : AND4_X1 port map( A1 => n513, A2 => n512, A3 => n511, A4 => n510, ZN
                           => n530);
   U1282 : AOI22_X1 port map( A1 => REG_29_21_port, A2 => n777, B1 => 
                           REG_31_21_port, B2 => n759, ZN => n517);
   U1283 : AOI22_X1 port map( A1 => REG_25_21_port, A2 => n813, B1 => 
                           REG_27_21_port, B2 => n795, ZN => n516);
   U1284 : AOI22_X1 port map( A1 => REG_28_21_port, A2 => n849, B1 => 
                           REG_30_21_port, B2 => n831, ZN => n515);
   U1285 : AOI22_X1 port map( A1 => REG_24_21_port, A2 => n885, B1 => 
                           REG_26_21_port, B2 => n867, ZN => n514);
   U1286 : AND4_X1 port map( A1 => n517, A2 => n516, A3 => n515, A4 => n514, ZN
                           => n529);
   U1287 : AOI22_X1 port map( A1 => REG_5_21_port, A2 => n777, B1 => 
                           REG_7_21_port, B2 => n759, ZN => n521);
   U1288 : AOI22_X1 port map( A1 => REG_1_21_port, A2 => n813, B1 => 
                           REG_3_21_port, B2 => n795, ZN => n520);
   U1289 : AOI22_X1 port map( A1 => REG_4_21_port, A2 => n849, B1 => 
                           REG_6_21_port, B2 => n831, ZN => n519);
   U1290 : AOI22_X1 port map( A1 => REG_0_21_port, A2 => n885, B1 => 
                           REG_2_21_port, B2 => n867, ZN => n518);
   U1291 : NAND4_X1 port map( A1 => n521, A2 => n520, A3 => n519, A4 => n518, 
                           ZN => n527);
   U1292 : AOI22_X1 port map( A1 => REG_13_21_port, A2 => n777, B1 => 
                           REG_15_21_port, B2 => n759, ZN => n525);
   U1293 : AOI22_X1 port map( A1 => REG_9_21_port, A2 => n813, B1 => 
                           REG_11_21_port, B2 => n795, ZN => n524);
   U1294 : AOI22_X1 port map( A1 => REG_12_21_port, A2 => n849, B1 => 
                           REG_14_21_port, B2 => n831, ZN => n523);
   U1295 : AOI22_X1 port map( A1 => REG_8_21_port, A2 => n885, B1 => 
                           REG_10_21_port, B2 => n867, ZN => n522);
   U1296 : NAND4_X1 port map( A1 => n525, A2 => n524, A3 => n523, A4 => n522, 
                           ZN => n526);
   U1297 : AOI22_X1 port map( A1 => n527, A2 => n899, B1 => n526, B2 => n895, 
                           ZN => n528);
   U1298 : OAI221_X1 port map( B1 => n907, B2 => n530, C1 => n904, C2 => n529, 
                           A => n528, ZN => N262);
   U1299 : AOI22_X1 port map( A1 => REG_21_22_port, A2 => n776, B1 => 
                           REG_23_22_port, B2 => n758, ZN => n534);
   U1300 : AOI22_X1 port map( A1 => REG_17_22_port, A2 => n812, B1 => 
                           REG_19_22_port, B2 => n794, ZN => n533);
   U1301 : AOI22_X1 port map( A1 => REG_20_22_port, A2 => n848, B1 => 
                           REG_22_22_port, B2 => n830, ZN => n532);
   U1302 : AOI22_X1 port map( A1 => REG_16_22_port, A2 => n884, B1 => 
                           REG_18_22_port, B2 => n866, ZN => n531);
   U1303 : AND4_X1 port map( A1 => n534, A2 => n533, A3 => n532, A4 => n531, ZN
                           => n551);
   U1304 : AOI22_X1 port map( A1 => REG_29_22_port, A2 => n776, B1 => 
                           REG_31_22_port, B2 => n758, ZN => n538);
   U1305 : AOI22_X1 port map( A1 => REG_25_22_port, A2 => n812, B1 => 
                           REG_27_22_port, B2 => n794, ZN => n537);
   U1306 : AOI22_X1 port map( A1 => REG_28_22_port, A2 => n848, B1 => 
                           REG_30_22_port, B2 => n830, ZN => n536);
   U1307 : AOI22_X1 port map( A1 => REG_24_22_port, A2 => n884, B1 => 
                           REG_26_22_port, B2 => n866, ZN => n535);
   U1308 : AND4_X1 port map( A1 => n538, A2 => n537, A3 => n536, A4 => n535, ZN
                           => n550);
   U1309 : AOI22_X1 port map( A1 => REG_5_22_port, A2 => n776, B1 => 
                           REG_7_22_port, B2 => n758, ZN => n542);
   U1310 : AOI22_X1 port map( A1 => REG_1_22_port, A2 => n812, B1 => 
                           REG_3_22_port, B2 => n794, ZN => n541);
   U1311 : AOI22_X1 port map( A1 => REG_4_22_port, A2 => n848, B1 => 
                           REG_6_22_port, B2 => n830, ZN => n540);
   U1312 : AOI22_X1 port map( A1 => REG_0_22_port, A2 => n884, B1 => 
                           REG_2_22_port, B2 => n866, ZN => n539);
   U1313 : NAND4_X1 port map( A1 => n542, A2 => n541, A3 => n540, A4 => n539, 
                           ZN => n548);
   U1314 : AOI22_X1 port map( A1 => REG_13_22_port, A2 => n776, B1 => 
                           REG_15_22_port, B2 => n758, ZN => n546);
   U1315 : AOI22_X1 port map( A1 => REG_9_22_port, A2 => n812, B1 => 
                           REG_11_22_port, B2 => n794, ZN => n545);
   U1316 : AOI22_X1 port map( A1 => REG_12_22_port, A2 => n848, B1 => 
                           REG_14_22_port, B2 => n830, ZN => n544);
   U1317 : AOI22_X1 port map( A1 => REG_8_22_port, A2 => n884, B1 => 
                           REG_10_22_port, B2 => n866, ZN => n543);
   U1318 : NAND4_X1 port map( A1 => n546, A2 => n545, A3 => n544, A4 => n543, 
                           ZN => n547);
   U1319 : AOI22_X1 port map( A1 => n548, A2 => n898, B1 => n547, B2 => n894, 
                           ZN => n549);
   U1320 : OAI221_X1 port map( B1 => n906, B2 => n551, C1 => n904, C2 => n550, 
                           A => n549, ZN => N261);
   U1321 : AOI22_X1 port map( A1 => REG_21_23_port, A2 => n776, B1 => 
                           REG_23_23_port, B2 => n758, ZN => n555);
   U1322 : AOI22_X1 port map( A1 => REG_17_23_port, A2 => n812, B1 => 
                           REG_19_23_port, B2 => n794, ZN => n554);
   U1323 : AOI22_X1 port map( A1 => REG_20_23_port, A2 => n848, B1 => 
                           REG_22_23_port, B2 => n830, ZN => n553);
   U1324 : AOI22_X1 port map( A1 => REG_16_23_port, A2 => n884, B1 => 
                           REG_18_23_port, B2 => n866, ZN => n552);
   U1325 : AND4_X1 port map( A1 => n555, A2 => n554, A3 => n553, A4 => n552, ZN
                           => n572);
   U1326 : AOI22_X1 port map( A1 => REG_29_23_port, A2 => n776, B1 => 
                           REG_31_23_port, B2 => n758, ZN => n559);
   U1327 : AOI22_X1 port map( A1 => REG_25_23_port, A2 => n812, B1 => 
                           REG_27_23_port, B2 => n794, ZN => n558);
   U1328 : AOI22_X1 port map( A1 => REG_28_23_port, A2 => n848, B1 => 
                           REG_30_23_port, B2 => n830, ZN => n557);
   U1329 : AOI22_X1 port map( A1 => REG_24_23_port, A2 => n884, B1 => 
                           REG_26_23_port, B2 => n866, ZN => n556);
   U1330 : AND4_X1 port map( A1 => n559, A2 => n558, A3 => n557, A4 => n556, ZN
                           => n571);
   U1331 : AOI22_X1 port map( A1 => REG_5_23_port, A2 => n776, B1 => 
                           REG_7_23_port, B2 => n758, ZN => n563);
   U1332 : AOI22_X1 port map( A1 => REG_1_23_port, A2 => n812, B1 => 
                           REG_3_23_port, B2 => n794, ZN => n562);
   U1333 : AOI22_X1 port map( A1 => REG_4_23_port, A2 => n848, B1 => 
                           REG_6_23_port, B2 => n830, ZN => n561);
   U1334 : AOI22_X1 port map( A1 => REG_0_23_port, A2 => n884, B1 => 
                           REG_2_23_port, B2 => n866, ZN => n560);
   U1335 : NAND4_X1 port map( A1 => n563, A2 => n562, A3 => n561, A4 => n560, 
                           ZN => n569);
   U1336 : AOI22_X1 port map( A1 => REG_13_23_port, A2 => n776, B1 => 
                           REG_15_23_port, B2 => n758, ZN => n567);
   U1337 : AOI22_X1 port map( A1 => REG_9_23_port, A2 => n812, B1 => 
                           REG_11_23_port, B2 => n794, ZN => n566);
   U1338 : AOI22_X1 port map( A1 => REG_12_23_port, A2 => n848, B1 => 
                           REG_14_23_port, B2 => n830, ZN => n565);
   U1339 : AOI22_X1 port map( A1 => REG_8_23_port, A2 => n884, B1 => 
                           REG_10_23_port, B2 => n866, ZN => n564);
   U1340 : NAND4_X1 port map( A1 => n567, A2 => n566, A3 => n565, A4 => n564, 
                           ZN => n568);
   U1341 : AOI22_X1 port map( A1 => n569, A2 => n898, B1 => n568, B2 => n894, 
                           ZN => n570);
   U1342 : OAI221_X1 port map( B1 => n906, B2 => n572, C1 => n904, C2 => n571, 
                           A => n570, ZN => N260);
   U1343 : AOI22_X1 port map( A1 => REG_21_24_port, A2 => n776, B1 => 
                           REG_23_24_port, B2 => n758, ZN => n576);
   U1344 : AOI22_X1 port map( A1 => REG_17_24_port, A2 => n812, B1 => 
                           REG_19_24_port, B2 => n794, ZN => n575);
   U1345 : AOI22_X1 port map( A1 => REG_20_24_port, A2 => n848, B1 => 
                           REG_22_24_port, B2 => n830, ZN => n574);
   U1346 : AOI22_X1 port map( A1 => REG_16_24_port, A2 => n884, B1 => 
                           REG_18_24_port, B2 => n866, ZN => n573);
   U1347 : AND4_X1 port map( A1 => n576, A2 => n575, A3 => n574, A4 => n573, ZN
                           => n593);
   U1348 : AOI22_X1 port map( A1 => REG_29_24_port, A2 => n776, B1 => 
                           REG_31_24_port, B2 => n758, ZN => n580);
   U1349 : AOI22_X1 port map( A1 => REG_25_24_port, A2 => n812, B1 => 
                           REG_27_24_port, B2 => n794, ZN => n579);
   U1350 : AOI22_X1 port map( A1 => REG_28_24_port, A2 => n848, B1 => 
                           REG_30_24_port, B2 => n830, ZN => n578);
   U1351 : AOI22_X1 port map( A1 => REG_24_24_port, A2 => n884, B1 => 
                           REG_26_24_port, B2 => n866, ZN => n577);
   U1352 : AND4_X1 port map( A1 => n580, A2 => n579, A3 => n578, A4 => n577, ZN
                           => n592);
   U1353 : AOI22_X1 port map( A1 => REG_5_24_port, A2 => n776, B1 => 
                           REG_7_24_port, B2 => n758, ZN => n584);
   U1354 : AOI22_X1 port map( A1 => REG_1_24_port, A2 => n812, B1 => 
                           REG_3_24_port, B2 => n794, ZN => n583);
   U1355 : AOI22_X1 port map( A1 => REG_4_24_port, A2 => n848, B1 => 
                           REG_6_24_port, B2 => n830, ZN => n582);
   U1356 : AOI22_X1 port map( A1 => REG_0_24_port, A2 => n884, B1 => 
                           REG_2_24_port, B2 => n866, ZN => n581);
   U1357 : NAND4_X1 port map( A1 => n584, A2 => n583, A3 => n582, A4 => n581, 
                           ZN => n590);
   U1358 : AOI22_X1 port map( A1 => REG_13_24_port, A2 => n775, B1 => 
                           REG_15_24_port, B2 => n757, ZN => n588);
   U1359 : AOI22_X1 port map( A1 => REG_9_24_port, A2 => n811, B1 => 
                           REG_11_24_port, B2 => n793, ZN => n587);
   U1360 : AOI22_X1 port map( A1 => REG_12_24_port, A2 => n847, B1 => 
                           REG_14_24_port, B2 => n829, ZN => n586);
   U1361 : AOI22_X1 port map( A1 => REG_8_24_port, A2 => n883, B1 => 
                           REG_10_24_port, B2 => n865, ZN => n585);
   U1362 : NAND4_X1 port map( A1 => n588, A2 => n587, A3 => n586, A4 => n585, 
                           ZN => n589);
   U1363 : AOI22_X1 port map( A1 => n590, A2 => n898, B1 => n589, B2 => n894, 
                           ZN => n591);
   U1364 : OAI221_X1 port map( B1 => n906, B2 => n593, C1 => n904, C2 => n592, 
                           A => n591, ZN => N259);
   U1365 : AOI22_X1 port map( A1 => REG_21_25_port, A2 => n775, B1 => 
                           REG_23_25_port, B2 => n757, ZN => n597);
   U1366 : AOI22_X1 port map( A1 => REG_17_25_port, A2 => n811, B1 => 
                           REG_19_25_port, B2 => n793, ZN => n596);
   U1367 : AOI22_X1 port map( A1 => REG_20_25_port, A2 => n847, B1 => 
                           REG_22_25_port, B2 => n829, ZN => n595);
   U1368 : AOI22_X1 port map( A1 => REG_16_25_port, A2 => n883, B1 => 
                           REG_18_25_port, B2 => n865, ZN => n594);
   U1369 : AND4_X1 port map( A1 => n597, A2 => n596, A3 => n595, A4 => n594, ZN
                           => n614);
   U1370 : AOI22_X1 port map( A1 => REG_29_25_port, A2 => n775, B1 => 
                           REG_31_25_port, B2 => n757, ZN => n601);
   U1371 : AOI22_X1 port map( A1 => REG_25_25_port, A2 => n811, B1 => 
                           REG_27_25_port, B2 => n793, ZN => n600);
   U1372 : AOI22_X1 port map( A1 => REG_28_25_port, A2 => n847, B1 => 
                           REG_30_25_port, B2 => n829, ZN => n599);
   U1373 : AOI22_X1 port map( A1 => REG_24_25_port, A2 => n883, B1 => 
                           REG_26_25_port, B2 => n865, ZN => n598);
   U1374 : AND4_X1 port map( A1 => n601, A2 => n600, A3 => n599, A4 => n598, ZN
                           => n613);
   U1375 : AOI22_X1 port map( A1 => REG_5_25_port, A2 => n775, B1 => 
                           REG_7_25_port, B2 => n757, ZN => n605);
   U1376 : AOI22_X1 port map( A1 => REG_1_25_port, A2 => n811, B1 => 
                           REG_3_25_port, B2 => n793, ZN => n604);
   U1377 : AOI22_X1 port map( A1 => REG_4_25_port, A2 => n847, B1 => 
                           REG_6_25_port, B2 => n829, ZN => n603);
   U1378 : AOI22_X1 port map( A1 => REG_0_25_port, A2 => n883, B1 => 
                           REG_2_25_port, B2 => n865, ZN => n602);
   U1379 : NAND4_X1 port map( A1 => n605, A2 => n604, A3 => n603, A4 => n602, 
                           ZN => n611);
   U1380 : AOI22_X1 port map( A1 => REG_13_25_port, A2 => n775, B1 => 
                           REG_15_25_port, B2 => n757, ZN => n609);
   U1381 : AOI22_X1 port map( A1 => REG_9_25_port, A2 => n811, B1 => 
                           REG_11_25_port, B2 => n793, ZN => n608);
   U1382 : AOI22_X1 port map( A1 => REG_12_25_port, A2 => n847, B1 => 
                           REG_14_25_port, B2 => n829, ZN => n607);
   U1383 : AOI22_X1 port map( A1 => REG_8_25_port, A2 => n883, B1 => 
                           REG_10_25_port, B2 => n865, ZN => n606);
   U1384 : NAND4_X1 port map( A1 => n609, A2 => n608, A3 => n607, A4 => n606, 
                           ZN => n610);
   U1385 : AOI22_X1 port map( A1 => n611, A2 => n898, B1 => n610, B2 => n894, 
                           ZN => n612);
   U1386 : OAI221_X1 port map( B1 => n906, B2 => n614, C1 => n904, C2 => n613, 
                           A => n612, ZN => N258);
   U1387 : AOI22_X1 port map( A1 => REG_21_26_port, A2 => n775, B1 => 
                           REG_23_26_port, B2 => n757, ZN => n618);
   U1388 : AOI22_X1 port map( A1 => REG_17_26_port, A2 => n811, B1 => 
                           REG_19_26_port, B2 => n793, ZN => n617);
   U1389 : AOI22_X1 port map( A1 => REG_20_26_port, A2 => n847, B1 => 
                           REG_22_26_port, B2 => n829, ZN => n616);
   U1390 : AOI22_X1 port map( A1 => REG_16_26_port, A2 => n883, B1 => 
                           REG_18_26_port, B2 => n865, ZN => n615);
   U1391 : AND4_X1 port map( A1 => n618, A2 => n617, A3 => n616, A4 => n615, ZN
                           => n635);
   U1392 : AOI22_X1 port map( A1 => REG_29_26_port, A2 => n775, B1 => 
                           REG_31_26_port, B2 => n757, ZN => n622);
   U1393 : AOI22_X1 port map( A1 => REG_25_26_port, A2 => n811, B1 => 
                           REG_27_26_port, B2 => n793, ZN => n621);
   U1394 : AOI22_X1 port map( A1 => REG_28_26_port, A2 => n847, B1 => 
                           REG_30_26_port, B2 => n829, ZN => n620);
   U1395 : AOI22_X1 port map( A1 => REG_24_26_port, A2 => n883, B1 => 
                           REG_26_26_port, B2 => n865, ZN => n619);
   U1396 : AND4_X1 port map( A1 => n622, A2 => n621, A3 => n620, A4 => n619, ZN
                           => n634);
   U1397 : AOI22_X1 port map( A1 => REG_5_26_port, A2 => n775, B1 => 
                           REG_7_26_port, B2 => n757, ZN => n626);
   U1398 : AOI22_X1 port map( A1 => REG_1_26_port, A2 => n811, B1 => 
                           REG_3_26_port, B2 => n793, ZN => n625);
   U1399 : AOI22_X1 port map( A1 => REG_4_26_port, A2 => n847, B1 => 
                           REG_6_26_port, B2 => n829, ZN => n624);
   U1400 : AOI22_X1 port map( A1 => REG_0_26_port, A2 => n883, B1 => 
                           REG_2_26_port, B2 => n865, ZN => n623);
   U1401 : NAND4_X1 port map( A1 => n626, A2 => n625, A3 => n624, A4 => n623, 
                           ZN => n632);
   U1402 : AOI22_X1 port map( A1 => REG_13_26_port, A2 => n775, B1 => 
                           REG_15_26_port, B2 => n757, ZN => n630);
   U1403 : AOI22_X1 port map( A1 => REG_9_26_port, A2 => n811, B1 => 
                           REG_11_26_port, B2 => n793, ZN => n629);
   U1404 : AOI22_X1 port map( A1 => REG_12_26_port, A2 => n847, B1 => 
                           REG_14_26_port, B2 => n829, ZN => n628);
   U1405 : AOI22_X1 port map( A1 => REG_8_26_port, A2 => n883, B1 => 
                           REG_10_26_port, B2 => n865, ZN => n627);
   U1406 : NAND4_X1 port map( A1 => n630, A2 => n629, A3 => n628, A4 => n627, 
                           ZN => n631);
   U1407 : AOI22_X1 port map( A1 => n632, A2 => n898, B1 => n631, B2 => n894, 
                           ZN => n633);
   U1408 : OAI221_X1 port map( B1 => n906, B2 => n635, C1 => n904, C2 => n634, 
                           A => n633, ZN => N257);
   U1409 : AOI22_X1 port map( A1 => REG_21_27_port, A2 => n775, B1 => 
                           REG_23_27_port, B2 => n757, ZN => n639);
   U1410 : AOI22_X1 port map( A1 => REG_17_27_port, A2 => n811, B1 => 
                           REG_19_27_port, B2 => n793, ZN => n638);
   U1411 : AOI22_X1 port map( A1 => REG_20_27_port, A2 => n847, B1 => 
                           REG_22_27_port, B2 => n829, ZN => n637);
   U1412 : AOI22_X1 port map( A1 => REG_16_27_port, A2 => n883, B1 => 
                           REG_18_27_port, B2 => n865, ZN => n636);
   U1413 : AND4_X1 port map( A1 => n639, A2 => n638, A3 => n637, A4 => n636, ZN
                           => n656);
   U1414 : AOI22_X1 port map( A1 => REG_29_27_port, A2 => n775, B1 => 
                           REG_31_27_port, B2 => n757, ZN => n643);
   U1415 : AOI22_X1 port map( A1 => REG_25_27_port, A2 => n811, B1 => 
                           REG_27_27_port, B2 => n793, ZN => n642);
   U1416 : AOI22_X1 port map( A1 => REG_28_27_port, A2 => n847, B1 => 
                           REG_30_27_port, B2 => n829, ZN => n641);
   U1417 : AOI22_X1 port map( A1 => REG_24_27_port, A2 => n883, B1 => 
                           REG_26_27_port, B2 => n865, ZN => n640);
   U1418 : AND4_X1 port map( A1 => n643, A2 => n642, A3 => n641, A4 => n640, ZN
                           => n655);
   U1419 : AOI22_X1 port map( A1 => REG_5_27_port, A2 => n774, B1 => 
                           REG_7_27_port, B2 => n756, ZN => n647);
   U1420 : AOI22_X1 port map( A1 => REG_1_27_port, A2 => n810, B1 => 
                           REG_3_27_port, B2 => n792, ZN => n646);
   U1421 : AOI22_X1 port map( A1 => REG_4_27_port, A2 => n846, B1 => 
                           REG_6_27_port, B2 => n828, ZN => n645);
   U1422 : AOI22_X1 port map( A1 => REG_0_27_port, A2 => n882, B1 => 
                           REG_2_27_port, B2 => n864, ZN => n644);
   U1423 : NAND4_X1 port map( A1 => n647, A2 => n646, A3 => n645, A4 => n644, 
                           ZN => n653);
   U1424 : AOI22_X1 port map( A1 => REG_13_27_port, A2 => n774, B1 => 
                           REG_15_27_port, B2 => n756, ZN => n651);
   U1425 : AOI22_X1 port map( A1 => REG_9_27_port, A2 => n810, B1 => 
                           REG_11_27_port, B2 => n792, ZN => n650);
   U1426 : AOI22_X1 port map( A1 => REG_12_27_port, A2 => n846, B1 => 
                           REG_14_27_port, B2 => n828, ZN => n649);
   U1427 : AOI22_X1 port map( A1 => REG_8_27_port, A2 => n882, B1 => 
                           REG_10_27_port, B2 => n864, ZN => n648);
   U1428 : NAND4_X1 port map( A1 => n651, A2 => n650, A3 => n649, A4 => n648, 
                           ZN => n652);
   U1429 : AOI22_X1 port map( A1 => n653, A2 => n898, B1 => n652, B2 => n894, 
                           ZN => n654);
   U1430 : OAI221_X1 port map( B1 => n906, B2 => n656, C1 => n904, C2 => n655, 
                           A => n654, ZN => N256);
   U1431 : AOI22_X1 port map( A1 => REG_21_28_port, A2 => n774, B1 => 
                           REG_23_28_port, B2 => n756, ZN => n660);
   U1432 : AOI22_X1 port map( A1 => REG_17_28_port, A2 => n810, B1 => 
                           REG_19_28_port, B2 => n792, ZN => n659);
   U1433 : AOI22_X1 port map( A1 => REG_20_28_port, A2 => n846, B1 => 
                           REG_22_28_port, B2 => n828, ZN => n658);
   U1434 : AOI22_X1 port map( A1 => REG_16_28_port, A2 => n882, B1 => 
                           REG_18_28_port, B2 => n864, ZN => n657);
   U1435 : AND4_X1 port map( A1 => n660, A2 => n659, A3 => n658, A4 => n657, ZN
                           => n677);
   U1436 : AOI22_X1 port map( A1 => REG_29_28_port, A2 => n774, B1 => 
                           REG_31_28_port, B2 => n756, ZN => n664);
   U1437 : AOI22_X1 port map( A1 => REG_25_28_port, A2 => n810, B1 => 
                           REG_27_28_port, B2 => n792, ZN => n663);
   U1438 : AOI22_X1 port map( A1 => REG_28_28_port, A2 => n846, B1 => 
                           REG_30_28_port, B2 => n828, ZN => n662);
   U1439 : AOI22_X1 port map( A1 => REG_24_28_port, A2 => n882, B1 => 
                           REG_26_28_port, B2 => n864, ZN => n661);
   U1440 : AND4_X1 port map( A1 => n664, A2 => n663, A3 => n662, A4 => n661, ZN
                           => n676);
   U1441 : AOI22_X1 port map( A1 => REG_5_28_port, A2 => n774, B1 => 
                           REG_7_28_port, B2 => n756, ZN => n668);
   U1442 : AOI22_X1 port map( A1 => REG_1_28_port, A2 => n810, B1 => 
                           REG_3_28_port, B2 => n792, ZN => n667);
   U1443 : AOI22_X1 port map( A1 => REG_4_28_port, A2 => n846, B1 => 
                           REG_6_28_port, B2 => n828, ZN => n666);
   U1444 : AOI22_X1 port map( A1 => REG_0_28_port, A2 => n882, B1 => 
                           REG_2_28_port, B2 => n864, ZN => n665);
   U1445 : NAND4_X1 port map( A1 => n668, A2 => n667, A3 => n666, A4 => n665, 
                           ZN => n674);
   U1446 : AOI22_X1 port map( A1 => REG_13_28_port, A2 => n774, B1 => 
                           REG_15_28_port, B2 => n756, ZN => n672);
   U1447 : AOI22_X1 port map( A1 => REG_9_28_port, A2 => n810, B1 => 
                           REG_11_28_port, B2 => n792, ZN => n671);
   U1448 : AOI22_X1 port map( A1 => REG_12_28_port, A2 => n846, B1 => 
                           REG_14_28_port, B2 => n828, ZN => n670);
   U1449 : AOI22_X1 port map( A1 => REG_8_28_port, A2 => n882, B1 => 
                           REG_10_28_port, B2 => n864, ZN => n669);
   U1450 : NAND4_X1 port map( A1 => n672, A2 => n671, A3 => n670, A4 => n669, 
                           ZN => n673);
   U1451 : AOI22_X1 port map( A1 => n674, A2 => n898, B1 => n673, B2 => n894, 
                           ZN => n675);
   U1452 : OAI221_X1 port map( B1 => n906, B2 => n677, C1 => n904, C2 => n676, 
                           A => n675, ZN => N255);
   U1453 : AOI22_X1 port map( A1 => REG_21_29_port, A2 => n774, B1 => 
                           REG_23_29_port, B2 => n756, ZN => n681);
   U1454 : AOI22_X1 port map( A1 => REG_17_29_port, A2 => n810, B1 => 
                           REG_19_29_port, B2 => n792, ZN => n680);
   U1455 : AOI22_X1 port map( A1 => REG_20_29_port, A2 => n846, B1 => 
                           REG_22_29_port, B2 => n828, ZN => n679);
   U1456 : AOI22_X1 port map( A1 => REG_16_29_port, A2 => n882, B1 => 
                           REG_18_29_port, B2 => n864, ZN => n678);
   U1457 : AND4_X1 port map( A1 => n681, A2 => n680, A3 => n679, A4 => n678, ZN
                           => n698);
   U1458 : AOI22_X1 port map( A1 => REG_29_29_port, A2 => n774, B1 => 
                           REG_31_29_port, B2 => n756, ZN => n685);
   U1459 : AOI22_X1 port map( A1 => REG_25_29_port, A2 => n810, B1 => 
                           REG_27_29_port, B2 => n792, ZN => n684);
   U1460 : AOI22_X1 port map( A1 => REG_28_29_port, A2 => n846, B1 => 
                           REG_30_29_port, B2 => n828, ZN => n683);
   U1461 : AOI22_X1 port map( A1 => REG_24_29_port, A2 => n882, B1 => 
                           REG_26_29_port, B2 => n864, ZN => n682);
   U1462 : AND4_X1 port map( A1 => n685, A2 => n684, A3 => n683, A4 => n682, ZN
                           => n697);
   U1463 : AOI22_X1 port map( A1 => REG_5_29_port, A2 => n774, B1 => 
                           REG_7_29_port, B2 => n756, ZN => n689);
   U1464 : AOI22_X1 port map( A1 => REG_1_29_port, A2 => n810, B1 => 
                           REG_3_29_port, B2 => n792, ZN => n688);
   U1465 : AOI22_X1 port map( A1 => REG_4_29_port, A2 => n846, B1 => 
                           REG_6_29_port, B2 => n828, ZN => n687);
   U1466 : AOI22_X1 port map( A1 => REG_0_29_port, A2 => n882, B1 => 
                           REG_2_29_port, B2 => n864, ZN => n686);
   U1467 : NAND4_X1 port map( A1 => n689, A2 => n688, A3 => n687, A4 => n686, 
                           ZN => n695);
   U1468 : AOI22_X1 port map( A1 => REG_13_29_port, A2 => n774, B1 => 
                           REG_15_29_port, B2 => n756, ZN => n693);
   U1469 : AOI22_X1 port map( A1 => REG_9_29_port, A2 => n810, B1 => 
                           REG_11_29_port, B2 => n792, ZN => n692);
   U1470 : AOI22_X1 port map( A1 => REG_12_29_port, A2 => n846, B1 => 
                           REG_14_29_port, B2 => n828, ZN => n691);
   U1471 : AOI22_X1 port map( A1 => REG_8_29_port, A2 => n882, B1 => 
                           REG_10_29_port, B2 => n864, ZN => n690);
   U1472 : NAND4_X1 port map( A1 => n693, A2 => n692, A3 => n691, A4 => n690, 
                           ZN => n694);
   U1473 : AOI22_X1 port map( A1 => n695, A2 => n898, B1 => n694, B2 => n894, 
                           ZN => n696);
   U1474 : OAI221_X1 port map( B1 => n906, B2 => n698, C1 => n904, C2 => n697, 
                           A => n696, ZN => N254);
   U1475 : AOI22_X1 port map( A1 => REG_21_30_port, A2 => n774, B1 => 
                           REG_23_30_port, B2 => n756, ZN => n702);
   U1476 : AOI22_X1 port map( A1 => REG_17_30_port, A2 => n810, B1 => 
                           REG_19_30_port, B2 => n792, ZN => n701);
   U1477 : AOI22_X1 port map( A1 => REG_20_30_port, A2 => n846, B1 => 
                           REG_22_30_port, B2 => n828, ZN => n700);
   U1478 : AOI22_X1 port map( A1 => REG_16_30_port, A2 => n882, B1 => 
                           REG_18_30_port, B2 => n864, ZN => n699);
   U1479 : AND4_X1 port map( A1 => n702, A2 => n701, A3 => n700, A4 => n699, ZN
                           => n719);
   U1480 : AOI22_X1 port map( A1 => REG_29_30_port, A2 => n773, B1 => 
                           REG_31_30_port, B2 => n755, ZN => n706);
   U1481 : AOI22_X1 port map( A1 => REG_25_30_port, A2 => n809, B1 => 
                           REG_27_30_port, B2 => n791, ZN => n705);
   U1482 : AOI22_X1 port map( A1 => REG_28_30_port, A2 => n845, B1 => 
                           REG_30_30_port, B2 => n827, ZN => n704);
   U1483 : AOI22_X1 port map( A1 => REG_24_30_port, A2 => n881, B1 => 
                           REG_26_30_port, B2 => n863, ZN => n703);
   U1484 : AND4_X1 port map( A1 => n706, A2 => n705, A3 => n704, A4 => n703, ZN
                           => n718);
   U1485 : AOI22_X1 port map( A1 => REG_5_30_port, A2 => n773, B1 => 
                           REG_7_30_port, B2 => n755, ZN => n710);
   U1486 : AOI22_X1 port map( A1 => REG_1_30_port, A2 => n809, B1 => 
                           REG_3_30_port, B2 => n791, ZN => n709);
   U1487 : AOI22_X1 port map( A1 => REG_4_30_port, A2 => n845, B1 => 
                           REG_6_30_port, B2 => n827, ZN => n708);
   U1488 : AOI22_X1 port map( A1 => REG_0_30_port, A2 => n881, B1 => 
                           REG_2_30_port, B2 => n863, ZN => n707);
   U1489 : NAND4_X1 port map( A1 => n710, A2 => n709, A3 => n708, A4 => n707, 
                           ZN => n716);
   U1490 : AOI22_X1 port map( A1 => REG_13_30_port, A2 => n773, B1 => 
                           REG_15_30_port, B2 => n755, ZN => n714);
   U1491 : AOI22_X1 port map( A1 => REG_9_30_port, A2 => n809, B1 => 
                           REG_11_30_port, B2 => n791, ZN => n713);
   U1492 : AOI22_X1 port map( A1 => REG_12_30_port, A2 => n845, B1 => 
                           REG_14_30_port, B2 => n827, ZN => n712);
   U1493 : AOI22_X1 port map( A1 => REG_8_30_port, A2 => n881, B1 => 
                           REG_10_30_port, B2 => n863, ZN => n711);
   U1494 : NAND4_X1 port map( A1 => n714, A2 => n713, A3 => n712, A4 => n711, 
                           ZN => n715);
   U1495 : AOI22_X1 port map( A1 => n716, A2 => n898, B1 => n715, B2 => n894, 
                           ZN => n717);
   U1496 : OAI221_X1 port map( B1 => n906, B2 => n719, C1 => n904, C2 => n718, 
                           A => n717, ZN => N253);
   U1497 : AOI22_X1 port map( A1 => REG_21_31_port, A2 => n773, B1 => 
                           REG_23_31_port, B2 => n755, ZN => n723);
   U1498 : AOI22_X1 port map( A1 => REG_17_31_port, A2 => n809, B1 => 
                           REG_19_31_port, B2 => n791, ZN => n722);
   U1499 : AOI22_X1 port map( A1 => REG_20_31_port, A2 => n845, B1 => 
                           REG_22_31_port, B2 => n827, ZN => n721);
   U1500 : AOI22_X1 port map( A1 => REG_16_31_port, A2 => n881, B1 => 
                           REG_18_31_port, B2 => n863, ZN => n720);
   U1501 : AND4_X1 port map( A1 => n723, A2 => n722, A3 => n721, A4 => n720, ZN
                           => n744);
   U1502 : AOI22_X1 port map( A1 => REG_29_31_port, A2 => n773, B1 => 
                           REG_31_31_port, B2 => n755, ZN => n727);
   U1503 : AOI22_X1 port map( A1 => REG_25_31_port, A2 => n809, B1 => 
                           REG_27_31_port, B2 => n791, ZN => n726);
   U1504 : AOI22_X1 port map( A1 => REG_28_31_port, A2 => n845, B1 => 
                           REG_30_31_port, B2 => n827, ZN => n725);
   U1505 : AOI22_X1 port map( A1 => REG_24_31_port, A2 => n881, B1 => 
                           REG_26_31_port, B2 => n863, ZN => n724);
   U1506 : AND4_X1 port map( A1 => n727, A2 => n726, A3 => n725, A4 => n724, ZN
                           => n742);
   U1507 : AOI22_X1 port map( A1 => REG_5_31_port, A2 => n773, B1 => 
                           REG_7_31_port, B2 => n755, ZN => n731);
   U1508 : AOI22_X1 port map( A1 => REG_1_31_port, A2 => n809, B1 => 
                           REG_3_31_port, B2 => n791, ZN => n730);
   U1509 : AOI22_X1 port map( A1 => REG_4_31_port, A2 => n845, B1 => 
                           REG_6_31_port, B2 => n827, ZN => n729);
   U1510 : AOI22_X1 port map( A1 => REG_0_31_port, A2 => n881, B1 => 
                           REG_2_31_port, B2 => n863, ZN => n728);
   U1511 : NAND4_X1 port map( A1 => n731, A2 => n730, A3 => n729, A4 => n728, 
                           ZN => n738);
   U1512 : AOI22_X1 port map( A1 => REG_13_31_port, A2 => n773, B1 => 
                           REG_15_31_port, B2 => n755, ZN => n735);
   U1513 : AOI22_X1 port map( A1 => REG_9_31_port, A2 => n809, B1 => 
                           REG_11_31_port, B2 => n791, ZN => n734);
   U1514 : AOI22_X1 port map( A1 => REG_12_31_port, A2 => n845, B1 => 
                           REG_14_31_port, B2 => n827, ZN => n733);
   U1515 : AOI22_X1 port map( A1 => REG_8_31_port, A2 => n881, B1 => 
                           REG_10_31_port, B2 => n863, ZN => n732);
   U1516 : NAND4_X1 port map( A1 => n735, A2 => n734, A3 => n733, A4 => n732, 
                           ZN => n736);
   U1517 : AOI22_X1 port map( A1 => n898, A2 => n738, B1 => n894, B2 => n736, 
                           ZN => n740);
   U1518 : OAI221_X1 port map( B1 => n744, B2 => n906, C1 => n742, C2 => n904, 
                           A => n740, ZN => N252);
   U1519 : NOR2_X1 port map( A1 => n1590, A2 => ADD_RD2(1), ZN => n909);
   U1520 : NOR2_X1 port map( A1 => n1590, A2 => n1591, ZN => n910);
   U1521 : AOI22_X1 port map( A1 => REG_21_0_port, A2 => n4, B1 => 
                           REG_23_0_port, B2 => n2, ZN => n916);
   U1522 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n911);
   U1523 : NOR2_X1 port map( A1 => n1591, A2 => ADD_RD2(2), ZN => n912);
   U1524 : AOI22_X1 port map( A1 => REG_17_0_port, A2 => n6, B1 => 
                           REG_19_0_port, B2 => n5, ZN => n915);
   U1525 : AOI22_X1 port map( A1 => REG_20_0_port, A2 => n7, B1 => 
                           REG_22_0_port, B2 => n3, ZN => n914);
   U1526 : AOI22_X1 port map( A1 => REG_16_0_port, A2 => n9, B1 => 
                           REG_18_0_port, B2 => n8, ZN => n913);
   U1527 : AND4_X1 port map( A1 => n916, A2 => n915, A3 => n914, A4 => n913, ZN
                           => n933);
   U1528 : AOI22_X1 port map( A1 => REG_29_0_port, A2 => n4, B1 => 
                           REG_31_0_port, B2 => n2, ZN => n920);
   U1529 : AOI22_X1 port map( A1 => REG_25_0_port, A2 => n6, B1 => 
                           REG_27_0_port, B2 => n5, ZN => n919);
   U1530 : AOI22_X1 port map( A1 => REG_28_0_port, A2 => n7, B1 => 
                           REG_30_0_port, B2 => n3, ZN => n918);
   U1531 : AOI22_X1 port map( A1 => REG_24_0_port, A2 => n9, B1 => 
                           REG_26_0_port, B2 => n8, ZN => n917);
   U1532 : AND4_X1 port map( A1 => n920, A2 => n919, A3 => n918, A4 => n917, ZN
                           => n932);
   U1533 : AOI22_X1 port map( A1 => REG_5_0_port, A2 => n4, B1 => REG_7_0_port,
                           B2 => n2, ZN => n924);
   U1534 : AOI22_X1 port map( A1 => REG_1_0_port, A2 => n6, B1 => REG_3_0_port,
                           B2 => n5, ZN => n923);
   U1535 : AOI22_X1 port map( A1 => REG_4_0_port, A2 => n7, B1 => REG_6_0_port,
                           B2 => n3, ZN => n922);
   U1536 : AOI22_X1 port map( A1 => REG_0_0_port, A2 => n9, B1 => REG_2_0_port,
                           B2 => n8, ZN => n921);
   U1537 : NAND4_X1 port map( A1 => n924, A2 => n923, A3 => n922, A4 => n921, 
                           ZN => n930);
   U1538 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n1583);
   U1539 : AOI22_X1 port map( A1 => REG_13_0_port, A2 => n4, B1 => 
                           REG_15_0_port, B2 => n2, ZN => n928);
   U1540 : AOI22_X1 port map( A1 => REG_9_0_port, A2 => n6, B1 => REG_11_0_port
                           , B2 => n5, ZN => n927);
   U1541 : AOI22_X1 port map( A1 => REG_12_0_port, A2 => n7, B1 => 
                           REG_14_0_port, B2 => n3, ZN => n926);
   U1542 : AOI22_X1 port map( A1 => REG_8_0_port, A2 => n9, B1 => REG_10_0_port
                           , B2 => n8, ZN => n925);
   U1543 : NAND4_X1 port map( A1 => n928, A2 => n927, A3 => n926, A4 => n925, 
                           ZN => n929);
   U1544 : AOI22_X1 port map( A1 => n930, A2 => n1619, B1 => n929, B2 => n1581,
                           ZN => n931);
   U1545 : OAI221_X1 port map( B1 => n1587, B2 => n933, C1 => n1585, C2 => n932
                           , A => n931, ZN => N315);
   U1546 : AOI22_X1 port map( A1 => REG_21_1_port, A2 => n4, B1 => 
                           REG_23_1_port, B2 => n2, ZN => n937);
   U1547 : AOI22_X1 port map( A1 => REG_17_1_port, A2 => n6, B1 => 
                           REG_19_1_port, B2 => n5, ZN => n936);
   U1548 : AOI22_X1 port map( A1 => REG_20_1_port, A2 => n7, B1 => 
                           REG_22_1_port, B2 => n3, ZN => n935);
   U1549 : AOI22_X1 port map( A1 => REG_16_1_port, A2 => n9, B1 => 
                           REG_18_1_port, B2 => n8, ZN => n934);
   U1550 : AND4_X1 port map( A1 => n937, A2 => n936, A3 => n935, A4 => n934, ZN
                           => n954);
   U1551 : AOI22_X1 port map( A1 => REG_29_1_port, A2 => n4, B1 => 
                           REG_31_1_port, B2 => n2, ZN => n941);
   U1552 : AOI22_X1 port map( A1 => REG_25_1_port, A2 => n6, B1 => 
                           REG_27_1_port, B2 => n5, ZN => n940);
   U1553 : AOI22_X1 port map( A1 => REG_28_1_port, A2 => n7, B1 => 
                           REG_30_1_port, B2 => n3, ZN => n939);
   U1554 : AOI22_X1 port map( A1 => REG_24_1_port, A2 => n9, B1 => 
                           REG_26_1_port, B2 => n8, ZN => n938);
   U1555 : AND4_X1 port map( A1 => n941, A2 => n940, A3 => n939, A4 => n938, ZN
                           => n953);
   U1556 : AOI22_X1 port map( A1 => REG_5_1_port, A2 => n4, B1 => REG_7_1_port,
                           B2 => n2, ZN => n945);
   U1557 : AOI22_X1 port map( A1 => REG_1_1_port, A2 => n6, B1 => REG_3_1_port,
                           B2 => n5, ZN => n944);
   U1558 : AOI22_X1 port map( A1 => REG_4_1_port, A2 => n7, B1 => REG_6_1_port,
                           B2 => n3, ZN => n943);
   U1559 : AOI22_X1 port map( A1 => REG_0_1_port, A2 => n9, B1 => REG_2_1_port,
                           B2 => n8, ZN => n942);
   U1560 : NAND4_X1 port map( A1 => n945, A2 => n944, A3 => n943, A4 => n942, 
                           ZN => n951);
   U1561 : AOI22_X1 port map( A1 => REG_13_1_port, A2 => n4, B1 => 
                           REG_15_1_port, B2 => n2, ZN => n949);
   U1562 : AOI22_X1 port map( A1 => REG_9_1_port, A2 => n6, B1 => REG_11_1_port
                           , B2 => n5, ZN => n948);
   U1563 : AOI22_X1 port map( A1 => REG_12_1_port, A2 => n7, B1 => 
                           REG_14_1_port, B2 => n3, ZN => n947);
   U1564 : AOI22_X1 port map( A1 => REG_8_1_port, A2 => n9, B1 => REG_10_1_port
                           , B2 => n8, ZN => n946);
   U1565 : NAND4_X1 port map( A1 => n949, A2 => n948, A3 => n947, A4 => n946, 
                           ZN => n950);
   U1566 : AOI22_X1 port map( A1 => n951, A2 => n1619, B1 => n950, B2 => n1581,
                           ZN => n952);
   U1567 : OAI221_X1 port map( B1 => n1587, B2 => n954, C1 => n1585, C2 => n953
                           , A => n952, ZN => N314);
   U1568 : AOI22_X1 port map( A1 => REG_21_2_port, A2 => n4, B1 => 
                           REG_23_2_port, B2 => n2, ZN => n958);
   U1569 : AOI22_X1 port map( A1 => REG_17_2_port, A2 => n6, B1 => 
                           REG_19_2_port, B2 => n5, ZN => n957);
   U1570 : AOI22_X1 port map( A1 => REG_20_2_port, A2 => n7, B1 => 
                           REG_22_2_port, B2 => n3, ZN => n956);
   U1571 : AOI22_X1 port map( A1 => REG_16_2_port, A2 => n9, B1 => 
                           REG_18_2_port, B2 => n8, ZN => n955);
   U1572 : AND4_X1 port map( A1 => n958, A2 => n957, A3 => n956, A4 => n955, ZN
                           => n975);
   U1573 : AOI22_X1 port map( A1 => REG_29_2_port, A2 => n4, B1 => 
                           REG_31_2_port, B2 => n2, ZN => n962);
   U1574 : AOI22_X1 port map( A1 => REG_25_2_port, A2 => n6, B1 => 
                           REG_27_2_port, B2 => n5, ZN => n961);
   U1575 : AOI22_X1 port map( A1 => REG_28_2_port, A2 => n7, B1 => 
                           REG_30_2_port, B2 => n3, ZN => n960);
   U1576 : AOI22_X1 port map( A1 => REG_24_2_port, A2 => n9, B1 => 
                           REG_26_2_port, B2 => n8, ZN => n959);
   U1577 : AND4_X1 port map( A1 => n962, A2 => n961, A3 => n960, A4 => n959, ZN
                           => n974);
   U1578 : AOI22_X1 port map( A1 => REG_5_2_port, A2 => n4, B1 => REG_7_2_port,
                           B2 => n2, ZN => n966);
   U1579 : AOI22_X1 port map( A1 => REG_1_2_port, A2 => n6, B1 => REG_3_2_port,
                           B2 => n5, ZN => n965);
   U1580 : AOI22_X1 port map( A1 => REG_4_2_port, A2 => n7, B1 => REG_6_2_port,
                           B2 => n3, ZN => n964);
   U1581 : AOI22_X1 port map( A1 => REG_0_2_port, A2 => n9, B1 => REG_2_2_port,
                           B2 => n8, ZN => n963);
   U1582 : NAND4_X1 port map( A1 => n966, A2 => n965, A3 => n964, A4 => n963, 
                           ZN => n972);
   U1583 : AOI22_X1 port map( A1 => REG_13_2_port, A2 => n4, B1 => 
                           REG_15_2_port, B2 => n2, ZN => n970);
   U1584 : AOI22_X1 port map( A1 => REG_9_2_port, A2 => n6, B1 => REG_11_2_port
                           , B2 => n5, ZN => n969);
   U1585 : AOI22_X1 port map( A1 => REG_12_2_port, A2 => n7, B1 => 
                           REG_14_2_port, B2 => n3, ZN => n968);
   U1586 : AOI22_X1 port map( A1 => REG_8_2_port, A2 => n9, B1 => REG_10_2_port
                           , B2 => n8, ZN => n967);
   U1587 : NAND4_X1 port map( A1 => n970, A2 => n969, A3 => n968, A4 => n967, 
                           ZN => n971);
   U1588 : AOI22_X1 port map( A1 => n972, A2 => n1619, B1 => n971, B2 => n1581,
                           ZN => n973);
   U1589 : OAI221_X1 port map( B1 => n1587, B2 => n975, C1 => n1585, C2 => n974
                           , A => n973, ZN => N313);
   U1590 : AOI22_X1 port map( A1 => REG_21_3_port, A2 => n4, B1 => 
                           REG_23_3_port, B2 => n2, ZN => n979);
   U1591 : AOI22_X1 port map( A1 => REG_17_3_port, A2 => n6, B1 => 
                           REG_19_3_port, B2 => n5, ZN => n978);
   U1592 : AOI22_X1 port map( A1 => REG_20_3_port, A2 => n7, B1 => 
                           REG_22_3_port, B2 => n3, ZN => n977);
   U1593 : AOI22_X1 port map( A1 => REG_16_3_port, A2 => n9, B1 => 
                           REG_18_3_port, B2 => n8, ZN => n976);
   U1594 : AND4_X1 port map( A1 => n979, A2 => n978, A3 => n977, A4 => n976, ZN
                           => n996);
   U1595 : AOI22_X1 port map( A1 => REG_29_3_port, A2 => n4, B1 => 
                           REG_31_3_port, B2 => n2, ZN => n983);
   U1596 : AOI22_X1 port map( A1 => REG_25_3_port, A2 => n6, B1 => 
                           REG_27_3_port, B2 => n5, ZN => n982);
   U1597 : AOI22_X1 port map( A1 => REG_28_3_port, A2 => n7, B1 => 
                           REG_30_3_port, B2 => n3, ZN => n981);
   U1598 : AOI22_X1 port map( A1 => REG_24_3_port, A2 => n9, B1 => 
                           REG_26_3_port, B2 => n8, ZN => n980);
   U1599 : AND4_X1 port map( A1 => n983, A2 => n982, A3 => n981, A4 => n980, ZN
                           => n995);
   U1600 : AOI22_X1 port map( A1 => REG_5_3_port, A2 => n4, B1 => REG_7_3_port,
                           B2 => n2, ZN => n987);
   U1601 : AOI22_X1 port map( A1 => REG_1_3_port, A2 => n6, B1 => REG_3_3_port,
                           B2 => n5, ZN => n986);
   U1602 : AOI22_X1 port map( A1 => REG_4_3_port, A2 => n7, B1 => REG_6_3_port,
                           B2 => n3, ZN => n985);
   U1603 : AOI22_X1 port map( A1 => REG_0_3_port, A2 => n9, B1 => REG_2_3_port,
                           B2 => n8, ZN => n984);
   U1604 : NAND4_X1 port map( A1 => n987, A2 => n986, A3 => n985, A4 => n984, 
                           ZN => n993);
   U1605 : AOI22_X1 port map( A1 => REG_13_3_port, A2 => n4, B1 => 
                           REG_15_3_port, B2 => n2, ZN => n991);
   U1606 : AOI22_X1 port map( A1 => REG_9_3_port, A2 => n6, B1 => REG_11_3_port
                           , B2 => n5, ZN => n990);
   U1607 : AOI22_X1 port map( A1 => REG_12_3_port, A2 => n7, B1 => 
                           REG_14_3_port, B2 => n3, ZN => n989);
   U1608 : AOI22_X1 port map( A1 => REG_8_3_port, A2 => n9, B1 => REG_10_3_port
                           , B2 => n8, ZN => n988);
   U1609 : NAND4_X1 port map( A1 => n991, A2 => n990, A3 => n989, A4 => n988, 
                           ZN => n992);
   U1610 : AOI22_X1 port map( A1 => n993, A2 => n1619, B1 => n992, B2 => n1581,
                           ZN => n994);
   U1611 : OAI221_X1 port map( B1 => n1587, B2 => n996, C1 => n1585, C2 => n995
                           , A => n994, ZN => N312);
   U1612 : AOI22_X1 port map( A1 => REG_21_4_port, A2 => n4, B1 => 
                           REG_23_4_port, B2 => n2, ZN => n1000);
   U1613 : AOI22_X1 port map( A1 => REG_17_4_port, A2 => n6, B1 => 
                           REG_19_4_port, B2 => n5, ZN => n999);
   U1614 : AOI22_X1 port map( A1 => REG_20_4_port, A2 => n7, B1 => 
                           REG_22_4_port, B2 => n3, ZN => n998);
   U1615 : AOI22_X1 port map( A1 => REG_16_4_port, A2 => n9, B1 => 
                           REG_18_4_port, B2 => n8, ZN => n997);
   U1616 : AND4_X1 port map( A1 => n1000, A2 => n999, A3 => n998, A4 => n997, 
                           ZN => n1017);
   U1617 : AOI22_X1 port map( A1 => REG_29_4_port, A2 => n4, B1 => 
                           REG_31_4_port, B2 => n2, ZN => n1004);
   U1618 : AOI22_X1 port map( A1 => REG_25_4_port, A2 => n6, B1 => 
                           REG_27_4_port, B2 => n5, ZN => n1003);
   U1619 : AOI22_X1 port map( A1 => REG_28_4_port, A2 => n7, B1 => 
                           REG_30_4_port, B2 => n3, ZN => n1002);
   U1620 : AOI22_X1 port map( A1 => REG_24_4_port, A2 => n9, B1 => 
                           REG_26_4_port, B2 => n8, ZN => n1001);
   U1621 : AND4_X1 port map( A1 => n1004, A2 => n1003, A3 => n1002, A4 => n1001
                           , ZN => n1016);
   U1622 : AOI22_X1 port map( A1 => REG_5_4_port, A2 => n4, B1 => REG_7_4_port,
                           B2 => n2, ZN => n1008);
   U1623 : AOI22_X1 port map( A1 => REG_1_4_port, A2 => n6, B1 => REG_3_4_port,
                           B2 => n5, ZN => n1007);
   U1624 : AOI22_X1 port map( A1 => REG_4_4_port, A2 => n7, B1 => REG_6_4_port,
                           B2 => n3, ZN => n1006);
   U1625 : AOI22_X1 port map( A1 => REG_0_4_port, A2 => n9, B1 => REG_2_4_port,
                           B2 => n8, ZN => n1005);
   U1626 : NAND4_X1 port map( A1 => n1008, A2 => n1007, A3 => n1006, A4 => 
                           n1005, ZN => n1014);
   U1627 : AOI22_X1 port map( A1 => REG_13_4_port, A2 => n4, B1 => 
                           REG_15_4_port, B2 => n2, ZN => n1012);
   U1628 : AOI22_X1 port map( A1 => REG_9_4_port, A2 => n6, B1 => REG_11_4_port
                           , B2 => n5, ZN => n1011);
   U1629 : AOI22_X1 port map( A1 => REG_12_4_port, A2 => n7, B1 => 
                           REG_14_4_port, B2 => n3, ZN => n1010);
   U1630 : AOI22_X1 port map( A1 => REG_8_4_port, A2 => n9, B1 => REG_10_4_port
                           , B2 => n8, ZN => n1009);
   U1631 : NAND4_X1 port map( A1 => n1012, A2 => n1011, A3 => n1010, A4 => 
                           n1009, ZN => n1013);
   U1632 : AOI22_X1 port map( A1 => n1014, A2 => n1619, B1 => n1013, B2 => 
                           n1581, ZN => n1015);
   U1633 : OAI221_X1 port map( B1 => n1587, B2 => n1017, C1 => n1585, C2 => 
                           n1016, A => n1015, ZN => N311);
   U1634 : AOI22_X1 port map( A1 => REG_21_5_port, A2 => n4, B1 => 
                           REG_23_5_port, B2 => n2, ZN => n1021);
   U1635 : AOI22_X1 port map( A1 => REG_17_5_port, A2 => n6, B1 => 
                           REG_19_5_port, B2 => n5, ZN => n1020);
   U1636 : AOI22_X1 port map( A1 => REG_20_5_port, A2 => n7, B1 => 
                           REG_22_5_port, B2 => n3, ZN => n1019);
   U1637 : AOI22_X1 port map( A1 => REG_16_5_port, A2 => n9, B1 => 
                           REG_18_5_port, B2 => n8, ZN => n1018);
   U1638 : AND4_X1 port map( A1 => n1021, A2 => n1020, A3 => n1019, A4 => n1018
                           , ZN => n1038);
   U1639 : AOI22_X1 port map( A1 => REG_29_5_port, A2 => n4, B1 => 
                           REG_31_5_port, B2 => n2, ZN => n1025);
   U1640 : AOI22_X1 port map( A1 => REG_25_5_port, A2 => n6, B1 => 
                           REG_27_5_port, B2 => n5, ZN => n1024);
   U1641 : AOI22_X1 port map( A1 => REG_28_5_port, A2 => n7, B1 => 
                           REG_30_5_port, B2 => n3, ZN => n1023);
   U1642 : AOI22_X1 port map( A1 => REG_24_5_port, A2 => n9, B1 => 
                           REG_26_5_port, B2 => n8, ZN => n1022);
   U1643 : AND4_X1 port map( A1 => n1025, A2 => n1024, A3 => n1023, A4 => n1022
                           , ZN => n1037);
   U1644 : AOI22_X1 port map( A1 => REG_5_5_port, A2 => n4, B1 => REG_7_5_port,
                           B2 => n2, ZN => n1029);
   U1645 : AOI22_X1 port map( A1 => REG_1_5_port, A2 => n6, B1 => REG_3_5_port,
                           B2 => n5, ZN => n1028);
   U1646 : AOI22_X1 port map( A1 => REG_4_5_port, A2 => n7, B1 => REG_6_5_port,
                           B2 => n3, ZN => n1027);
   U1647 : AOI22_X1 port map( A1 => REG_0_5_port, A2 => n9, B1 => REG_2_5_port,
                           B2 => n8, ZN => n1026);
   U1648 : NAND4_X1 port map( A1 => n1029, A2 => n1028, A3 => n1027, A4 => 
                           n1026, ZN => n1035);
   U1649 : AOI22_X1 port map( A1 => REG_13_5_port, A2 => n4, B1 => 
                           REG_15_5_port, B2 => n2, ZN => n1033);
   U1650 : AOI22_X1 port map( A1 => REG_9_5_port, A2 => n6, B1 => REG_11_5_port
                           , B2 => n5, ZN => n1032);
   U1651 : AOI22_X1 port map( A1 => REG_12_5_port, A2 => n7, B1 => 
                           REG_14_5_port, B2 => n3, ZN => n1031);
   U1652 : AOI22_X1 port map( A1 => REG_8_5_port, A2 => n9, B1 => REG_10_5_port
                           , B2 => n8, ZN => n1030);
   U1653 : NAND4_X1 port map( A1 => n1033, A2 => n1032, A3 => n1031, A4 => 
                           n1030, ZN => n1034);
   U1654 : AOI22_X1 port map( A1 => n1035, A2 => n1619, B1 => n1034, B2 => 
                           n1581, ZN => n1036);
   U1655 : OAI221_X1 port map( B1 => n1587, B2 => n1038, C1 => n1585, C2 => 
                           n1037, A => n1036, ZN => N310);
   U1656 : AOI22_X1 port map( A1 => REG_21_6_port, A2 => n4, B1 => 
                           REG_23_6_port, B2 => n2, ZN => n1042);
   U1657 : AOI22_X1 port map( A1 => REG_17_6_port, A2 => n6, B1 => 
                           REG_19_6_port, B2 => n5, ZN => n1041);
   U1658 : AOI22_X1 port map( A1 => REG_20_6_port, A2 => n7, B1 => 
                           REG_22_6_port, B2 => n3, ZN => n1040);
   U1659 : AOI22_X1 port map( A1 => REG_16_6_port, A2 => n9, B1 => 
                           REG_18_6_port, B2 => n8, ZN => n1039);
   U1660 : AND4_X1 port map( A1 => n1042, A2 => n1041, A3 => n1040, A4 => n1039
                           , ZN => n1059);
   U1661 : AOI22_X1 port map( A1 => REG_29_6_port, A2 => n4, B1 => 
                           REG_31_6_port, B2 => n2, ZN => n1046);
   U1662 : AOI22_X1 port map( A1 => REG_25_6_port, A2 => n6, B1 => 
                           REG_27_6_port, B2 => n5, ZN => n1045);
   U1663 : AOI22_X1 port map( A1 => REG_28_6_port, A2 => n7, B1 => 
                           REG_30_6_port, B2 => n3, ZN => n1044);
   U1664 : AOI22_X1 port map( A1 => REG_24_6_port, A2 => n9, B1 => 
                           REG_26_6_port, B2 => n8, ZN => n1043);
   U1665 : AND4_X1 port map( A1 => n1046, A2 => n1045, A3 => n1044, A4 => n1043
                           , ZN => n1058);
   U1666 : AOI22_X1 port map( A1 => REG_5_6_port, A2 => n4, B1 => REG_7_6_port,
                           B2 => n2, ZN => n1050);
   U1667 : AOI22_X1 port map( A1 => REG_1_6_port, A2 => n6, B1 => REG_3_6_port,
                           B2 => n5, ZN => n1049);
   U1668 : AOI22_X1 port map( A1 => REG_4_6_port, A2 => n7, B1 => REG_6_6_port,
                           B2 => n3, ZN => n1048);
   U1669 : AOI22_X1 port map( A1 => REG_0_6_port, A2 => n9, B1 => REG_2_6_port,
                           B2 => n8, ZN => n1047);
   U1670 : NAND4_X1 port map( A1 => n1050, A2 => n1049, A3 => n1048, A4 => 
                           n1047, ZN => n1056);
   U1671 : AOI22_X1 port map( A1 => REG_13_6_port, A2 => n4, B1 => 
                           REG_15_6_port, B2 => n2, ZN => n1054);
   U1672 : AOI22_X1 port map( A1 => REG_9_6_port, A2 => n6, B1 => REG_11_6_port
                           , B2 => n5, ZN => n1053);
   U1673 : AOI22_X1 port map( A1 => REG_12_6_port, A2 => n7, B1 => 
                           REG_14_6_port, B2 => n3, ZN => n1052);
   U1674 : AOI22_X1 port map( A1 => REG_8_6_port, A2 => n9, B1 => REG_10_6_port
                           , B2 => n8, ZN => n1051);
   U1675 : NAND4_X1 port map( A1 => n1054, A2 => n1053, A3 => n1052, A4 => 
                           n1051, ZN => n1055);
   U1676 : AOI22_X1 port map( A1 => n1056, A2 => n1619, B1 => n1055, B2 => 
                           n1581, ZN => n1057);
   U1677 : OAI221_X1 port map( B1 => n1587, B2 => n1059, C1 => n1585, C2 => 
                           n1058, A => n1057, ZN => N309);
   U1678 : AOI22_X1 port map( A1 => REG_21_7_port, A2 => n4, B1 => 
                           REG_23_7_port, B2 => n2, ZN => n1063);
   U1679 : AOI22_X1 port map( A1 => REG_17_7_port, A2 => n6, B1 => 
                           REG_19_7_port, B2 => n5, ZN => n1062);
   U1680 : AOI22_X1 port map( A1 => REG_20_7_port, A2 => n7, B1 => 
                           REG_22_7_port, B2 => n3, ZN => n1061);
   U1681 : AOI22_X1 port map( A1 => REG_16_7_port, A2 => n9, B1 => 
                           REG_18_7_port, B2 => n8, ZN => n1060);
   U1682 : AND4_X1 port map( A1 => n1063, A2 => n1062, A3 => n1061, A4 => n1060
                           , ZN => n1080);
   U1683 : AOI22_X1 port map( A1 => REG_29_7_port, A2 => n4, B1 => 
                           REG_31_7_port, B2 => n2, ZN => n1067);
   U1684 : AOI22_X1 port map( A1 => REG_25_7_port, A2 => n6, B1 => 
                           REG_27_7_port, B2 => n5, ZN => n1066);
   U1685 : AOI22_X1 port map( A1 => REG_28_7_port, A2 => n7, B1 => 
                           REG_30_7_port, B2 => n3, ZN => n1065);
   U1686 : AOI22_X1 port map( A1 => REG_24_7_port, A2 => n9, B1 => 
                           REG_26_7_port, B2 => n8, ZN => n1064);
   U1687 : AND4_X1 port map( A1 => n1067, A2 => n1066, A3 => n1065, A4 => n1064
                           , ZN => n1079);
   U1688 : AOI22_X1 port map( A1 => REG_5_7_port, A2 => n4, B1 => REG_7_7_port,
                           B2 => n2, ZN => n1071);
   U1689 : AOI22_X1 port map( A1 => REG_1_7_port, A2 => n6, B1 => REG_3_7_port,
                           B2 => n5, ZN => n1070);
   U1690 : AOI22_X1 port map( A1 => REG_4_7_port, A2 => n7, B1 => REG_6_7_port,
                           B2 => n3, ZN => n1069);
   U1691 : AOI22_X1 port map( A1 => REG_0_7_port, A2 => n9, B1 => REG_2_7_port,
                           B2 => n8, ZN => n1068);
   U1692 : NAND4_X1 port map( A1 => n1071, A2 => n1070, A3 => n1069, A4 => 
                           n1068, ZN => n1077);
   U1693 : AOI22_X1 port map( A1 => REG_13_7_port, A2 => n4, B1 => 
                           REG_15_7_port, B2 => n2, ZN => n1075);
   U1694 : AOI22_X1 port map( A1 => REG_9_7_port, A2 => n6, B1 => REG_11_7_port
                           , B2 => n5, ZN => n1074);
   U1695 : AOI22_X1 port map( A1 => REG_12_7_port, A2 => n7, B1 => 
                           REG_14_7_port, B2 => n3, ZN => n1073);
   U1696 : AOI22_X1 port map( A1 => REG_8_7_port, A2 => n9, B1 => REG_10_7_port
                           , B2 => n8, ZN => n1072);
   U1697 : NAND4_X1 port map( A1 => n1075, A2 => n1074, A3 => n1073, A4 => 
                           n1072, ZN => n1076);
   U1698 : AOI22_X1 port map( A1 => n1077, A2 => n1619, B1 => n1076, B2 => 
                           n1581, ZN => n1078);
   U1699 : OAI221_X1 port map( B1 => n1587, B2 => n1080, C1 => n1585, C2 => 
                           n1079, A => n1078, ZN => N308);
   U1700 : AOI22_X1 port map( A1 => REG_21_8_port, A2 => n4, B1 => 
                           REG_23_8_port, B2 => n2, ZN => n1084);
   U1701 : AOI22_X1 port map( A1 => REG_17_8_port, A2 => n6, B1 => 
                           REG_19_8_port, B2 => n5, ZN => n1083);
   U1702 : AOI22_X1 port map( A1 => REG_20_8_port, A2 => n7, B1 => 
                           REG_22_8_port, B2 => n3, ZN => n1082);
   U1703 : AOI22_X1 port map( A1 => REG_16_8_port, A2 => n9, B1 => 
                           REG_18_8_port, B2 => n8, ZN => n1081);
   U1704 : AND4_X1 port map( A1 => n1084, A2 => n1083, A3 => n1082, A4 => n1081
                           , ZN => n1101);
   U1705 : AOI22_X1 port map( A1 => REG_29_8_port, A2 => n4, B1 => 
                           REG_31_8_port, B2 => n2, ZN => n1088);
   U1706 : AOI22_X1 port map( A1 => REG_25_8_port, A2 => n6, B1 => 
                           REG_27_8_port, B2 => n1600, ZN => n1087);
   U1707 : AOI22_X1 port map( A1 => REG_28_8_port, A2 => n7, B1 => 
                           REG_30_8_port, B2 => n3, ZN => n1086);
   U1708 : AOI22_X1 port map( A1 => REG_24_8_port, A2 => n9, B1 => 
                           REG_26_8_port, B2 => n8, ZN => n1085);
   U1709 : AND4_X1 port map( A1 => n1088, A2 => n1087, A3 => n1086, A4 => n1085
                           , ZN => n1100);
   U1710 : AOI22_X1 port map( A1 => REG_5_8_port, A2 => n4, B1 => REG_7_8_port,
                           B2 => n2, ZN => n1092);
   U1711 : AOI22_X1 port map( A1 => REG_1_8_port, A2 => n6, B1 => REG_3_8_port,
                           B2 => n1600, ZN => n1091);
   U1712 : AOI22_X1 port map( A1 => REG_4_8_port, A2 => n7, B1 => REG_6_8_port,
                           B2 => n3, ZN => n1090);
   U1713 : AOI22_X1 port map( A1 => REG_0_8_port, A2 => n9, B1 => REG_2_8_port,
                           B2 => n8, ZN => n1089);
   U1714 : NAND4_X1 port map( A1 => n1092, A2 => n1091, A3 => n1090, A4 => 
                           n1089, ZN => n1098);
   U1715 : AOI22_X1 port map( A1 => REG_13_8_port, A2 => n4, B1 => 
                           REG_15_8_port, B2 => n2, ZN => n1096);
   U1716 : AOI22_X1 port map( A1 => REG_9_8_port, A2 => n6, B1 => REG_11_8_port
                           , B2 => n1600, ZN => n1095);
   U1717 : AOI22_X1 port map( A1 => REG_12_8_port, A2 => n7, B1 => 
                           REG_14_8_port, B2 => n3, ZN => n1094);
   U1718 : AOI22_X1 port map( A1 => REG_8_8_port, A2 => n9, B1 => REG_10_8_port
                           , B2 => n8, ZN => n1093);
   U1719 : NAND4_X1 port map( A1 => n1096, A2 => n1095, A3 => n1094, A4 => 
                           n1093, ZN => n1097);
   U1720 : AOI22_X1 port map( A1 => n1098, A2 => n1619, B1 => n1097, B2 => 
                           n1581, ZN => n1099);
   U1721 : OAI221_X1 port map( B1 => n1587, B2 => n1101, C1 => n1585, C2 => 
                           n1100, A => n1099, ZN => N307);
   U1722 : AOI22_X1 port map( A1 => REG_21_9_port, A2 => n4, B1 => 
                           REG_23_9_port, B2 => n2, ZN => n1105);
   U1723 : AOI22_X1 port map( A1 => REG_17_9_port, A2 => n6, B1 => 
                           REG_19_9_port, B2 => n1600, ZN => n1104);
   U1724 : AOI22_X1 port map( A1 => REG_20_9_port, A2 => n7, B1 => 
                           REG_22_9_port, B2 => n3, ZN => n1103);
   U1725 : AOI22_X1 port map( A1 => REG_16_9_port, A2 => n9, B1 => 
                           REG_18_9_port, B2 => n8, ZN => n1102);
   U1726 : AND4_X1 port map( A1 => n1105, A2 => n1104, A3 => n1103, A4 => n1102
                           , ZN => n1122);
   U1727 : AOI22_X1 port map( A1 => REG_29_9_port, A2 => n4, B1 => 
                           REG_31_9_port, B2 => n2, ZN => n1109);
   U1728 : AOI22_X1 port map( A1 => REG_25_9_port, A2 => n6, B1 => 
                           REG_27_9_port, B2 => n1600, ZN => n1108);
   U1729 : AOI22_X1 port map( A1 => REG_28_9_port, A2 => n7, B1 => 
                           REG_30_9_port, B2 => n3, ZN => n1107);
   U1730 : AOI22_X1 port map( A1 => REG_24_9_port, A2 => n9, B1 => 
                           REG_26_9_port, B2 => n8, ZN => n1106);
   U1731 : AND4_X1 port map( A1 => n1109, A2 => n1108, A3 => n1107, A4 => n1106
                           , ZN => n1121);
   U1732 : AOI22_X1 port map( A1 => REG_5_9_port, A2 => n4, B1 => REG_7_9_port,
                           B2 => n2, ZN => n1113);
   U1733 : AOI22_X1 port map( A1 => REG_1_9_port, A2 => n6, B1 => REG_3_9_port,
                           B2 => n1600, ZN => n1112);
   U1734 : AOI22_X1 port map( A1 => REG_4_9_port, A2 => n7, B1 => REG_6_9_port,
                           B2 => n3, ZN => n1111);
   U1735 : AOI22_X1 port map( A1 => REG_0_9_port, A2 => n9, B1 => REG_2_9_port,
                           B2 => n8, ZN => n1110);
   U1736 : NAND4_X1 port map( A1 => n1113, A2 => n1112, A3 => n1111, A4 => 
                           n1110, ZN => n1119);
   U1737 : AOI22_X1 port map( A1 => REG_13_9_port, A2 => n4, B1 => 
                           REG_15_9_port, B2 => n2, ZN => n1117);
   U1738 : AOI22_X1 port map( A1 => REG_9_9_port, A2 => n6, B1 => REG_11_9_port
                           , B2 => n1600, ZN => n1116);
   U1739 : AOI22_X1 port map( A1 => REG_12_9_port, A2 => n7, B1 => 
                           REG_14_9_port, B2 => n3, ZN => n1115);
   U1740 : AOI22_X1 port map( A1 => REG_8_9_port, A2 => n9, B1 => REG_10_9_port
                           , B2 => n8, ZN => n1114);
   U1741 : NAND4_X1 port map( A1 => n1117, A2 => n1116, A3 => n1115, A4 => 
                           n1114, ZN => n1118);
   U1742 : AOI22_X1 port map( A1 => n1119, A2 => n1619, B1 => n1118, B2 => 
                           n1581, ZN => n1120);
   U1743 : OAI221_X1 port map( B1 => n1587, B2 => n1122, C1 => n1585, C2 => 
                           n1121, A => n1120, ZN => N306);
   U1744 : AOI22_X1 port map( A1 => REG_21_10_port, A2 => n4, B1 => 
                           REG_23_10_port, B2 => n2, ZN => n1126);
   U1745 : AOI22_X1 port map( A1 => REG_17_10_port, A2 => n6, B1 => 
                           REG_19_10_port, B2 => n1600, ZN => n1125);
   U1746 : AOI22_X1 port map( A1 => REG_20_10_port, A2 => n7, B1 => 
                           REG_22_10_port, B2 => n3, ZN => n1124);
   U1747 : AOI22_X1 port map( A1 => REG_16_10_port, A2 => n9, B1 => 
                           REG_18_10_port, B2 => n8, ZN => n1123);
   U1748 : AND4_X1 port map( A1 => n1126, A2 => n1125, A3 => n1124, A4 => n1123
                           , ZN => n1143);
   U1749 : AOI22_X1 port map( A1 => REG_29_10_port, A2 => n4, B1 => 
                           REG_31_10_port, B2 => n2, ZN => n1130);
   U1750 : AOI22_X1 port map( A1 => REG_25_10_port, A2 => n6, B1 => 
                           REG_27_10_port, B2 => n1600, ZN => n1129);
   U1751 : AOI22_X1 port map( A1 => REG_28_10_port, A2 => n7, B1 => 
                           REG_30_10_port, B2 => n3, ZN => n1128);
   U1752 : AOI22_X1 port map( A1 => REG_24_10_port, A2 => n9, B1 => 
                           REG_26_10_port, B2 => n8, ZN => n1127);
   U1753 : AND4_X1 port map( A1 => n1130, A2 => n1129, A3 => n1128, A4 => n1127
                           , ZN => n1142);
   U1754 : AOI22_X1 port map( A1 => REG_5_10_port, A2 => n4, B1 => 
                           REG_7_10_port, B2 => n2, ZN => n1134);
   U1755 : AOI22_X1 port map( A1 => REG_1_10_port, A2 => n6, B1 => 
                           REG_3_10_port, B2 => n1600, ZN => n1133);
   U1756 : AOI22_X1 port map( A1 => REG_4_10_port, A2 => n7, B1 => 
                           REG_6_10_port, B2 => n3, ZN => n1132);
   U1757 : AOI22_X1 port map( A1 => REG_0_10_port, A2 => n9, B1 => 
                           REG_2_10_port, B2 => n8, ZN => n1131);
   U1758 : NAND4_X1 port map( A1 => n1134, A2 => n1133, A3 => n1132, A4 => 
                           n1131, ZN => n1140);
   U1759 : AOI22_X1 port map( A1 => REG_13_10_port, A2 => n4, B1 => 
                           REG_15_10_port, B2 => n2, ZN => n1138);
   U1760 : AOI22_X1 port map( A1 => REG_9_10_port, A2 => n6, B1 => 
                           REG_11_10_port, B2 => n1600, ZN => n1137);
   U1761 : AOI22_X1 port map( A1 => REG_12_10_port, A2 => n7, B1 => 
                           REG_14_10_port, B2 => n3, ZN => n1136);
   U1762 : AOI22_X1 port map( A1 => REG_8_10_port, A2 => n9, B1 => 
                           REG_10_10_port, B2 => n8, ZN => n1135);
   U1763 : NAND4_X1 port map( A1 => n1138, A2 => n1137, A3 => n1136, A4 => 
                           n1135, ZN => n1139);
   U1764 : AOI22_X1 port map( A1 => n1140, A2 => n1619, B1 => n1139, B2 => 
                           n1581, ZN => n1141);
   U1765 : OAI221_X1 port map( B1 => n1587, B2 => n1143, C1 => n1585, C2 => 
                           n1142, A => n1141, ZN => N305);
   U1766 : AOI22_X1 port map( A1 => REG_21_11_port, A2 => n4, B1 => 
                           REG_23_11_port, B2 => n1597, ZN => n1147);
   U1767 : AOI22_X1 port map( A1 => REG_17_11_port, A2 => n1604, B1 => 
                           REG_19_11_port, B2 => n5, ZN => n1146);
   U1768 : AOI22_X1 port map( A1 => REG_20_11_port, A2 => n7, B1 => 
                           REG_22_11_port, B2 => n1609, ZN => n1145);
   U1769 : AOI22_X1 port map( A1 => REG_16_11_port, A2 => n1617, B1 => 
                           REG_18_11_port, B2 => n8, ZN => n1144);
   U1770 : AND4_X1 port map( A1 => n1147, A2 => n1146, A3 => n1145, A4 => n1144
                           , ZN => n1164);
   U1771 : AOI22_X1 port map( A1 => REG_29_11_port, A2 => n4, B1 => 
                           REG_31_11_port, B2 => n1597, ZN => n1151);
   U1772 : AOI22_X1 port map( A1 => REG_25_11_port, A2 => n1604, B1 => 
                           REG_27_11_port, B2 => n5, ZN => n1150);
   U1773 : AOI22_X1 port map( A1 => REG_28_11_port, A2 => n7, B1 => 
                           REG_30_11_port, B2 => n1609, ZN => n1149);
   U1774 : AOI22_X1 port map( A1 => REG_24_11_port, A2 => n1617, B1 => 
                           REG_26_11_port, B2 => n8, ZN => n1148);
   U1775 : AND4_X1 port map( A1 => n1151, A2 => n1150, A3 => n1149, A4 => n1148
                           , ZN => n1163);
   U1776 : AOI22_X1 port map( A1 => REG_5_11_port, A2 => n4, B1 => 
                           REG_7_11_port, B2 => n1597, ZN => n1155);
   U1777 : AOI22_X1 port map( A1 => REG_1_11_port, A2 => n1604, B1 => 
                           REG_3_11_port, B2 => n5, ZN => n1154);
   U1778 : AOI22_X1 port map( A1 => REG_4_11_port, A2 => n7, B1 => 
                           REG_6_11_port, B2 => n1609, ZN => n1153);
   U1779 : AOI22_X1 port map( A1 => REG_0_11_port, A2 => n1617, B1 => 
                           REG_2_11_port, B2 => n8, ZN => n1152);
   U1780 : NAND4_X1 port map( A1 => n1155, A2 => n1154, A3 => n1153, A4 => 
                           n1152, ZN => n1161);
   U1781 : AOI22_X1 port map( A1 => REG_13_11_port, A2 => n4, B1 => 
                           REG_15_11_port, B2 => n1597, ZN => n1159);
   U1782 : AOI22_X1 port map( A1 => REG_9_11_port, A2 => n1604, B1 => 
                           REG_11_11_port, B2 => n5, ZN => n1158);
   U1783 : AOI22_X1 port map( A1 => REG_12_11_port, A2 => n7, B1 => 
                           REG_14_11_port, B2 => n1609, ZN => n1157);
   U1784 : AOI22_X1 port map( A1 => REG_8_11_port, A2 => n1617, B1 => 
                           REG_10_11_port, B2 => n8, ZN => n1156);
   U1785 : NAND4_X1 port map( A1 => n1159, A2 => n1158, A3 => n1157, A4 => 
                           n1156, ZN => n1160);
   U1786 : AOI22_X1 port map( A1 => n1161, A2 => n1619, B1 => n1160, B2 => 
                           n1618, ZN => n1162);
   U1787 : OAI221_X1 port map( B1 => n1587, B2 => n1164, C1 => n1585, C2 => 
                           n1163, A => n1162, ZN => N304);
   U1788 : AOI22_X1 port map( A1 => REG_21_12_port, A2 => n4, B1 => 
                           REG_23_12_port, B2 => n1597, ZN => n1168);
   U1789 : AOI22_X1 port map( A1 => REG_17_12_port, A2 => n1604, B1 => 
                           REG_19_12_port, B2 => n5, ZN => n1167);
   U1790 : AOI22_X1 port map( A1 => REG_20_12_port, A2 => n7, B1 => 
                           REG_22_12_port, B2 => n1609, ZN => n1166);
   U1791 : AOI22_X1 port map( A1 => REG_16_12_port, A2 => n1617, B1 => 
                           REG_18_12_port, B2 => n8, ZN => n1165);
   U1792 : AND4_X1 port map( A1 => n1168, A2 => n1167, A3 => n1166, A4 => n1165
                           , ZN => n1185);
   U1793 : AOI22_X1 port map( A1 => REG_29_12_port, A2 => n4, B1 => 
                           REG_31_12_port, B2 => n1597, ZN => n1172);
   U1794 : AOI22_X1 port map( A1 => REG_25_12_port, A2 => n1604, B1 => 
                           REG_27_12_port, B2 => n5, ZN => n1171);
   U1795 : AOI22_X1 port map( A1 => REG_28_12_port, A2 => n7, B1 => 
                           REG_30_12_port, B2 => n1609, ZN => n1170);
   U1796 : AOI22_X1 port map( A1 => REG_24_12_port, A2 => n1617, B1 => 
                           REG_26_12_port, B2 => n8, ZN => n1169);
   U1797 : AND4_X1 port map( A1 => n1172, A2 => n1171, A3 => n1170, A4 => n1169
                           , ZN => n1184);
   U1798 : AOI22_X1 port map( A1 => REG_5_12_port, A2 => n4, B1 => 
                           REG_7_12_port, B2 => n1597, ZN => n1176);
   U1799 : AOI22_X1 port map( A1 => REG_1_12_port, A2 => n1604, B1 => 
                           REG_3_12_port, B2 => n5, ZN => n1175);
   U1800 : AOI22_X1 port map( A1 => REG_4_12_port, A2 => n7, B1 => 
                           REG_6_12_port, B2 => n1609, ZN => n1174);
   U1801 : AOI22_X1 port map( A1 => REG_0_12_port, A2 => n1617, B1 => 
                           REG_2_12_port, B2 => n8, ZN => n1173);
   U1802 : NAND4_X1 port map( A1 => n1176, A2 => n1175, A3 => n1174, A4 => 
                           n1173, ZN => n1182);
   U1803 : AOI22_X1 port map( A1 => REG_13_12_port, A2 => n4, B1 => 
                           REG_15_12_port, B2 => n1597, ZN => n1180);
   U1804 : AOI22_X1 port map( A1 => REG_9_12_port, A2 => n1604, B1 => 
                           REG_11_12_port, B2 => n5, ZN => n1179);
   U1805 : AOI22_X1 port map( A1 => REG_12_12_port, A2 => n7, B1 => 
                           REG_14_12_port, B2 => n1609, ZN => n1178);
   U1806 : AOI22_X1 port map( A1 => REG_8_12_port, A2 => n1617, B1 => 
                           REG_10_12_port, B2 => n8, ZN => n1177);
   U1807 : NAND4_X1 port map( A1 => n1180, A2 => n1179, A3 => n1178, A4 => 
                           n1177, ZN => n1181);
   U1808 : AOI22_X1 port map( A1 => n1182, A2 => n1619, B1 => n1181, B2 => 
                           n1618, ZN => n1183);
   U1809 : OAI221_X1 port map( B1 => n1587, B2 => n1185, C1 => n1585, C2 => 
                           n1184, A => n1183, ZN => N303);
   U1810 : AOI22_X1 port map( A1 => REG_21_13_port, A2 => n4, B1 => 
                           REG_23_13_port, B2 => n1597, ZN => n1189);
   U1811 : AOI22_X1 port map( A1 => REG_17_13_port, A2 => n1604, B1 => 
                           REG_19_13_port, B2 => n5, ZN => n1188);
   U1812 : AOI22_X1 port map( A1 => REG_20_13_port, A2 => n7, B1 => 
                           REG_22_13_port, B2 => n1609, ZN => n1187);
   U1813 : AOI22_X1 port map( A1 => REG_16_13_port, A2 => n1617, B1 => 
                           REG_18_13_port, B2 => n8, ZN => n1186);
   U1814 : AND4_X1 port map( A1 => n1189, A2 => n1188, A3 => n1187, A4 => n1186
                           , ZN => n1206);
   U1815 : AOI22_X1 port map( A1 => REG_29_13_port, A2 => n4, B1 => 
                           REG_31_13_port, B2 => n1597, ZN => n1193);
   U1816 : AOI22_X1 port map( A1 => REG_25_13_port, A2 => n1604, B1 => 
                           REG_27_13_port, B2 => n5, ZN => n1192);
   U1817 : AOI22_X1 port map( A1 => REG_28_13_port, A2 => n7, B1 => 
                           REG_30_13_port, B2 => n1609, ZN => n1191);
   U1818 : AOI22_X1 port map( A1 => REG_24_13_port, A2 => n1617, B1 => 
                           REG_26_13_port, B2 => n8, ZN => n1190);
   U1819 : AND4_X1 port map( A1 => n1193, A2 => n1192, A3 => n1191, A4 => n1190
                           , ZN => n1205);
   U1820 : AOI22_X1 port map( A1 => REG_5_13_port, A2 => n4, B1 => 
                           REG_7_13_port, B2 => n1597, ZN => n1197);
   U1821 : AOI22_X1 port map( A1 => REG_1_13_port, A2 => n1604, B1 => 
                           REG_3_13_port, B2 => n5, ZN => n1196);
   U1822 : AOI22_X1 port map( A1 => REG_4_13_port, A2 => n7, B1 => 
                           REG_6_13_port, B2 => n1609, ZN => n1195);
   U1823 : AOI22_X1 port map( A1 => REG_0_13_port, A2 => n1617, B1 => 
                           REG_2_13_port, B2 => n8, ZN => n1194);
   U1824 : NAND4_X1 port map( A1 => n1197, A2 => n1196, A3 => n1195, A4 => 
                           n1194, ZN => n1203);
   U1825 : AOI22_X1 port map( A1 => REG_13_13_port, A2 => n4, B1 => 
                           REG_15_13_port, B2 => n1596, ZN => n1201);
   U1826 : AOI22_X1 port map( A1 => REG_9_13_port, A2 => n1603, B1 => 
                           REG_11_13_port, B2 => n5, ZN => n1200);
   U1827 : AOI22_X1 port map( A1 => REG_12_13_port, A2 => n7, B1 => 
                           REG_14_13_port, B2 => n1609, ZN => n1199);
   U1828 : AOI22_X1 port map( A1 => REG_8_13_port, A2 => n1617, B1 => 
                           REG_10_13_port, B2 => n8, ZN => n1198);
   U1829 : NAND4_X1 port map( A1 => n1201, A2 => n1200, A3 => n1199, A4 => 
                           n1198, ZN => n1202);
   U1830 : AOI22_X1 port map( A1 => n1203, A2 => n1619, B1 => n1202, B2 => 
                           n1618, ZN => n1204);
   U1831 : OAI221_X1 port map( B1 => n1587, B2 => n1206, C1 => n1585, C2 => 
                           n1205, A => n1204, ZN => N302);
   U1832 : AOI22_X1 port map( A1 => REG_21_14_port, A2 => n4, B1 => 
                           REG_23_14_port, B2 => n1596, ZN => n1210);
   U1833 : AOI22_X1 port map( A1 => REG_17_14_port, A2 => n1603, B1 => 
                           REG_19_14_port, B2 => n5, ZN => n1209);
   U1834 : AOI22_X1 port map( A1 => REG_20_14_port, A2 => n7, B1 => 
                           REG_22_14_port, B2 => n1609, ZN => n1208);
   U1835 : AOI22_X1 port map( A1 => REG_16_14_port, A2 => n1617, B1 => 
                           REG_18_14_port, B2 => n8, ZN => n1207);
   U1836 : AND4_X1 port map( A1 => n1210, A2 => n1209, A3 => n1208, A4 => n1207
                           , ZN => n1227);
   U1837 : AOI22_X1 port map( A1 => REG_29_14_port, A2 => n4, B1 => 
                           REG_31_14_port, B2 => n1596, ZN => n1214);
   U1838 : AOI22_X1 port map( A1 => REG_25_14_port, A2 => n1603, B1 => 
                           REG_27_14_port, B2 => n5, ZN => n1213);
   U1839 : AOI22_X1 port map( A1 => REG_28_14_port, A2 => n7, B1 => 
                           REG_30_14_port, B2 => n1609, ZN => n1212);
   U1840 : AOI22_X1 port map( A1 => REG_24_14_port, A2 => n1617, B1 => 
                           REG_26_14_port, B2 => n8, ZN => n1211);
   U1841 : AND4_X1 port map( A1 => n1214, A2 => n1213, A3 => n1212, A4 => n1211
                           , ZN => n1226);
   U1842 : AOI22_X1 port map( A1 => REG_5_14_port, A2 => n4, B1 => 
                           REG_7_14_port, B2 => n1596, ZN => n1218);
   U1843 : AOI22_X1 port map( A1 => REG_1_14_port, A2 => n1603, B1 => 
                           REG_3_14_port, B2 => n5, ZN => n1217);
   U1844 : AOI22_X1 port map( A1 => REG_4_14_port, A2 => n7, B1 => 
                           REG_6_14_port, B2 => n1609, ZN => n1216);
   U1845 : AOI22_X1 port map( A1 => REG_0_14_port, A2 => n1617, B1 => 
                           REG_2_14_port, B2 => n8, ZN => n1215);
   U1846 : NAND4_X1 port map( A1 => n1218, A2 => n1217, A3 => n1216, A4 => 
                           n1215, ZN => n1224);
   U1847 : AOI22_X1 port map( A1 => REG_13_14_port, A2 => n4, B1 => 
                           REG_15_14_port, B2 => n1596, ZN => n1222);
   U1848 : AOI22_X1 port map( A1 => REG_9_14_port, A2 => n1603, B1 => 
                           REG_11_14_port, B2 => n5, ZN => n1221);
   U1849 : AOI22_X1 port map( A1 => REG_12_14_port, A2 => n7, B1 => 
                           REG_14_14_port, B2 => n1609, ZN => n1220);
   U1850 : AOI22_X1 port map( A1 => REG_8_14_port, A2 => n1617, B1 => 
                           REG_10_14_port, B2 => n8, ZN => n1219);
   U1851 : NAND4_X1 port map( A1 => n1222, A2 => n1221, A3 => n1220, A4 => 
                           n1219, ZN => n1223);
   U1852 : AOI22_X1 port map( A1 => n1224, A2 => n1619, B1 => n1223, B2 => 
                           n1618, ZN => n1225);
   U1853 : OAI221_X1 port map( B1 => n1587, B2 => n1227, C1 => n1585, C2 => 
                           n1226, A => n1225, ZN => N301);
   U1854 : AOI22_X1 port map( A1 => REG_21_15_port, A2 => n4, B1 => 
                           REG_23_15_port, B2 => n1596, ZN => n1231);
   U1855 : AOI22_X1 port map( A1 => REG_17_15_port, A2 => n1603, B1 => 
                           REG_19_15_port, B2 => n5, ZN => n1230);
   U1856 : AOI22_X1 port map( A1 => REG_20_15_port, A2 => n7, B1 => 
                           REG_22_15_port, B2 => n1609, ZN => n1229);
   U1857 : AOI22_X1 port map( A1 => REG_16_15_port, A2 => n1617, B1 => 
                           REG_18_15_port, B2 => n8, ZN => n1228);
   U1858 : AND4_X1 port map( A1 => n1231, A2 => n1230, A3 => n1229, A4 => n1228
                           , ZN => n1248);
   U1859 : AOI22_X1 port map( A1 => REG_29_15_port, A2 => n4, B1 => 
                           REG_31_15_port, B2 => n1596, ZN => n1235);
   U1860 : AOI22_X1 port map( A1 => REG_25_15_port, A2 => n1603, B1 => 
                           REG_27_15_port, B2 => n5, ZN => n1234);
   U1861 : AOI22_X1 port map( A1 => REG_28_15_port, A2 => n7, B1 => 
                           REG_30_15_port, B2 => n1609, ZN => n1233);
   U1862 : AOI22_X1 port map( A1 => REG_24_15_port, A2 => n1617, B1 => 
                           REG_26_15_port, B2 => n8, ZN => n1232);
   U1863 : AND4_X1 port map( A1 => n1235, A2 => n1234, A3 => n1233, A4 => n1232
                           , ZN => n1247);
   U1864 : AOI22_X1 port map( A1 => REG_5_15_port, A2 => n4, B1 => 
                           REG_7_15_port, B2 => n1596, ZN => n1239);
   U1865 : AOI22_X1 port map( A1 => REG_1_15_port, A2 => n1603, B1 => 
                           REG_3_15_port, B2 => n5, ZN => n1238);
   U1866 : AOI22_X1 port map( A1 => REG_4_15_port, A2 => n7, B1 => 
                           REG_6_15_port, B2 => n1609, ZN => n1237);
   U1867 : AOI22_X1 port map( A1 => REG_0_15_port, A2 => n1617, B1 => 
                           REG_2_15_port, B2 => n8, ZN => n1236);
   U1868 : NAND4_X1 port map( A1 => n1239, A2 => n1238, A3 => n1237, A4 => 
                           n1236, ZN => n1245);
   U1869 : AOI22_X1 port map( A1 => REG_13_15_port, A2 => n4, B1 => 
                           REG_15_15_port, B2 => n1596, ZN => n1243);
   U1870 : AOI22_X1 port map( A1 => REG_9_15_port, A2 => n1603, B1 => 
                           REG_11_15_port, B2 => n5, ZN => n1242);
   U1871 : AOI22_X1 port map( A1 => REG_12_15_port, A2 => n7, B1 => 
                           REG_14_15_port, B2 => n1609, ZN => n1241);
   U1872 : AOI22_X1 port map( A1 => REG_8_15_port, A2 => n1617, B1 => 
                           REG_10_15_port, B2 => n8, ZN => n1240);
   U1873 : NAND4_X1 port map( A1 => n1243, A2 => n1242, A3 => n1241, A4 => 
                           n1240, ZN => n1244);
   U1874 : AOI22_X1 port map( A1 => n1245, A2 => n1619, B1 => n1244, B2 => 
                           n1618, ZN => n1246);
   U1875 : OAI221_X1 port map( B1 => n1587, B2 => n1248, C1 => n1585, C2 => 
                           n1247, A => n1246, ZN => N300);
   U1876 : AOI22_X1 port map( A1 => REG_21_16_port, A2 => n4, B1 => 
                           REG_23_16_port, B2 => n1596, ZN => n1252);
   U1877 : AOI22_X1 port map( A1 => REG_17_16_port, A2 => n1603, B1 => 
                           REG_19_16_port, B2 => n5, ZN => n1251);
   U1878 : AOI22_X1 port map( A1 => REG_20_16_port, A2 => n7, B1 => 
                           REG_22_16_port, B2 => n1609, ZN => n1250);
   U1879 : AOI22_X1 port map( A1 => REG_16_16_port, A2 => n1617, B1 => 
                           REG_18_16_port, B2 => n8, ZN => n1249);
   U1880 : AND4_X1 port map( A1 => n1252, A2 => n1251, A3 => n1250, A4 => n1249
                           , ZN => n1269);
   U1881 : AOI22_X1 port map( A1 => REG_29_16_port, A2 => n4, B1 => 
                           REG_31_16_port, B2 => n1596, ZN => n1256);
   U1882 : AOI22_X1 port map( A1 => REG_25_16_port, A2 => n1603, B1 => 
                           REG_27_16_port, B2 => n5, ZN => n1255);
   U1883 : AOI22_X1 port map( A1 => REG_28_16_port, A2 => n7, B1 => 
                           REG_30_16_port, B2 => n1609, ZN => n1254);
   U1884 : AOI22_X1 port map( A1 => REG_24_16_port, A2 => n1617, B1 => 
                           REG_26_16_port, B2 => n8, ZN => n1253);
   U1885 : AND4_X1 port map( A1 => n1256, A2 => n1255, A3 => n1254, A4 => n1253
                           , ZN => n1268);
   U1886 : AOI22_X1 port map( A1 => REG_5_16_port, A2 => n1598, B1 => 
                           REG_7_16_port, B2 => n1593, ZN => n1260);
   U1887 : AOI22_X1 port map( A1 => REG_1_16_port, A2 => n1602, B1 => 
                           REG_3_16_port, B2 => n5, ZN => n1259);
   U1888 : AOI22_X1 port map( A1 => REG_4_16_port, A2 => n7, B1 => 
                           REG_6_16_port, B2 => n1605, ZN => n1258);
   U1889 : AOI22_X1 port map( A1 => REG_0_16_port, A2 => n1616, B1 => 
                           REG_2_16_port, B2 => n1611, ZN => n1257);
   U1890 : NAND4_X1 port map( A1 => n1260, A2 => n1259, A3 => n1258, A4 => 
                           n1257, ZN => n1266);
   U1891 : AOI22_X1 port map( A1 => REG_13_16_port, A2 => n1598, B1 => 
                           REG_15_16_port, B2 => n1593, ZN => n1264);
   U1892 : AOI22_X1 port map( A1 => REG_9_16_port, A2 => n1602, B1 => 
                           REG_11_16_port, B2 => n5, ZN => n1263);
   U1893 : AOI22_X1 port map( A1 => REG_12_16_port, A2 => n7, B1 => 
                           REG_14_16_port, B2 => n1605, ZN => n1262);
   U1894 : AOI22_X1 port map( A1 => REG_8_16_port, A2 => n1616, B1 => 
                           REG_10_16_port, B2 => n1611, ZN => n1261);
   U1895 : NAND4_X1 port map( A1 => n1264, A2 => n1263, A3 => n1262, A4 => 
                           n1261, ZN => n1265);
   U1896 : AOI22_X1 port map( A1 => n1266, A2 => n1619, B1 => n1265, B2 => 
                           n1618, ZN => n1267);
   U1897 : OAI221_X1 port map( B1 => n1587, B2 => n1269, C1 => n1585, C2 => 
                           n1268, A => n1267, ZN => N299);
   U1898 : AOI22_X1 port map( A1 => REG_21_17_port, A2 => n1598, B1 => 
                           REG_23_17_port, B2 => n1593, ZN => n1273);
   U1899 : AOI22_X1 port map( A1 => REG_17_17_port, A2 => n1602, B1 => 
                           REG_19_17_port, B2 => n5, ZN => n1272);
   U1900 : AOI22_X1 port map( A1 => REG_20_17_port, A2 => n7, B1 => 
                           REG_22_17_port, B2 => n1605, ZN => n1271);
   U1901 : AOI22_X1 port map( A1 => REG_16_17_port, A2 => n1616, B1 => 
                           REG_18_17_port, B2 => n1611, ZN => n1270);
   U1902 : AND4_X1 port map( A1 => n1273, A2 => n1272, A3 => n1271, A4 => n1270
                           , ZN => n1290);
   U1903 : AOI22_X1 port map( A1 => REG_29_17_port, A2 => n1598, B1 => 
                           REG_31_17_port, B2 => n1593, ZN => n1277);
   U1904 : AOI22_X1 port map( A1 => REG_25_17_port, A2 => n1602, B1 => 
                           REG_27_17_port, B2 => n5, ZN => n1276);
   U1905 : AOI22_X1 port map( A1 => REG_28_17_port, A2 => n7, B1 => 
                           REG_30_17_port, B2 => n1605, ZN => n1275);
   U1906 : AOI22_X1 port map( A1 => REG_24_17_port, A2 => n1616, B1 => 
                           REG_26_17_port, B2 => n1611, ZN => n1274);
   U1907 : AND4_X1 port map( A1 => n1277, A2 => n1276, A3 => n1275, A4 => n1274
                           , ZN => n1289);
   U1908 : AOI22_X1 port map( A1 => REG_5_17_port, A2 => n1598, B1 => 
                           REG_7_17_port, B2 => n1593, ZN => n1281);
   U1909 : AOI22_X1 port map( A1 => REG_1_17_port, A2 => n1602, B1 => 
                           REG_3_17_port, B2 => n5, ZN => n1280);
   U1910 : AOI22_X1 port map( A1 => REG_4_17_port, A2 => n7, B1 => 
                           REG_6_17_port, B2 => n1605, ZN => n1279);
   U1911 : AOI22_X1 port map( A1 => REG_0_17_port, A2 => n1616, B1 => 
                           REG_2_17_port, B2 => n1611, ZN => n1278);
   U1912 : NAND4_X1 port map( A1 => n1281, A2 => n1280, A3 => n1279, A4 => 
                           n1278, ZN => n1287);
   U1913 : AOI22_X1 port map( A1 => REG_13_17_port, A2 => n1598, B1 => 
                           REG_15_17_port, B2 => n1593, ZN => n1285);
   U1914 : AOI22_X1 port map( A1 => REG_9_17_port, A2 => n1602, B1 => 
                           REG_11_17_port, B2 => n5, ZN => n1284);
   U1915 : AOI22_X1 port map( A1 => REG_12_17_port, A2 => n7, B1 => 
                           REG_14_17_port, B2 => n1605, ZN => n1283);
   U1916 : AOI22_X1 port map( A1 => REG_8_17_port, A2 => n1616, B1 => 
                           REG_10_17_port, B2 => n1611, ZN => n1282);
   U1917 : NAND4_X1 port map( A1 => n1285, A2 => n1284, A3 => n1283, A4 => 
                           n1282, ZN => n1286);
   U1918 : AOI22_X1 port map( A1 => n1287, A2 => n1619, B1 => n1286, B2 => 
                           n1618, ZN => n1288);
   U1919 : OAI221_X1 port map( B1 => n1587, B2 => n1290, C1 => n1585, C2 => 
                           n1289, A => n1288, ZN => N298);
   U1920 : AOI22_X1 port map( A1 => REG_21_18_port, A2 => n1598, B1 => 
                           REG_23_18_port, B2 => n1593, ZN => n1294);
   U1921 : AOI22_X1 port map( A1 => REG_17_18_port, A2 => n1602, B1 => 
                           REG_19_18_port, B2 => n5, ZN => n1293);
   U1922 : AOI22_X1 port map( A1 => REG_20_18_port, A2 => n7, B1 => 
                           REG_22_18_port, B2 => n1605, ZN => n1292);
   U1923 : AOI22_X1 port map( A1 => REG_16_18_port, A2 => n1616, B1 => 
                           REG_18_18_port, B2 => n1611, ZN => n1291);
   U1924 : AND4_X1 port map( A1 => n1294, A2 => n1293, A3 => n1292, A4 => n1291
                           , ZN => n1311);
   U1925 : AOI22_X1 port map( A1 => REG_29_18_port, A2 => n1598, B1 => 
                           REG_31_18_port, B2 => n1593, ZN => n1298);
   U1926 : AOI22_X1 port map( A1 => REG_25_18_port, A2 => n1602, B1 => 
                           REG_27_18_port, B2 => n5, ZN => n1297);
   U1927 : AOI22_X1 port map( A1 => REG_28_18_port, A2 => n7, B1 => 
                           REG_30_18_port, B2 => n1605, ZN => n1296);
   U1928 : AOI22_X1 port map( A1 => REG_24_18_port, A2 => n1616, B1 => 
                           REG_26_18_port, B2 => n1611, ZN => n1295);
   U1929 : AND4_X1 port map( A1 => n1298, A2 => n1297, A3 => n1296, A4 => n1295
                           , ZN => n1310);
   U1930 : AOI22_X1 port map( A1 => REG_5_18_port, A2 => n1598, B1 => 
                           REG_7_18_port, B2 => n1593, ZN => n1302);
   U1931 : AOI22_X1 port map( A1 => REG_1_18_port, A2 => n1602, B1 => 
                           REG_3_18_port, B2 => n5, ZN => n1301);
   U1932 : AOI22_X1 port map( A1 => REG_4_18_port, A2 => n7, B1 => 
                           REG_6_18_port, B2 => n1605, ZN => n1300);
   U1933 : AOI22_X1 port map( A1 => REG_0_18_port, A2 => n1616, B1 => 
                           REG_2_18_port, B2 => n1611, ZN => n1299);
   U1934 : NAND4_X1 port map( A1 => n1302, A2 => n1301, A3 => n1300, A4 => 
                           n1299, ZN => n1308);
   U1935 : AOI22_X1 port map( A1 => REG_13_18_port, A2 => n1598, B1 => 
                           REG_15_18_port, B2 => n1593, ZN => n1306);
   U1936 : AOI22_X1 port map( A1 => REG_9_18_port, A2 => n1602, B1 => 
                           REG_11_18_port, B2 => n5, ZN => n1305);
   U1937 : AOI22_X1 port map( A1 => REG_12_18_port, A2 => n7, B1 => 
                           REG_14_18_port, B2 => n1605, ZN => n1304);
   U1938 : AOI22_X1 port map( A1 => REG_8_18_port, A2 => n1616, B1 => 
                           REG_10_18_port, B2 => n1611, ZN => n1303);
   U1939 : NAND4_X1 port map( A1 => n1306, A2 => n1305, A3 => n1304, A4 => 
                           n1303, ZN => n1307);
   U1940 : AOI22_X1 port map( A1 => n1308, A2 => n1619, B1 => n1307, B2 => 
                           n1618, ZN => n1309);
   U1941 : OAI221_X1 port map( B1 => n1587, B2 => n1311, C1 => n1585, C2 => 
                           n1310, A => n1309, ZN => N297);
   U1942 : AOI22_X1 port map( A1 => REG_21_19_port, A2 => n1598, B1 => 
                           REG_23_19_port, B2 => n1593, ZN => n1315);
   U1943 : AOI22_X1 port map( A1 => REG_17_19_port, A2 => n1602, B1 => 
                           REG_19_19_port, B2 => n5, ZN => n1314);
   U1944 : AOI22_X1 port map( A1 => REG_20_19_port, A2 => n7, B1 => 
                           REG_22_19_port, B2 => n1605, ZN => n1313);
   U1945 : AOI22_X1 port map( A1 => REG_16_19_port, A2 => n1616, B1 => 
                           REG_18_19_port, B2 => n1611, ZN => n1312);
   U1946 : AND4_X1 port map( A1 => n1315, A2 => n1314, A3 => n1313, A4 => n1312
                           , ZN => n1332);
   U1947 : AOI22_X1 port map( A1 => REG_29_19_port, A2 => n1598, B1 => 
                           REG_31_19_port, B2 => n1593, ZN => n1319);
   U1948 : AOI22_X1 port map( A1 => REG_25_19_port, A2 => n1602, B1 => 
                           REG_27_19_port, B2 => n5, ZN => n1318);
   U1949 : AOI22_X1 port map( A1 => REG_28_19_port, A2 => n1610, B1 => 
                           REG_30_19_port, B2 => n1605, ZN => n1317);
   U1950 : AOI22_X1 port map( A1 => REG_24_19_port, A2 => n1615, B1 => 
                           REG_26_19_port, B2 => n1611, ZN => n1316);
   U1951 : AND4_X1 port map( A1 => n1319, A2 => n1318, A3 => n1317, A4 => n1316
                           , ZN => n1331);
   U1952 : AOI22_X1 port map( A1 => REG_5_19_port, A2 => n1598, B1 => 
                           REG_7_19_port, B2 => n1593, ZN => n1323);
   U1953 : AOI22_X1 port map( A1 => REG_1_19_port, A2 => n1602, B1 => 
                           REG_3_19_port, B2 => n5, ZN => n1322);
   U1954 : AOI22_X1 port map( A1 => REG_4_19_port, A2 => n1610, B1 => 
                           REG_6_19_port, B2 => n1605, ZN => n1321);
   U1955 : AOI22_X1 port map( A1 => REG_0_19_port, A2 => n1615, B1 => 
                           REG_2_19_port, B2 => n1611, ZN => n1320);
   U1956 : NAND4_X1 port map( A1 => n1323, A2 => n1322, A3 => n1321, A4 => 
                           n1320, ZN => n1329);
   U1957 : AOI22_X1 port map( A1 => REG_13_19_port, A2 => n1598, B1 => 
                           REG_15_19_port, B2 => n1593, ZN => n1327);
   U1958 : AOI22_X1 port map( A1 => REG_9_19_port, A2 => n1602, B1 => 
                           REG_11_19_port, B2 => n5, ZN => n1326);
   U1959 : AOI22_X1 port map( A1 => REG_12_19_port, A2 => n1610, B1 => 
                           REG_14_19_port, B2 => n1605, ZN => n1325);
   U1960 : AOI22_X1 port map( A1 => REG_8_19_port, A2 => n1615, B1 => 
                           REG_10_19_port, B2 => n1611, ZN => n1324);
   U1961 : NAND4_X1 port map( A1 => n1327, A2 => n1326, A3 => n1325, A4 => 
                           n1324, ZN => n1328);
   U1962 : AOI22_X1 port map( A1 => n1329, A2 => n1619, B1 => n1328, B2 => 
                           n1618, ZN => n1330);
   U1963 : OAI221_X1 port map( B1 => n1587, B2 => n1332, C1 => n1585, C2 => 
                           n1331, A => n1330, ZN => N296);
   U1964 : AOI22_X1 port map( A1 => REG_21_20_port, A2 => n1598, B1 => 
                           REG_23_20_port, B2 => n1593, ZN => n1336);
   U1965 : AOI22_X1 port map( A1 => REG_17_20_port, A2 => n1602, B1 => 
                           REG_19_20_port, B2 => n5, ZN => n1335);
   U1966 : AOI22_X1 port map( A1 => REG_20_20_port, A2 => n1610, B1 => 
                           REG_22_20_port, B2 => n1605, ZN => n1334);
   U1967 : AOI22_X1 port map( A1 => REG_16_20_port, A2 => n1615, B1 => 
                           REG_18_20_port, B2 => n1611, ZN => n1333);
   U1968 : AND4_X1 port map( A1 => n1336, A2 => n1335, A3 => n1334, A4 => n1333
                           , ZN => n1353);
   U1969 : AOI22_X1 port map( A1 => REG_29_20_port, A2 => n1598, B1 => 
                           REG_31_20_port, B2 => n1593, ZN => n1340);
   U1970 : AOI22_X1 port map( A1 => REG_25_20_port, A2 => n1602, B1 => 
                           REG_27_20_port, B2 => n5, ZN => n1339);
   U1971 : AOI22_X1 port map( A1 => REG_28_20_port, A2 => n1610, B1 => 
                           REG_30_20_port, B2 => n1605, ZN => n1338);
   U1972 : AOI22_X1 port map( A1 => REG_24_20_port, A2 => n1615, B1 => 
                           REG_26_20_port, B2 => n1611, ZN => n1337);
   U1973 : AND4_X1 port map( A1 => n1340, A2 => n1339, A3 => n1338, A4 => n1337
                           , ZN => n1352);
   U1974 : AOI22_X1 port map( A1 => REG_5_20_port, A2 => n1598, B1 => 
                           REG_7_20_port, B2 => n1593, ZN => n1344);
   U1975 : AOI22_X1 port map( A1 => REG_1_20_port, A2 => n1602, B1 => 
                           REG_3_20_port, B2 => n5, ZN => n1343);
   U1976 : AOI22_X1 port map( A1 => REG_4_20_port, A2 => n1610, B1 => 
                           REG_6_20_port, B2 => n1605, ZN => n1342);
   U1977 : AOI22_X1 port map( A1 => REG_0_20_port, A2 => n1615, B1 => 
                           REG_2_20_port, B2 => n1611, ZN => n1341);
   U1978 : NAND4_X1 port map( A1 => n1344, A2 => n1343, A3 => n1342, A4 => 
                           n1341, ZN => n1350);
   U1979 : AOI22_X1 port map( A1 => REG_13_20_port, A2 => n1598, B1 => 
                           REG_15_20_port, B2 => n1593, ZN => n1348);
   U1980 : AOI22_X1 port map( A1 => REG_9_20_port, A2 => n1602, B1 => 
                           REG_11_20_port, B2 => n5, ZN => n1347);
   U1981 : AOI22_X1 port map( A1 => REG_12_20_port, A2 => n1610, B1 => 
                           REG_14_20_port, B2 => n1605, ZN => n1346);
   U1982 : AOI22_X1 port map( A1 => REG_8_20_port, A2 => n1615, B1 => 
                           REG_10_20_port, B2 => n1611, ZN => n1345);
   U1983 : NAND4_X1 port map( A1 => n1348, A2 => n1347, A3 => n1346, A4 => 
                           n1345, ZN => n1349);
   U1984 : AOI22_X1 port map( A1 => n1350, A2 => n1619, B1 => n1349, B2 => 
                           n1618, ZN => n1351);
   U1985 : OAI221_X1 port map( B1 => n1587, B2 => n1353, C1 => n1585, C2 => 
                           n1352, A => n1351, ZN => N295);
   U1986 : AOI22_X1 port map( A1 => REG_21_21_port, A2 => n1598, B1 => 
                           REG_23_21_port, B2 => n1593, ZN => n1357);
   U1987 : AOI22_X1 port map( A1 => REG_17_21_port, A2 => n1602, B1 => 
                           REG_19_21_port, B2 => n5, ZN => n1356);
   U1988 : AOI22_X1 port map( A1 => REG_20_21_port, A2 => n1610, B1 => 
                           REG_22_21_port, B2 => n1605, ZN => n1355);
   U1989 : AOI22_X1 port map( A1 => REG_16_21_port, A2 => n1615, B1 => 
                           REG_18_21_port, B2 => n1611, ZN => n1354);
   U1990 : AND4_X1 port map( A1 => n1357, A2 => n1356, A3 => n1355, A4 => n1354
                           , ZN => n1374);
   U1991 : AOI22_X1 port map( A1 => REG_29_21_port, A2 => n1598, B1 => 
                           REG_31_21_port, B2 => n1593, ZN => n1361);
   U1992 : AOI22_X1 port map( A1 => REG_25_21_port, A2 => n1602, B1 => 
                           REG_27_21_port, B2 => n5, ZN => n1360);
   U1993 : AOI22_X1 port map( A1 => REG_28_21_port, A2 => n1610, B1 => 
                           REG_30_21_port, B2 => n1605, ZN => n1359);
   U1994 : AOI22_X1 port map( A1 => REG_24_21_port, A2 => n1615, B1 => 
                           REG_26_21_port, B2 => n1611, ZN => n1358);
   U1995 : AND4_X1 port map( A1 => n1361, A2 => n1360, A3 => n1359, A4 => n1358
                           , ZN => n1373);
   U1996 : AOI22_X1 port map( A1 => REG_5_21_port, A2 => n1598, B1 => 
                           REG_7_21_port, B2 => n1593, ZN => n1365);
   U1997 : AOI22_X1 port map( A1 => REG_1_21_port, A2 => n1602, B1 => 
                           REG_3_21_port, B2 => n5, ZN => n1364);
   U1998 : AOI22_X1 port map( A1 => REG_4_21_port, A2 => n1610, B1 => 
                           REG_6_21_port, B2 => n1605, ZN => n1363);
   U1999 : AOI22_X1 port map( A1 => REG_0_21_port, A2 => n1615, B1 => 
                           REG_2_21_port, B2 => n1611, ZN => n1362);
   U2000 : NAND4_X1 port map( A1 => n1365, A2 => n1364, A3 => n1363, A4 => 
                           n1362, ZN => n1371);
   U2001 : AOI22_X1 port map( A1 => REG_13_21_port, A2 => n1598, B1 => 
                           REG_15_21_port, B2 => n1593, ZN => n1369);
   U2002 : AOI22_X1 port map( A1 => REG_9_21_port, A2 => n1602, B1 => 
                           REG_11_21_port, B2 => n5, ZN => n1368);
   U2003 : AOI22_X1 port map( A1 => REG_12_21_port, A2 => n1610, B1 => 
                           REG_14_21_port, B2 => n1605, ZN => n1367);
   U2004 : AOI22_X1 port map( A1 => REG_8_21_port, A2 => n1615, B1 => 
                           REG_10_21_port, B2 => n1611, ZN => n1366);
   U2005 : NAND4_X1 port map( A1 => n1369, A2 => n1368, A3 => n1367, A4 => 
                           n1366, ZN => n1370);
   U2006 : AOI22_X1 port map( A1 => n1371, A2 => n1619, B1 => n1370, B2 => 
                           n1618, ZN => n1372);
   U2007 : OAI221_X1 port map( B1 => n1587, B2 => n1374, C1 => n1585, C2 => 
                           n1373, A => n1372, ZN => N294);
   U2008 : AOI22_X1 port map( A1 => REG_21_22_port, A2 => n1598, B1 => 
                           REG_23_22_port, B2 => n1593, ZN => n1378);
   U2009 : AOI22_X1 port map( A1 => REG_17_22_port, A2 => n1602, B1 => 
                           REG_19_22_port, B2 => n1599, ZN => n1377);
   U2010 : AOI22_X1 port map( A1 => REG_20_22_port, A2 => n1610, B1 => 
                           REG_22_22_port, B2 => n1605, ZN => n1376);
   U2011 : AOI22_X1 port map( A1 => REG_16_22_port, A2 => n1614, B1 => 
                           REG_18_22_port, B2 => n1611, ZN => n1375);
   U2012 : AND4_X1 port map( A1 => n1378, A2 => n1377, A3 => n1376, A4 => n1375
                           , ZN => n1395);
   U2013 : AOI22_X1 port map( A1 => REG_29_22_port, A2 => n1598, B1 => 
                           REG_31_22_port, B2 => n1593, ZN => n1382);
   U2014 : AOI22_X1 port map( A1 => REG_25_22_port, A2 => n1602, B1 => 
                           REG_27_22_port, B2 => n1599, ZN => n1381);
   U2015 : AOI22_X1 port map( A1 => REG_28_22_port, A2 => n1610, B1 => 
                           REG_30_22_port, B2 => n1605, ZN => n1380);
   U2016 : AOI22_X1 port map( A1 => REG_24_22_port, A2 => n1614, B1 => 
                           REG_26_22_port, B2 => n1611, ZN => n1379);
   U2017 : AND4_X1 port map( A1 => n1382, A2 => n1381, A3 => n1380, A4 => n1379
                           , ZN => n1394);
   U2018 : AOI22_X1 port map( A1 => REG_5_22_port, A2 => n1598, B1 => 
                           REG_7_22_port, B2 => n1593, ZN => n1386);
   U2019 : AOI22_X1 port map( A1 => REG_1_22_port, A2 => n1602, B1 => 
                           REG_3_22_port, B2 => n1599, ZN => n1385);
   U2020 : AOI22_X1 port map( A1 => REG_4_22_port, A2 => n1610, B1 => 
                           REG_6_22_port, B2 => n1605, ZN => n1384);
   U2021 : AOI22_X1 port map( A1 => REG_0_22_port, A2 => n1614, B1 => 
                           REG_2_22_port, B2 => n1611, ZN => n1383);
   U2022 : NAND4_X1 port map( A1 => n1386, A2 => n1385, A3 => n1384, A4 => 
                           n1383, ZN => n1392);
   U2023 : AOI22_X1 port map( A1 => REG_13_22_port, A2 => n1598, B1 => 
                           REG_15_22_port, B2 => n1593, ZN => n1390);
   U2024 : AOI22_X1 port map( A1 => REG_9_22_port, A2 => n1602, B1 => 
                           REG_11_22_port, B2 => n1599, ZN => n1389);
   U2025 : AOI22_X1 port map( A1 => REG_12_22_port, A2 => n1610, B1 => 
                           REG_14_22_port, B2 => n1605, ZN => n1388);
   U2026 : AOI22_X1 port map( A1 => REG_8_22_port, A2 => n1614, B1 => 
                           REG_10_22_port, B2 => n1611, ZN => n1387);
   U2027 : NAND4_X1 port map( A1 => n1390, A2 => n1389, A3 => n1388, A4 => 
                           n1387, ZN => n1391);
   U2028 : AOI22_X1 port map( A1 => n1392, A2 => n1619, B1 => n1391, B2 => 
                           n1581, ZN => n1393);
   U2029 : OAI221_X1 port map( B1 => n1587, B2 => n1395, C1 => n1585, C2 => 
                           n1394, A => n1393, ZN => N293);
   U2030 : AOI22_X1 port map( A1 => REG_21_23_port, A2 => n1598, B1 => 
                           REG_23_23_port, B2 => n1593, ZN => n1399);
   U2031 : AOI22_X1 port map( A1 => REG_17_23_port, A2 => n1602, B1 => 
                           REG_19_23_port, B2 => n1599, ZN => n1398);
   U2032 : AOI22_X1 port map( A1 => REG_20_23_port, A2 => n1610, B1 => 
                           REG_22_23_port, B2 => n1605, ZN => n1397);
   U2033 : AOI22_X1 port map( A1 => REG_16_23_port, A2 => n1614, B1 => 
                           REG_18_23_port, B2 => n1611, ZN => n1396);
   U2034 : AND4_X1 port map( A1 => n1399, A2 => n1398, A3 => n1397, A4 => n1396
                           , ZN => n1416);
   U2035 : AOI22_X1 port map( A1 => REG_29_23_port, A2 => n1598, B1 => 
                           REG_31_23_port, B2 => n1593, ZN => n1403);
   U2036 : AOI22_X1 port map( A1 => REG_25_23_port, A2 => n1602, B1 => 
                           REG_27_23_port, B2 => n1599, ZN => n1402);
   U2037 : AOI22_X1 port map( A1 => REG_28_23_port, A2 => n1610, B1 => 
                           REG_30_23_port, B2 => n1605, ZN => n1401);
   U2038 : AOI22_X1 port map( A1 => REG_24_23_port, A2 => n1614, B1 => 
                           REG_26_23_port, B2 => n1611, ZN => n1400);
   U2039 : AND4_X1 port map( A1 => n1403, A2 => n1402, A3 => n1401, A4 => n1400
                           , ZN => n1415);
   U2040 : AOI22_X1 port map( A1 => REG_5_23_port, A2 => n1598, B1 => 
                           REG_7_23_port, B2 => n1593, ZN => n1407);
   U2041 : AOI22_X1 port map( A1 => REG_1_23_port, A2 => n1602, B1 => 
                           REG_3_23_port, B2 => n1599, ZN => n1406);
   U2042 : AOI22_X1 port map( A1 => REG_4_23_port, A2 => n1610, B1 => 
                           REG_6_23_port, B2 => n1605, ZN => n1405);
   U2043 : AOI22_X1 port map( A1 => REG_0_23_port, A2 => n1614, B1 => 
                           REG_2_23_port, B2 => n1611, ZN => n1404);
   U2044 : NAND4_X1 port map( A1 => n1407, A2 => n1406, A3 => n1405, A4 => 
                           n1404, ZN => n1413);
   U2045 : AOI22_X1 port map( A1 => REG_13_23_port, A2 => n1598, B1 => 
                           REG_15_23_port, B2 => n1593, ZN => n1411);
   U2046 : AOI22_X1 port map( A1 => REG_9_23_port, A2 => n1602, B1 => 
                           REG_11_23_port, B2 => n1599, ZN => n1410);
   U2047 : AOI22_X1 port map( A1 => REG_12_23_port, A2 => n1610, B1 => 
                           REG_14_23_port, B2 => n1605, ZN => n1409);
   U2048 : AOI22_X1 port map( A1 => REG_8_23_port, A2 => n1614, B1 => 
                           REG_10_23_port, B2 => n1611, ZN => n1408);
   U2049 : NAND4_X1 port map( A1 => n1411, A2 => n1410, A3 => n1409, A4 => 
                           n1408, ZN => n1412);
   U2050 : AOI22_X1 port map( A1 => n1413, A2 => n1619, B1 => n1412, B2 => 
                           n1581, ZN => n1414);
   U2051 : OAI221_X1 port map( B1 => n1587, B2 => n1416, C1 => n1585, C2 => 
                           n1415, A => n1414, ZN => N292);
   U2052 : AOI22_X1 port map( A1 => REG_21_24_port, A2 => n1598, B1 => 
                           REG_23_24_port, B2 => n1593, ZN => n1420);
   U2053 : AOI22_X1 port map( A1 => REG_17_24_port, A2 => n1602, B1 => 
                           REG_19_24_port, B2 => n1599, ZN => n1419);
   U2054 : AOI22_X1 port map( A1 => REG_20_24_port, A2 => n1610, B1 => 
                           REG_22_24_port, B2 => n1605, ZN => n1418);
   U2055 : AOI22_X1 port map( A1 => REG_16_24_port, A2 => n1614, B1 => 
                           REG_18_24_port, B2 => n1611, ZN => n1417);
   U2056 : AND4_X1 port map( A1 => n1420, A2 => n1419, A3 => n1418, A4 => n1417
                           , ZN => n1437);
   U2057 : AOI22_X1 port map( A1 => REG_29_24_port, A2 => n1598, B1 => 
                           REG_31_24_port, B2 => n1593, ZN => n1424);
   U2058 : AOI22_X1 port map( A1 => REG_25_24_port, A2 => n1602, B1 => 
                           REG_27_24_port, B2 => n1599, ZN => n1423);
   U2059 : AOI22_X1 port map( A1 => REG_28_24_port, A2 => n1610, B1 => 
                           REG_30_24_port, B2 => n1605, ZN => n1422);
   U2060 : AOI22_X1 port map( A1 => REG_24_24_port, A2 => n1614, B1 => 
                           REG_26_24_port, B2 => n1611, ZN => n1421);
   U2061 : AND4_X1 port map( A1 => n1424, A2 => n1423, A3 => n1422, A4 => n1421
                           , ZN => n1436);
   U2062 : AOI22_X1 port map( A1 => REG_5_24_port, A2 => n1598, B1 => 
                           REG_7_24_port, B2 => n1593, ZN => n1428);
   U2063 : AOI22_X1 port map( A1 => REG_1_24_port, A2 => n1602, B1 => 
                           REG_3_24_port, B2 => n1599, ZN => n1427);
   U2064 : AOI22_X1 port map( A1 => REG_4_24_port, A2 => n1610, B1 => 
                           REG_6_24_port, B2 => n1605, ZN => n1426);
   U2065 : AOI22_X1 port map( A1 => REG_0_24_port, A2 => n1614, B1 => 
                           REG_2_24_port, B2 => n1611, ZN => n1425);
   U2066 : NAND4_X1 port map( A1 => n1428, A2 => n1427, A3 => n1426, A4 => 
                           n1425, ZN => n1434);
   U2067 : AOI22_X1 port map( A1 => REG_13_24_port, A2 => n1598, B1 => 
                           REG_15_24_port, B2 => n1595, ZN => n1432);
   U2068 : AOI22_X1 port map( A1 => REG_9_24_port, A2 => n1601, B1 => 
                           REG_11_24_port, B2 => n1599, ZN => n1431);
   U2069 : AOI22_X1 port map( A1 => REG_12_24_port, A2 => n1610, B1 => 
                           REG_14_24_port, B2 => n1608, ZN => n1430);
   U2070 : AOI22_X1 port map( A1 => REG_8_24_port, A2 => n1612, B1 => 
                           REG_10_24_port, B2 => n8, ZN => n1429);
   U2071 : NAND4_X1 port map( A1 => n1432, A2 => n1431, A3 => n1430, A4 => 
                           n1429, ZN => n1433);
   U2072 : AOI22_X1 port map( A1 => n1434, A2 => n1619, B1 => n1433, B2 => 
                           n1581, ZN => n1435);
   U2073 : OAI221_X1 port map( B1 => n1587, B2 => n1437, C1 => n1585, C2 => 
                           n1436, A => n1435, ZN => N291);
   U2074 : AOI22_X1 port map( A1 => REG_21_25_port, A2 => n1598, B1 => 
                           REG_23_25_port, B2 => n1595, ZN => n1441);
   U2075 : AOI22_X1 port map( A1 => REG_17_25_port, A2 => n1601, B1 => 
                           REG_19_25_port, B2 => n1599, ZN => n1440);
   U2076 : AOI22_X1 port map( A1 => REG_20_25_port, A2 => n1610, B1 => 
                           REG_22_25_port, B2 => n1608, ZN => n1439);
   U2077 : AOI22_X1 port map( A1 => REG_16_25_port, A2 => n1612, B1 => 
                           REG_18_25_port, B2 => n8, ZN => n1438);
   U2078 : AND4_X1 port map( A1 => n1441, A2 => n1440, A3 => n1439, A4 => n1438
                           , ZN => n1458);
   U2079 : AOI22_X1 port map( A1 => REG_29_25_port, A2 => n1598, B1 => 
                           REG_31_25_port, B2 => n1595, ZN => n1445);
   U2080 : AOI22_X1 port map( A1 => REG_25_25_port, A2 => n1601, B1 => 
                           REG_27_25_port, B2 => n1599, ZN => n1444);
   U2081 : AOI22_X1 port map( A1 => REG_28_25_port, A2 => n1610, B1 => 
                           REG_30_25_port, B2 => n1608, ZN => n1443);
   U2082 : AOI22_X1 port map( A1 => REG_24_25_port, A2 => n1612, B1 => 
                           REG_26_25_port, B2 => n8, ZN => n1442);
   U2083 : AND4_X1 port map( A1 => n1445, A2 => n1444, A3 => n1443, A4 => n1442
                           , ZN => n1457);
   U2084 : AOI22_X1 port map( A1 => REG_5_25_port, A2 => n1598, B1 => 
                           REG_7_25_port, B2 => n1595, ZN => n1449);
   U2085 : AOI22_X1 port map( A1 => REG_1_25_port, A2 => n1601, B1 => 
                           REG_3_25_port, B2 => n1599, ZN => n1448);
   U2086 : AOI22_X1 port map( A1 => REG_4_25_port, A2 => n1610, B1 => 
                           REG_6_25_port, B2 => n1608, ZN => n1447);
   U2087 : AOI22_X1 port map( A1 => REG_0_25_port, A2 => n1612, B1 => 
                           REG_2_25_port, B2 => n8, ZN => n1446);
   U2088 : NAND4_X1 port map( A1 => n1449, A2 => n1448, A3 => n1447, A4 => 
                           n1446, ZN => n1455);
   U2089 : AOI22_X1 port map( A1 => REG_13_25_port, A2 => n1598, B1 => 
                           REG_15_25_port, B2 => n1595, ZN => n1453);
   U2090 : AOI22_X1 port map( A1 => REG_9_25_port, A2 => n1601, B1 => 
                           REG_11_25_port, B2 => n1599, ZN => n1452);
   U2091 : AOI22_X1 port map( A1 => REG_12_25_port, A2 => n1610, B1 => 
                           REG_14_25_port, B2 => n1608, ZN => n1451);
   U2092 : AOI22_X1 port map( A1 => REG_8_25_port, A2 => n1612, B1 => 
                           REG_10_25_port, B2 => n8, ZN => n1450);
   U2093 : NAND4_X1 port map( A1 => n1453, A2 => n1452, A3 => n1451, A4 => 
                           n1450, ZN => n1454);
   U2094 : AOI22_X1 port map( A1 => n1455, A2 => n1619, B1 => n1454, B2 => 
                           n1581, ZN => n1456);
   U2095 : OAI221_X1 port map( B1 => n1587, B2 => n1458, C1 => n1585, C2 => 
                           n1457, A => n1456, ZN => N290);
   U2096 : AOI22_X1 port map( A1 => REG_21_26_port, A2 => n1598, B1 => 
                           REG_23_26_port, B2 => n1595, ZN => n1462);
   U2097 : AOI22_X1 port map( A1 => REG_17_26_port, A2 => n1601, B1 => 
                           REG_19_26_port, B2 => n1599, ZN => n1461);
   U2098 : AOI22_X1 port map( A1 => REG_20_26_port, A2 => n1610, B1 => 
                           REG_22_26_port, B2 => n1608, ZN => n1460);
   U2099 : AOI22_X1 port map( A1 => REG_16_26_port, A2 => n1612, B1 => 
                           REG_18_26_port, B2 => n8, ZN => n1459);
   U2100 : AND4_X1 port map( A1 => n1462, A2 => n1461, A3 => n1460, A4 => n1459
                           , ZN => n1479);
   U2101 : AOI22_X1 port map( A1 => REG_29_26_port, A2 => n1598, B1 => 
                           REG_31_26_port, B2 => n1595, ZN => n1466);
   U2102 : AOI22_X1 port map( A1 => REG_25_26_port, A2 => n1601, B1 => 
                           REG_27_26_port, B2 => n1599, ZN => n1465);
   U2103 : AOI22_X1 port map( A1 => REG_28_26_port, A2 => n1610, B1 => 
                           REG_30_26_port, B2 => n1608, ZN => n1464);
   U2104 : AOI22_X1 port map( A1 => REG_24_26_port, A2 => n1612, B1 => 
                           REG_26_26_port, B2 => n8, ZN => n1463);
   U2105 : AND4_X1 port map( A1 => n1466, A2 => n1465, A3 => n1464, A4 => n1463
                           , ZN => n1478);
   U2106 : AOI22_X1 port map( A1 => REG_5_26_port, A2 => n1598, B1 => 
                           REG_7_26_port, B2 => n1595, ZN => n1470);
   U2107 : AOI22_X1 port map( A1 => REG_1_26_port, A2 => n1601, B1 => 
                           REG_3_26_port, B2 => n1599, ZN => n1469);
   U2108 : AOI22_X1 port map( A1 => REG_4_26_port, A2 => n1610, B1 => 
                           REG_6_26_port, B2 => n1608, ZN => n1468);
   U2109 : AOI22_X1 port map( A1 => REG_0_26_port, A2 => n1612, B1 => 
                           REG_2_26_port, B2 => n8, ZN => n1467);
   U2110 : NAND4_X1 port map( A1 => n1470, A2 => n1469, A3 => n1468, A4 => 
                           n1467, ZN => n1476);
   U2111 : AOI22_X1 port map( A1 => REG_13_26_port, A2 => n1598, B1 => 
                           REG_15_26_port, B2 => n1595, ZN => n1474);
   U2112 : AOI22_X1 port map( A1 => REG_9_26_port, A2 => n1601, B1 => 
                           REG_11_26_port, B2 => n1599, ZN => n1473);
   U2113 : AOI22_X1 port map( A1 => REG_12_26_port, A2 => n1610, B1 => 
                           REG_14_26_port, B2 => n1608, ZN => n1472);
   U2114 : AOI22_X1 port map( A1 => REG_8_26_port, A2 => n1612, B1 => 
                           REG_10_26_port, B2 => n8, ZN => n1471);
   U2115 : NAND4_X1 port map( A1 => n1474, A2 => n1473, A3 => n1472, A4 => 
                           n1471, ZN => n1475);
   U2116 : AOI22_X1 port map( A1 => n1476, A2 => n1619, B1 => n1475, B2 => 
                           n1581, ZN => n1477);
   U2117 : OAI221_X1 port map( B1 => n1587, B2 => n1479, C1 => n1585, C2 => 
                           n1478, A => n1477, ZN => N289);
   U2118 : AOI22_X1 port map( A1 => REG_21_27_port, A2 => n1598, B1 => 
                           REG_23_27_port, B2 => n1595, ZN => n1483);
   U2119 : AOI22_X1 port map( A1 => REG_17_27_port, A2 => n1601, B1 => 
                           REG_19_27_port, B2 => n1599, ZN => n1482);
   U2120 : AOI22_X1 port map( A1 => REG_20_27_port, A2 => n1610, B1 => 
                           REG_22_27_port, B2 => n1608, ZN => n1481);
   U2121 : AOI22_X1 port map( A1 => REG_16_27_port, A2 => n1612, B1 => 
                           REG_18_27_port, B2 => n8, ZN => n1480);
   U2122 : AND4_X1 port map( A1 => n1483, A2 => n1482, A3 => n1481, A4 => n1480
                           , ZN => n1500);
   U2123 : AOI22_X1 port map( A1 => REG_29_27_port, A2 => n1598, B1 => 
                           REG_31_27_port, B2 => n1595, ZN => n1487);
   U2124 : AOI22_X1 port map( A1 => REG_25_27_port, A2 => n1601, B1 => 
                           REG_27_27_port, B2 => n1599, ZN => n1486);
   U2125 : AOI22_X1 port map( A1 => REG_28_27_port, A2 => n1610, B1 => 
                           REG_30_27_port, B2 => n1608, ZN => n1485);
   U2126 : AOI22_X1 port map( A1 => REG_24_27_port, A2 => n1612, B1 => 
                           REG_26_27_port, B2 => n8, ZN => n1484);
   U2127 : AND4_X1 port map( A1 => n1487, A2 => n1486, A3 => n1485, A4 => n1484
                           , ZN => n1499);
   U2128 : AOI22_X1 port map( A1 => REG_5_27_port, A2 => n1598, B1 => 
                           REG_7_27_port, B2 => n1595, ZN => n1491);
   U2129 : AOI22_X1 port map( A1 => REG_1_27_port, A2 => n1601, B1 => 
                           REG_3_27_port, B2 => n1599, ZN => n1490);
   U2130 : AOI22_X1 port map( A1 => REG_4_27_port, A2 => n1610, B1 => 
                           REG_6_27_port, B2 => n1607, ZN => n1489);
   U2131 : AOI22_X1 port map( A1 => REG_0_27_port, A2 => n1612, B1 => 
                           REG_2_27_port, B2 => n8, ZN => n1488);
   U2132 : NAND4_X1 port map( A1 => n1491, A2 => n1490, A3 => n1489, A4 => 
                           n1488, ZN => n1497);
   U2133 : AOI22_X1 port map( A1 => REG_13_27_port, A2 => n1598, B1 => 
                           REG_15_27_port, B2 => n1595, ZN => n1495);
   U2134 : AOI22_X1 port map( A1 => REG_9_27_port, A2 => n1601, B1 => 
                           REG_11_27_port, B2 => n1599, ZN => n1494);
   U2135 : AOI22_X1 port map( A1 => REG_12_27_port, A2 => n1610, B1 => 
                           REG_14_27_port, B2 => n1607, ZN => n1493);
   U2136 : AOI22_X1 port map( A1 => REG_8_27_port, A2 => n1612, B1 => 
                           REG_10_27_port, B2 => n8, ZN => n1492);
   U2137 : NAND4_X1 port map( A1 => n1495, A2 => n1494, A3 => n1493, A4 => 
                           n1492, ZN => n1496);
   U2138 : AOI22_X1 port map( A1 => n1497, A2 => n1619, B1 => n1496, B2 => 
                           n1581, ZN => n1498);
   U2139 : OAI221_X1 port map( B1 => n1587, B2 => n1500, C1 => n1585, C2 => 
                           n1499, A => n1498, ZN => N288);
   U2140 : AOI22_X1 port map( A1 => REG_21_28_port, A2 => n1598, B1 => 
                           REG_23_28_port, B2 => n1595, ZN => n1504);
   U2141 : AOI22_X1 port map( A1 => REG_17_28_port, A2 => n1601, B1 => 
                           REG_19_28_port, B2 => n1599, ZN => n1503);
   U2142 : AOI22_X1 port map( A1 => REG_20_28_port, A2 => n1610, B1 => 
                           REG_22_28_port, B2 => n1607, ZN => n1502);
   U2143 : AOI22_X1 port map( A1 => REG_16_28_port, A2 => n1612, B1 => 
                           REG_18_28_port, B2 => n8, ZN => n1501);
   U2144 : AND4_X1 port map( A1 => n1504, A2 => n1503, A3 => n1502, A4 => n1501
                           , ZN => n1521);
   U2145 : AOI22_X1 port map( A1 => REG_29_28_port, A2 => n1598, B1 => 
                           REG_31_28_port, B2 => n1595, ZN => n1508);
   U2146 : AOI22_X1 port map( A1 => REG_25_28_port, A2 => n1601, B1 => 
                           REG_27_28_port, B2 => n1599, ZN => n1507);
   U2147 : AOI22_X1 port map( A1 => REG_28_28_port, A2 => n1610, B1 => 
                           REG_30_28_port, B2 => n1607, ZN => n1506);
   U2148 : AOI22_X1 port map( A1 => REG_24_28_port, A2 => n1612, B1 => 
                           REG_26_28_port, B2 => n8, ZN => n1505);
   U2149 : AND4_X1 port map( A1 => n1508, A2 => n1507, A3 => n1506, A4 => n1505
                           , ZN => n1520);
   U2150 : AOI22_X1 port map( A1 => REG_5_28_port, A2 => n1598, B1 => 
                           REG_7_28_port, B2 => n1595, ZN => n1512);
   U2151 : AOI22_X1 port map( A1 => REG_1_28_port, A2 => n1601, B1 => 
                           REG_3_28_port, B2 => n1599, ZN => n1511);
   U2152 : AOI22_X1 port map( A1 => REG_4_28_port, A2 => n1610, B1 => 
                           REG_6_28_port, B2 => n1607, ZN => n1510);
   U2153 : AOI22_X1 port map( A1 => REG_0_28_port, A2 => n1612, B1 => 
                           REG_2_28_port, B2 => n8, ZN => n1509);
   U2154 : NAND4_X1 port map( A1 => n1512, A2 => n1511, A3 => n1510, A4 => 
                           n1509, ZN => n1518);
   U2155 : AOI22_X1 port map( A1 => REG_13_28_port, A2 => n1598, B1 => 
                           REG_15_28_port, B2 => n1595, ZN => n1516);
   U2156 : AOI22_X1 port map( A1 => REG_9_28_port, A2 => n1601, B1 => 
                           REG_11_28_port, B2 => n1599, ZN => n1515);
   U2157 : AOI22_X1 port map( A1 => REG_12_28_port, A2 => n1610, B1 => 
                           REG_14_28_port, B2 => n1607, ZN => n1514);
   U2158 : AOI22_X1 port map( A1 => REG_8_28_port, A2 => n1612, B1 => 
                           REG_10_28_port, B2 => n8, ZN => n1513);
   U2159 : NAND4_X1 port map( A1 => n1516, A2 => n1515, A3 => n1514, A4 => 
                           n1513, ZN => n1517);
   U2160 : AOI22_X1 port map( A1 => n1518, A2 => n1619, B1 => n1517, B2 => 
                           n1581, ZN => n1519);
   U2161 : OAI221_X1 port map( B1 => n1587, B2 => n1521, C1 => n1585, C2 => 
                           n1520, A => n1519, ZN => N287);
   U2162 : AOI22_X1 port map( A1 => REG_21_29_port, A2 => n1598, B1 => 
                           REG_23_29_port, B2 => n1595, ZN => n1525);
   U2163 : AOI22_X1 port map( A1 => REG_17_29_port, A2 => n1601, B1 => 
                           REG_19_29_port, B2 => n1599, ZN => n1524);
   U2164 : AOI22_X1 port map( A1 => REG_20_29_port, A2 => n1610, B1 => 
                           REG_22_29_port, B2 => n1607, ZN => n1523);
   U2165 : AOI22_X1 port map( A1 => REG_16_29_port, A2 => n1612, B1 => 
                           REG_18_29_port, B2 => n8, ZN => n1522);
   U2166 : AND4_X1 port map( A1 => n1525, A2 => n1524, A3 => n1523, A4 => n1522
                           , ZN => n1542);
   U2167 : AOI22_X1 port map( A1 => REG_29_29_port, A2 => n1598, B1 => 
                           REG_31_29_port, B2 => n1595, ZN => n1529);
   U2168 : AOI22_X1 port map( A1 => REG_25_29_port, A2 => n1601, B1 => 
                           REG_27_29_port, B2 => n1599, ZN => n1528);
   U2169 : AOI22_X1 port map( A1 => REG_28_29_port, A2 => n1610, B1 => 
                           REG_30_29_port, B2 => n1607, ZN => n1527);
   U2170 : AOI22_X1 port map( A1 => REG_24_29_port, A2 => n1612, B1 => 
                           REG_26_29_port, B2 => n8, ZN => n1526);
   U2171 : AND4_X1 port map( A1 => n1529, A2 => n1528, A3 => n1527, A4 => n1526
                           , ZN => n1541);
   U2172 : AOI22_X1 port map( A1 => REG_5_29_port, A2 => n1598, B1 => 
                           REG_7_29_port, B2 => n1595, ZN => n1533);
   U2173 : AOI22_X1 port map( A1 => REG_1_29_port, A2 => n1601, B1 => 
                           REG_3_29_port, B2 => n1599, ZN => n1532);
   U2174 : AOI22_X1 port map( A1 => REG_4_29_port, A2 => n1610, B1 => 
                           REG_6_29_port, B2 => n1607, ZN => n1531);
   U2175 : AOI22_X1 port map( A1 => REG_0_29_port, A2 => n1612, B1 => 
                           REG_2_29_port, B2 => n8, ZN => n1530);
   U2176 : NAND4_X1 port map( A1 => n1533, A2 => n1532, A3 => n1531, A4 => 
                           n1530, ZN => n1539);
   U2177 : AOI22_X1 port map( A1 => REG_13_29_port, A2 => n1598, B1 => 
                           REG_15_29_port, B2 => n1595, ZN => n1537);
   U2178 : AOI22_X1 port map( A1 => REG_9_29_port, A2 => n1601, B1 => 
                           REG_11_29_port, B2 => n1599, ZN => n1536);
   U2179 : AOI22_X1 port map( A1 => REG_12_29_port, A2 => n1610, B1 => 
                           REG_14_29_port, B2 => n1607, ZN => n1535);
   U2180 : AOI22_X1 port map( A1 => REG_8_29_port, A2 => n1612, B1 => 
                           REG_10_29_port, B2 => n8, ZN => n1534);
   U2181 : NAND4_X1 port map( A1 => n1537, A2 => n1536, A3 => n1535, A4 => 
                           n1534, ZN => n1538);
   U2182 : AOI22_X1 port map( A1 => n1539, A2 => n1619, B1 => n1538, B2 => 
                           n1581, ZN => n1540);
   U2183 : OAI221_X1 port map( B1 => n1587, B2 => n1542, C1 => n1585, C2 => 
                           n1541, A => n1540, ZN => N286);
   U2184 : AOI22_X1 port map( A1 => REG_21_30_port, A2 => n1598, B1 => 
                           REG_23_30_port, B2 => n1595, ZN => n1546);
   U2185 : AOI22_X1 port map( A1 => REG_17_30_port, A2 => n1601, B1 => 
                           REG_19_30_port, B2 => n1599, ZN => n1545);
   U2186 : AOI22_X1 port map( A1 => REG_20_30_port, A2 => n1610, B1 => 
                           REG_22_30_port, B2 => n1607, ZN => n1544);
   U2187 : AOI22_X1 port map( A1 => REG_16_30_port, A2 => n1612, B1 => 
                           REG_18_30_port, B2 => n8, ZN => n1543);
   U2188 : AND4_X1 port map( A1 => n1546, A2 => n1545, A3 => n1544, A4 => n1543
                           , ZN => n1563);
   U2189 : AOI22_X1 port map( A1 => REG_29_30_port, A2 => n1598, B1 => 
                           REG_31_30_port, B2 => n1594, ZN => n1550);
   U2190 : AOI22_X1 port map( A1 => REG_25_30_port, A2 => n1601, B1 => 
                           REG_27_30_port, B2 => n1599, ZN => n1549);
   U2191 : AOI22_X1 port map( A1 => REG_28_30_port, A2 => n1610, B1 => 
                           REG_30_30_port, B2 => n1606, ZN => n1548);
   U2192 : AOI22_X1 port map( A1 => REG_24_30_port, A2 => n1613, B1 => 
                           REG_26_30_port, B2 => n8, ZN => n1547);
   U2193 : AND4_X1 port map( A1 => n1550, A2 => n1549, A3 => n1548, A4 => n1547
                           , ZN => n1562);
   U2194 : AOI22_X1 port map( A1 => REG_5_30_port, A2 => n1598, B1 => 
                           REG_7_30_port, B2 => n1594, ZN => n1554);
   U2195 : AOI22_X1 port map( A1 => REG_1_30_port, A2 => n1601, B1 => 
                           REG_3_30_port, B2 => n1599, ZN => n1553);
   U2196 : AOI22_X1 port map( A1 => REG_4_30_port, A2 => n1610, B1 => 
                           REG_6_30_port, B2 => n1606, ZN => n1552);
   U2197 : AOI22_X1 port map( A1 => REG_0_30_port, A2 => n1613, B1 => 
                           REG_2_30_port, B2 => n8, ZN => n1551);
   U2198 : NAND4_X1 port map( A1 => n1554, A2 => n1553, A3 => n1552, A4 => 
                           n1551, ZN => n1560);
   U2199 : AOI22_X1 port map( A1 => REG_13_30_port, A2 => n1598, B1 => 
                           REG_15_30_port, B2 => n1594, ZN => n1558);
   U2200 : AOI22_X1 port map( A1 => REG_9_30_port, A2 => n1601, B1 => 
                           REG_11_30_port, B2 => n1599, ZN => n1557);
   U2201 : AOI22_X1 port map( A1 => REG_12_30_port, A2 => n1610, B1 => 
                           REG_14_30_port, B2 => n1606, ZN => n1556);
   U2202 : AOI22_X1 port map( A1 => REG_8_30_port, A2 => n1613, B1 => 
                           REG_10_30_port, B2 => n8, ZN => n1555);
   U2203 : NAND4_X1 port map( A1 => n1558, A2 => n1557, A3 => n1556, A4 => 
                           n1555, ZN => n1559);
   U2204 : AOI22_X1 port map( A1 => n1560, A2 => n1619, B1 => n1559, B2 => 
                           n1581, ZN => n1561);
   U2205 : OAI221_X1 port map( B1 => n1587, B2 => n1563, C1 => n1585, C2 => 
                           n1562, A => n1561, ZN => N285);
   U2206 : AOI22_X1 port map( A1 => REG_21_31_port, A2 => n1598, B1 => 
                           REG_23_31_port, B2 => n1594, ZN => n1567);
   U2207 : AOI22_X1 port map( A1 => REG_17_31_port, A2 => n1601, B1 => 
                           REG_19_31_port, B2 => n1599, ZN => n1566);
   U2208 : AOI22_X1 port map( A1 => REG_20_31_port, A2 => n1610, B1 => 
                           REG_22_31_port, B2 => n1606, ZN => n1565);
   U2209 : AOI22_X1 port map( A1 => REG_16_31_port, A2 => n1613, B1 => 
                           REG_18_31_port, B2 => n8, ZN => n1564);
   U2210 : AND4_X1 port map( A1 => n1567, A2 => n1566, A3 => n1565, A4 => n1564
                           , ZN => n1588);
   U2211 : AOI22_X1 port map( A1 => REG_29_31_port, A2 => n1598, B1 => 
                           REG_31_31_port, B2 => n1594, ZN => n1571);
   U2212 : AOI22_X1 port map( A1 => REG_25_31_port, A2 => n1601, B1 => 
                           REG_27_31_port, B2 => n1599, ZN => n1570);
   U2213 : AOI22_X1 port map( A1 => REG_28_31_port, A2 => n1610, B1 => 
                           REG_30_31_port, B2 => n1606, ZN => n1569);
   U2214 : AOI22_X1 port map( A1 => REG_24_31_port, A2 => n1613, B1 => 
                           REG_26_31_port, B2 => n8, ZN => n1568);
   U2215 : AND4_X1 port map( A1 => n1571, A2 => n1570, A3 => n1569, A4 => n1568
                           , ZN => n1586);
   U2216 : AOI22_X1 port map( A1 => REG_5_31_port, A2 => n1598, B1 => 
                           REG_7_31_port, B2 => n1594, ZN => n1575);
   U2217 : AOI22_X1 port map( A1 => REG_1_31_port, A2 => n1601, B1 => 
                           REG_3_31_port, B2 => n1599, ZN => n1574);
   U2218 : AOI22_X1 port map( A1 => REG_4_31_port, A2 => n1610, B1 => 
                           REG_6_31_port, B2 => n1606, ZN => n1573);
   U2219 : AOI22_X1 port map( A1 => REG_0_31_port, A2 => n1613, B1 => 
                           REG_2_31_port, B2 => n8, ZN => n1572);
   U2220 : NAND4_X1 port map( A1 => n1575, A2 => n1574, A3 => n1573, A4 => 
                           n1572, ZN => n1582);
   U2221 : AOI22_X1 port map( A1 => REG_13_31_port, A2 => n1598, B1 => 
                           REG_15_31_port, B2 => n1594, ZN => n1579);
   U2222 : AOI22_X1 port map( A1 => REG_9_31_port, A2 => n1601, B1 => 
                           REG_11_31_port, B2 => n1599, ZN => n1578);
   U2223 : AOI22_X1 port map( A1 => REG_12_31_port, A2 => n1610, B1 => 
                           REG_14_31_port, B2 => n1606, ZN => n1577);
   U2224 : AOI22_X1 port map( A1 => REG_8_31_port, A2 => n1613, B1 => 
                           REG_10_31_port, B2 => n8, ZN => n1576);
   U2225 : NAND4_X1 port map( A1 => n1579, A2 => n1578, A3 => n1577, A4 => 
                           n1576, ZN => n1580);
   U2226 : AOI22_X1 port map( A1 => n1619, A2 => n1582, B1 => n1581, B2 => 
                           n1580, ZN => n1584);
   U2227 : OAI221_X1 port map( B1 => n1588, B2 => n1587, C1 => n1586, C2 => 
                           n1585, A => n1584, ZN => N284);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_6 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_6;

architecture SYN_STRUCTURAL of LDR_N32_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_192
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_193
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_194
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_195
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_196
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_197
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_198
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_199
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_200
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_201
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_202
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_203
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_204
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_205
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_206
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_207
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_208
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_209
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_210
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_211
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_212
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_213
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_214
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_215
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_216
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_217
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_218
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_219
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_220
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_221
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_222
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_223
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_223 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_222 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_221 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_220 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_219 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_218 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_217 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_216 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_215 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_214 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_213 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_212 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_211 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_210 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_209 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_208 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_207 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_206 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_205 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_204 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_203 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_202 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_201 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9))
                           ;
   LDI_8 : LD_200 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8))
                           ;
   LDI_7 : LD_199 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7))
                           ;
   LDI_6 : LD_198 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6))
                           ;
   LDI_5 : LD_197 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5))
                           ;
   LDI_4 : LD_196 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4))
                           ;
   LDI_3 : LD_195 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3))
                           ;
   LDI_2 : LD_194 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2))
                           ;
   LDI_1 : LD_193 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1))
                           ;
   LDI_0 : LD_192 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0))
                           ;
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_4;

architecture SYN_BEHAVIORAL of MUX21_N32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => S, Z => n6);
   U2 : BUF_X1 port map( A => S, Z => n7);
   U3 : BUF_X1 port map( A => n7, Z => n2);
   U4 : BUF_X1 port map( A => n7, Z => n1);
   U5 : INV_X1 port map( A => n6, ZN => n5);
   U6 : INV_X1 port map( A => n6, ZN => n4);
   U7 : BUF_X1 port map( A => n7, Z => n3);
   U8 : INV_X1 port map( A => n54, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n1, ZN => 
                           n54);
   U10 : INV_X1 port map( A => n65, ZN => Y(0));
   U11 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n1, ZN => 
                           n65);
   U12 : INV_X1 port map( A => n43, ZN => Y(2));
   U13 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n2, ZN => 
                           n43);
   U14 : INV_X1 port map( A => n40, ZN => Y(3));
   U15 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => B(3), B2 => n3, ZN => 
                           n40);
   U16 : INV_X1 port map( A => n42, ZN => Y(30));
   U17 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n2, ZN =>
                           n42);
   U18 : INV_X1 port map( A => n44, ZN => Y(29));
   U19 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n2, ZN =>
                           n44);
   U20 : INV_X1 port map( A => n45, ZN => Y(28));
   U21 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n2, ZN =>
                           n45);
   U22 : INV_X1 port map( A => n46, ZN => Y(27));
   U23 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n2, ZN =>
                           n46);
   U24 : INV_X1 port map( A => n47, ZN => Y(26));
   U25 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n2, ZN =>
                           n47);
   U26 : INV_X1 port map( A => n48, ZN => Y(25));
   U27 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n2, ZN =>
                           n48);
   U28 : INV_X1 port map( A => n49, ZN => Y(24));
   U29 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n2, ZN =>
                           n49);
   U30 : INV_X1 port map( A => n50, ZN => Y(23));
   U31 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n2, ZN =>
                           n50);
   U32 : INV_X1 port map( A => n51, ZN => Y(22));
   U33 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n2, ZN =>
                           n51);
   U34 : INV_X1 port map( A => n52, ZN => Y(21));
   U35 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n2, ZN =>
                           n52);
   U36 : INV_X1 port map( A => n53, ZN => Y(20));
   U37 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n2, ZN =>
                           n53);
   U38 : INV_X1 port map( A => n55, ZN => Y(19));
   U39 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n1, ZN =>
                           n55);
   U40 : INV_X1 port map( A => n56, ZN => Y(18));
   U41 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n1, ZN =>
                           n56);
   U42 : INV_X1 port map( A => n57, ZN => Y(17));
   U43 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n1, ZN =>
                           n57);
   U44 : INV_X1 port map( A => n58, ZN => Y(16));
   U45 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n1, ZN =>
                           n58);
   U46 : INV_X1 port map( A => n59, ZN => Y(15));
   U47 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n1, ZN =>
                           n59);
   U48 : INV_X1 port map( A => n60, ZN => Y(14));
   U49 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n1, ZN =>
                           n60);
   U50 : INV_X1 port map( A => n61, ZN => Y(13));
   U51 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n1, ZN =>
                           n61);
   U52 : INV_X1 port map( A => n62, ZN => Y(12));
   U53 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n1, ZN =>
                           n62);
   U54 : INV_X1 port map( A => n63, ZN => Y(11));
   U55 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n1, ZN =>
                           n63);
   U56 : INV_X1 port map( A => n64, ZN => Y(10));
   U57 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n1, ZN =>
                           n64);
   U58 : INV_X1 port map( A => n35, ZN => Y(8));
   U59 : AOI22_X1 port map( A1 => A(8), A2 => n4, B1 => B(8), B2 => n3, ZN => 
                           n35);
   U60 : INV_X1 port map( A => n36, ZN => Y(7));
   U61 : AOI22_X1 port map( A1 => A(7), A2 => n5, B1 => B(7), B2 => n3, ZN => 
                           n36);
   U62 : INV_X1 port map( A => n37, ZN => Y(6));
   U63 : AOI22_X1 port map( A1 => A(6), A2 => n4, B1 => B(6), B2 => n3, ZN => 
                           n37);
   U64 : INV_X1 port map( A => n38, ZN => Y(5));
   U65 : AOI22_X1 port map( A1 => A(5), A2 => n5, B1 => B(5), B2 => n3, ZN => 
                           n38);
   U66 : INV_X1 port map( A => n39, ZN => Y(4));
   U67 : AOI22_X1 port map( A1 => A(4), A2 => n4, B1 => B(4), B2 => n3, ZN => 
                           n39);
   U68 : INV_X1 port map( A => n41, ZN => Y(31));
   U69 : AOI22_X1 port map( A1 => A(31), A2 => n5, B1 => B(31), B2 => n3, ZN =>
                           n41);
   U70 : INV_X1 port map( A => n34, ZN => Y(9));
   U71 : AOI22_X1 port map( A1 => A(9), A2 => n4, B1 => n3, B2 => B(9), ZN => 
                           n34);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFDR_N32 is

   port( CLK, RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 
         0);  REGOUT : out std_logic_vector (31 downto 0));

end FFDR_N32;

architecture SYN_STRUCTURAL of FFDR_N32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FFD_0
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_1
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_2
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_3
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_4
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_5
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_6
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_7
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_8
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_9
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_10
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_11
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_12
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_13
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_14
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_15
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_16
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_17
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_18
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_19
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_20
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_21
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_22
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_23
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_24
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_25
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_26
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_27
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_28
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_29
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_30
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_31
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   FFI_31 : FFD_31 port map( CLK => CLK, RST => n3, EN => EN, D => REGIN(31), Q
                           => REGOUT(31));
   FFI_30 : FFD_30 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(30), Q
                           => REGOUT(30));
   FFI_29 : FFD_29 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(29), Q
                           => REGOUT(29));
   FFI_28 : FFD_28 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(28), Q
                           => REGOUT(28));
   FFI_27 : FFD_27 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(27), Q
                           => REGOUT(27));
   FFI_26 : FFD_26 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(26), Q
                           => REGOUT(26));
   FFI_25 : FFD_25 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(25), Q
                           => REGOUT(25));
   FFI_24 : FFD_24 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(24), Q
                           => REGOUT(24));
   FFI_23 : FFD_23 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(23), Q
                           => REGOUT(23));
   FFI_22 : FFD_22 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(22), Q
                           => REGOUT(22));
   FFI_21 : FFD_21 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(21), Q
                           => REGOUT(21));
   FFI_20 : FFD_20 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(20), Q
                           => REGOUT(20));
   FFI_19 : FFD_19 port map( CLK => CLK, RST => n1, EN => EN, D => REGIN(19), Q
                           => REGOUT(19));
   FFI_18 : FFD_18 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(18), Q
                           => REGOUT(18));
   FFI_17 : FFD_17 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(17), Q
                           => REGOUT(17));
   FFI_16 : FFD_16 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(16), Q
                           => REGOUT(16));
   FFI_15 : FFD_15 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(15), Q
                           => REGOUT(15));
   FFI_14 : FFD_14 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(14), Q
                           => REGOUT(14));
   FFI_13 : FFD_13 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(13), Q
                           => REGOUT(13));
   FFI_12 : FFD_12 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(12), Q
                           => REGOUT(12));
   FFI_11 : FFD_11 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(11), Q
                           => REGOUT(11));
   FFI_10 : FFD_10 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(10), Q
                           => REGOUT(10));
   FFI_9 : FFD_9 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(9), Q =>
                           REGOUT(9));
   FFI_8 : FFD_8 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(8), Q =>
                           REGOUT(8));
   FFI_7 : FFD_7 port map( CLK => CLK, RST => n2, EN => EN, D => REGIN(7), Q =>
                           REGOUT(7));
   FFI_6 : FFD_6 port map( CLK => CLK, RST => n3, EN => EN, D => REGIN(6), Q =>
                           REGOUT(6));
   FFI_5 : FFD_5 port map( CLK => CLK, RST => n3, EN => EN, D => REGIN(5), Q =>
                           REGOUT(5));
   FFI_4 : FFD_4 port map( CLK => CLK, RST => n3, EN => EN, D => REGIN(4), Q =>
                           REGOUT(4));
   FFI_3 : FFD_3 port map( CLK => CLK, RST => n3, EN => EN, D => REGIN(3), Q =>
                           REGOUT(3));
   FFI_2 : FFD_2 port map( CLK => CLK, RST => n3, EN => EN, D => REGIN(2), Q =>
                           REGOUT(2));
   FFI_1 : FFD_1 port map( CLK => CLK, RST => n3, EN => EN, D => REGIN(1), Q =>
                           REGOUT(1));
   FFI_0 : FFD_0 port map( CLK => CLK, RST => n3, EN => EN, D => REGIN(0), Q =>
                           REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32 is

   port( CLK, RST : in std_logic;  IR_IN, DRAM_OUT : in std_logic_vector (31 
         downto 0);  IR_LATCH_EN, PC_LATCH_EN, NPC_LATCH_EN, RF_WE, 
         RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, 
         ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
         std_logic_vector (0 to 6);  LMD_LATCH_EN, JUMP_EN, JUMP_COND, 
         WB_MUX_SEL, JAL_MUX_SEL : in std_logic;  IR_OUT, PC_OUT, ALU_OUT, 
         DRAM_IN : out std_logic_vector (31 downto 0));

end DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32;

architecture SYN_DLX_DATAPATH_ARCH of 
   DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component 
      DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component MUX21_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component LDR_N32_0
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component LD_224
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LDR_N32_1
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component FU_N5
      port( RS1, RS2, RD_MEM, RD_WB : in std_logic_vector (4 downto 0);  
            RF_WE_MEM, RF_WE_WB : in std_logic;  FORWARD_A, FORWARD_B : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component ZERO_DETECTOR_N32_1
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic);
   end component;
   
   component MUX21_L_320
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component ALU_N32_NB8
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
            std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);
            Z : out std_logic);
   end component;
   
   component MUX21_N32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_N32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX41_N32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX41_N32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component LDR_N32_2
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component LDR_N32_3
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component LDR_N32_4
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REGADDR_N32_OPC6_REG5
      port( INSTR : in std_logic_vector (31 downto 0);  RS1, RS2, RD : out 
            std_logic_vector (4 downto 0));
   end component;
   
   component SIGNEX_N32_OPC6_REG5
      port( INSTR : in std_logic_vector (31 downto 0);  IMM : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component RF_N32_NA5
      port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
            ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component LDR_N32_5
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component LDR_N32_6
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_N32_4
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component FFDR_N32
      port( CLK, RST, EN : in std_logic;  REGIN : in std_logic_vector (31 
            downto 0);  REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, IR_OUT_31_port, IR_OUT_30_port, 
      IR_OUT_29_port, IR_OUT_28_port, IR_OUT_27_port, IR_OUT_26_port, 
      IR_OUT_25_port, IR_OUT_24_port, IR_OUT_23_port, IR_OUT_22_port, 
      IR_OUT_21_port, IR_OUT_20_port, IR_OUT_19_port, IR_OUT_18_port, 
      IR_OUT_17_port, IR_OUT_16_port, IR_OUT_15_port, IR_OUT_14_port, 
      IR_OUT_13_port, IR_OUT_12_port, IR_OUT_11_port, IR_OUT_10_port, 
      IR_OUT_9_port, IR_OUT_8_port, IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port
      , IR_OUT_4_port, IR_OUT_3_port, IR_OUT_2_port, IR_OUT_1_port, 
      IR_OUT_0_port, PC_OUT_31_port, PC_OUT_30_port, PC_OUT_29_port, 
      PC_OUT_28_port, PC_OUT_27_port, PC_OUT_26_port, PC_OUT_25_port, 
      PC_OUT_24_port, PC_OUT_23_port, PC_OUT_22_port, PC_OUT_21_port, 
      PC_OUT_20_port, PC_OUT_19_port, PC_OUT_18_port, PC_OUT_17_port, 
      PC_OUT_16_port, PC_OUT_15_port, PC_OUT_14_port, PC_OUT_13_port, 
      PC_OUT_12_port, PC_OUT_11_port, PC_OUT_10_port, PC_OUT_9_port, 
      PC_OUT_8_port, PC_OUT_7_port, PC_OUT_6_port, PC_OUT_5_port, PC_OUT_4_port
      , PC_OUT_3_port, PC_OUT_2_port, PC_OUT_1_port, PC_OUT_0_port, 
      ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, ALU_OUT_28_port, 
      ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, ALU_OUT_24_port, 
      ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, ALU_OUT_20_port, 
      ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, ALU_OUT_16_port, 
      ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, ALU_OUT_12_port, 
      ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, ALU_OUT_8_port, 
      ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, ALU_OUT_4_port, 
      ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, ALU_OUT_0_port, 
      IF_ID_NPC_31_port, IF_ID_NPC_30_port, IF_ID_NPC_29_port, 
      IF_ID_NPC_28_port, IF_ID_NPC_27_port, IF_ID_NPC_26_port, 
      IF_ID_NPC_25_port, IF_ID_NPC_24_port, IF_ID_NPC_23_port, 
      IF_ID_NPC_22_port, IF_ID_NPC_21_port, IF_ID_NPC_20_port, 
      IF_ID_NPC_19_port, IF_ID_NPC_18_port, IF_ID_NPC_17_port, 
      IF_ID_NPC_16_port, IF_ID_NPC_15_port, IF_ID_NPC_14_port, 
      IF_ID_NPC_13_port, IF_ID_NPC_12_port, IF_ID_NPC_11_port, 
      IF_ID_NPC_10_port, IF_ID_NPC_9_port, IF_ID_NPC_8_port, IF_ID_NPC_7_port, 
      IF_ID_NPC_6_port, IF_ID_NPC_5_port, IF_ID_NPC_4_port, IF_ID_NPC_3_port, 
      IF_ID_NPC_2_port, IF_ID_NPC_1_port, IF_ID_NPC_0_port, IF_ID_IR_31_port, 
      IF_ID_IR_30_port, IF_ID_IR_29_port, IF_ID_IR_28_port, IF_ID_IR_27_port, 
      IF_ID_IR_26_port, IF_ID_IR_25_port, IF_ID_IR_24_port, IF_ID_IR_23_port, 
      IF_ID_IR_22_port, IF_ID_IR_21_port, IF_ID_IR_20_port, IF_ID_IR_19_port, 
      IF_ID_IR_18_port, IF_ID_IR_17_port, IF_ID_IR_16_port, IF_ID_IR_15_port, 
      IF_ID_IR_14_port, IF_ID_IR_13_port, IF_ID_IR_12_port, IF_ID_IR_11_port, 
      IF_ID_IR_10_port, IF_ID_IR_9_port, IF_ID_IR_8_port, IF_ID_IR_7_port, 
      IF_ID_IR_6_port, IF_ID_IR_5_port, IF_ID_IR_4_port, IF_ID_IR_3_port, 
      IF_ID_IR_2_port, IF_ID_IR_1_port, IF_ID_IR_0_port, ID_EX_NPC_31_port, 
      ID_EX_NPC_30_port, ID_EX_NPC_29_port, ID_EX_NPC_28_port, 
      ID_EX_NPC_27_port, ID_EX_NPC_26_port, ID_EX_NPC_25_port, 
      ID_EX_NPC_24_port, ID_EX_NPC_23_port, ID_EX_NPC_22_port, 
      ID_EX_NPC_21_port, ID_EX_NPC_20_port, ID_EX_NPC_19_port, 
      ID_EX_NPC_18_port, ID_EX_NPC_17_port, ID_EX_NPC_16_port, 
      ID_EX_NPC_15_port, ID_EX_NPC_14_port, ID_EX_NPC_13_port, 
      ID_EX_NPC_12_port, ID_EX_NPC_11_port, ID_EX_NPC_10_port, ID_EX_NPC_9_port
      , ID_EX_NPC_8_port, ID_EX_NPC_7_port, ID_EX_NPC_6_port, ID_EX_NPC_5_port,
      ID_EX_NPC_4_port, ID_EX_NPC_3_port, ID_EX_NPC_2_port, ID_EX_NPC_1_port, 
      ID_EX_NPC_0_port, ID_EX_RF_WE, ID_EX_RS1_4_port, ID_EX_RS1_3_port, 
      ID_EX_RS1_2_port, ID_EX_RS1_1_port, ID_EX_RS1_0_port, ID_EX_RS2_4_port, 
      ID_EX_RS2_3_port, ID_EX_RS2_2_port, ID_EX_RS2_1_port, ID_EX_RS2_0_port, 
      ID_EX_RD_4_port, ID_EX_RD_3_port, ID_EX_RD_2_port, ID_EX_RD_1_port, 
      ID_EX_RD_0_port, ID_EX_RF_OUT1_31_port, ID_EX_RF_OUT1_30_port, 
      ID_EX_RF_OUT1_29_port, ID_EX_RF_OUT1_28_port, ID_EX_RF_OUT1_27_port, 
      ID_EX_RF_OUT1_26_port, ID_EX_RF_OUT1_25_port, ID_EX_RF_OUT1_24_port, 
      ID_EX_RF_OUT1_23_port, ID_EX_RF_OUT1_22_port, ID_EX_RF_OUT1_21_port, 
      ID_EX_RF_OUT1_20_port, ID_EX_RF_OUT1_19_port, ID_EX_RF_OUT1_18_port, 
      ID_EX_RF_OUT1_17_port, ID_EX_RF_OUT1_16_port, ID_EX_RF_OUT1_15_port, 
      ID_EX_RF_OUT1_14_port, ID_EX_RF_OUT1_13_port, ID_EX_RF_OUT1_12_port, 
      ID_EX_RF_OUT1_11_port, ID_EX_RF_OUT1_10_port, ID_EX_RF_OUT1_9_port, 
      ID_EX_RF_OUT1_8_port, ID_EX_RF_OUT1_7_port, ID_EX_RF_OUT1_6_port, 
      ID_EX_RF_OUT1_5_port, ID_EX_RF_OUT1_4_port, ID_EX_RF_OUT1_3_port, 
      ID_EX_RF_OUT1_2_port, ID_EX_RF_OUT1_1_port, ID_EX_RF_OUT1_0_port, 
      ID_EX_RF_OUT2_31_port, ID_EX_RF_OUT2_30_port, ID_EX_RF_OUT2_29_port, 
      ID_EX_RF_OUT2_28_port, ID_EX_RF_OUT2_27_port, ID_EX_RF_OUT2_26_port, 
      ID_EX_RF_OUT2_25_port, ID_EX_RF_OUT2_24_port, ID_EX_RF_OUT2_23_port, 
      ID_EX_RF_OUT2_22_port, ID_EX_RF_OUT2_21_port, ID_EX_RF_OUT2_20_port, 
      ID_EX_RF_OUT2_19_port, ID_EX_RF_OUT2_18_port, ID_EX_RF_OUT2_17_port, 
      ID_EX_RF_OUT2_16_port, ID_EX_RF_OUT2_15_port, ID_EX_RF_OUT2_14_port, 
      ID_EX_RF_OUT2_13_port, ID_EX_RF_OUT2_12_port, ID_EX_RF_OUT2_11_port, 
      ID_EX_RF_OUT2_10_port, ID_EX_RF_OUT2_9_port, ID_EX_RF_OUT2_8_port, 
      ID_EX_RF_OUT2_7_port, ID_EX_RF_OUT2_6_port, ID_EX_RF_OUT2_5_port, 
      ID_EX_RF_OUT2_4_port, ID_EX_RF_OUT2_3_port, ID_EX_RF_OUT2_2_port, 
      ID_EX_RF_OUT2_1_port, ID_EX_RF_OUT2_0_port, ID_EX_IMM_31_port, 
      ID_EX_IMM_30_port, ID_EX_IMM_29_port, ID_EX_IMM_28_port, 
      ID_EX_IMM_27_port, ID_EX_IMM_26_port, ID_EX_IMM_25_port, 
      ID_EX_IMM_24_port, ID_EX_IMM_23_port, ID_EX_IMM_22_port, 
      ID_EX_IMM_21_port, ID_EX_IMM_20_port, ID_EX_IMM_19_port, 
      ID_EX_IMM_18_port, ID_EX_IMM_17_port, ID_EX_IMM_16_port, 
      ID_EX_IMM_15_port, ID_EX_IMM_14_port, ID_EX_IMM_13_port, 
      ID_EX_IMM_12_port, ID_EX_IMM_11_port, ID_EX_IMM_10_port, ID_EX_IMM_9_port
      , ID_EX_IMM_8_port, ID_EX_IMM_7_port, ID_EX_IMM_6_port, ID_EX_IMM_5_port,
      ID_EX_IMM_4_port, ID_EX_IMM_3_port, ID_EX_IMM_2_port, ID_EX_IMM_1_port, 
      ID_EX_IMM_0_port, EX_MEM_NPC_31_port, EX_MEM_NPC_30_port, 
      EX_MEM_NPC_29_port, EX_MEM_NPC_28_port, EX_MEM_NPC_27_port, 
      EX_MEM_NPC_26_port, EX_MEM_NPC_25_port, EX_MEM_NPC_24_port, 
      EX_MEM_NPC_23_port, EX_MEM_NPC_22_port, EX_MEM_NPC_21_port, 
      EX_MEM_NPC_20_port, EX_MEM_NPC_19_port, EX_MEM_NPC_18_port, 
      EX_MEM_NPC_17_port, EX_MEM_NPC_16_port, EX_MEM_NPC_15_port, 
      EX_MEM_NPC_14_port, EX_MEM_NPC_13_port, EX_MEM_NPC_12_port, 
      EX_MEM_NPC_11_port, EX_MEM_NPC_10_port, EX_MEM_NPC_9_port, 
      EX_MEM_NPC_8_port, EX_MEM_NPC_7_port, EX_MEM_NPC_6_port, 
      EX_MEM_NPC_5_port, EX_MEM_NPC_4_port, EX_MEM_NPC_3_port, 
      EX_MEM_NPC_2_port, EX_MEM_NPC_1_port, EX_MEM_NPC_0_port, EX_MEM_RF_WE, 
      EX_MEM_BRANCH_DETECT, EX_MEM_RD_4_port, EX_MEM_RD_3_port, 
      EX_MEM_RD_2_port, EX_MEM_RD_1_port, EX_MEM_RD_0_port, MEM_WB_NPC_31_port,
      MEM_WB_NPC_30_port, MEM_WB_NPC_29_port, MEM_WB_NPC_28_port, 
      MEM_WB_NPC_27_port, MEM_WB_NPC_26_port, MEM_WB_NPC_25_port, 
      MEM_WB_NPC_24_port, MEM_WB_NPC_23_port, MEM_WB_NPC_22_port, 
      MEM_WB_NPC_21_port, MEM_WB_NPC_20_port, MEM_WB_NPC_19_port, 
      MEM_WB_NPC_18_port, MEM_WB_NPC_17_port, MEM_WB_NPC_16_port, 
      MEM_WB_NPC_15_port, MEM_WB_NPC_14_port, MEM_WB_NPC_13_port, 
      MEM_WB_NPC_12_port, MEM_WB_NPC_11_port, MEM_WB_NPC_10_port, 
      MEM_WB_NPC_9_port, MEM_WB_NPC_8_port, MEM_WB_NPC_7_port, 
      MEM_WB_NPC_6_port, MEM_WB_NPC_5_port, MEM_WB_NPC_4_port, 
      MEM_WB_NPC_3_port, MEM_WB_NPC_2_port, MEM_WB_NPC_1_port, 
      MEM_WB_NPC_0_port, MEM_WB_RF_WE, MEM_WB_ALU_OUTPUT_31_port, 
      MEM_WB_ALU_OUTPUT_30_port, MEM_WB_ALU_OUTPUT_29_port, 
      MEM_WB_ALU_OUTPUT_28_port, MEM_WB_ALU_OUTPUT_27_port, 
      MEM_WB_ALU_OUTPUT_26_port, MEM_WB_ALU_OUTPUT_25_port, 
      MEM_WB_ALU_OUTPUT_24_port, MEM_WB_ALU_OUTPUT_23_port, 
      MEM_WB_ALU_OUTPUT_22_port, MEM_WB_ALU_OUTPUT_21_port, 
      MEM_WB_ALU_OUTPUT_20_port, MEM_WB_ALU_OUTPUT_19_port, 
      MEM_WB_ALU_OUTPUT_18_port, MEM_WB_ALU_OUTPUT_17_port, 
      MEM_WB_ALU_OUTPUT_16_port, MEM_WB_ALU_OUTPUT_15_port, 
      MEM_WB_ALU_OUTPUT_14_port, MEM_WB_ALU_OUTPUT_13_port, 
      MEM_WB_ALU_OUTPUT_12_port, MEM_WB_ALU_OUTPUT_11_port, 
      MEM_WB_ALU_OUTPUT_10_port, MEM_WB_ALU_OUTPUT_9_port, 
      MEM_WB_ALU_OUTPUT_8_port, MEM_WB_ALU_OUTPUT_7_port, 
      MEM_WB_ALU_OUTPUT_6_port, MEM_WB_ALU_OUTPUT_5_port, 
      MEM_WB_ALU_OUTPUT_4_port, MEM_WB_ALU_OUTPUT_3_port, 
      MEM_WB_ALU_OUTPUT_2_port, MEM_WB_ALU_OUTPUT_1_port, 
      MEM_WB_ALU_OUTPUT_0_port, MEM_WB_DRAM_OUTPUT_31_port, 
      MEM_WB_DRAM_OUTPUT_30_port, MEM_WB_DRAM_OUTPUT_29_port, 
      MEM_WB_DRAM_OUTPUT_28_port, MEM_WB_DRAM_OUTPUT_27_port, 
      MEM_WB_DRAM_OUTPUT_26_port, MEM_WB_DRAM_OUTPUT_25_port, 
      MEM_WB_DRAM_OUTPUT_24_port, MEM_WB_DRAM_OUTPUT_23_port, 
      MEM_WB_DRAM_OUTPUT_22_port, MEM_WB_DRAM_OUTPUT_21_port, 
      MEM_WB_DRAM_OUTPUT_20_port, MEM_WB_DRAM_OUTPUT_19_port, 
      MEM_WB_DRAM_OUTPUT_18_port, MEM_WB_DRAM_OUTPUT_17_port, 
      MEM_WB_DRAM_OUTPUT_16_port, MEM_WB_DRAM_OUTPUT_15_port, 
      MEM_WB_DRAM_OUTPUT_14_port, MEM_WB_DRAM_OUTPUT_13_port, 
      MEM_WB_DRAM_OUTPUT_12_port, MEM_WB_DRAM_OUTPUT_11_port, 
      MEM_WB_DRAM_OUTPUT_10_port, MEM_WB_DRAM_OUTPUT_9_port, 
      MEM_WB_DRAM_OUTPUT_8_port, MEM_WB_DRAM_OUTPUT_7_port, 
      MEM_WB_DRAM_OUTPUT_6_port, MEM_WB_DRAM_OUTPUT_5_port, 
      MEM_WB_DRAM_OUTPUT_4_port, MEM_WB_DRAM_OUTPUT_3_port, 
      MEM_WB_DRAM_OUTPUT_2_port, MEM_WB_DRAM_OUTPUT_1_port, 
      MEM_WB_DRAM_OUTPUT_0_port, MEM_WB_RD_4_port, MEM_WB_RD_3_port, 
      MEM_WB_RD_2_port, MEM_WB_RD_1_port, MEM_WB_RD_0_port, 
      IF_ID_NPC_NEXT_31_port, IF_ID_NPC_NEXT_30_port, IF_ID_NPC_NEXT_29_port, 
      IF_ID_NPC_NEXT_28_port, IF_ID_NPC_NEXT_27_port, IF_ID_NPC_NEXT_26_port, 
      IF_ID_NPC_NEXT_25_port, IF_ID_NPC_NEXT_24_port, IF_ID_NPC_NEXT_23_port, 
      IF_ID_NPC_NEXT_22_port, IF_ID_NPC_NEXT_21_port, IF_ID_NPC_NEXT_20_port, 
      IF_ID_NPC_NEXT_19_port, IF_ID_NPC_NEXT_18_port, IF_ID_NPC_NEXT_17_port, 
      IF_ID_NPC_NEXT_16_port, IF_ID_NPC_NEXT_15_port, IF_ID_NPC_NEXT_14_port, 
      IF_ID_NPC_NEXT_13_port, IF_ID_NPC_NEXT_12_port, IF_ID_NPC_NEXT_11_port, 
      IF_ID_NPC_NEXT_10_port, IF_ID_NPC_NEXT_9_port, IF_ID_NPC_NEXT_8_port, 
      IF_ID_NPC_NEXT_7_port, IF_ID_NPC_NEXT_6_port, IF_ID_NPC_NEXT_5_port, 
      IF_ID_NPC_NEXT_4_port, IF_ID_NPC_NEXT_3_port, IF_ID_NPC_NEXT_2_port, 
      IF_ID_NPC_NEXT_1_port, IF_ID_NPC_NEXT_0_port, ID_EX_RS1_NEXT_4_port, 
      ID_EX_RS1_NEXT_3_port, ID_EX_RS1_NEXT_2_port, ID_EX_RS1_NEXT_1_port, 
      ID_EX_RS1_NEXT_0_port, ID_EX_RS2_NEXT_4_port, ID_EX_RS2_NEXT_3_port, 
      ID_EX_RS2_NEXT_2_port, ID_EX_RS2_NEXT_1_port, ID_EX_RS2_NEXT_0_port, 
      ID_EX_RD_NEXT_4_port, ID_EX_RD_NEXT_3_port, ID_EX_RD_NEXT_2_port, 
      ID_EX_RD_NEXT_1_port, ID_EX_RD_NEXT_0_port, ID_EX_RF_OUT1_NEXT_31_port, 
      ID_EX_RF_OUT1_NEXT_30_port, ID_EX_RF_OUT1_NEXT_29_port, 
      ID_EX_RF_OUT1_NEXT_28_port, ID_EX_RF_OUT1_NEXT_27_port, 
      ID_EX_RF_OUT1_NEXT_26_port, ID_EX_RF_OUT1_NEXT_25_port, 
      ID_EX_RF_OUT1_NEXT_24_port, ID_EX_RF_OUT1_NEXT_23_port, 
      ID_EX_RF_OUT1_NEXT_22_port, ID_EX_RF_OUT1_NEXT_21_port, 
      ID_EX_RF_OUT1_NEXT_20_port, ID_EX_RF_OUT1_NEXT_19_port, 
      ID_EX_RF_OUT1_NEXT_18_port, ID_EX_RF_OUT1_NEXT_17_port, 
      ID_EX_RF_OUT1_NEXT_16_port, ID_EX_RF_OUT1_NEXT_15_port, 
      ID_EX_RF_OUT1_NEXT_14_port, ID_EX_RF_OUT1_NEXT_13_port, 
      ID_EX_RF_OUT1_NEXT_12_port, ID_EX_RF_OUT1_NEXT_11_port, 
      ID_EX_RF_OUT1_NEXT_10_port, ID_EX_RF_OUT1_NEXT_9_port, 
      ID_EX_RF_OUT1_NEXT_8_port, ID_EX_RF_OUT1_NEXT_7_port, 
      ID_EX_RF_OUT1_NEXT_6_port, ID_EX_RF_OUT1_NEXT_5_port, 
      ID_EX_RF_OUT1_NEXT_4_port, ID_EX_RF_OUT1_NEXT_3_port, 
      ID_EX_RF_OUT1_NEXT_2_port, ID_EX_RF_OUT1_NEXT_1_port, 
      ID_EX_RF_OUT1_NEXT_0_port, ID_EX_RF_OUT2_NEXT_31_port, 
      ID_EX_RF_OUT2_NEXT_30_port, ID_EX_RF_OUT2_NEXT_29_port, 
      ID_EX_RF_OUT2_NEXT_28_port, ID_EX_RF_OUT2_NEXT_27_port, 
      ID_EX_RF_OUT2_NEXT_26_port, ID_EX_RF_OUT2_NEXT_25_port, 
      ID_EX_RF_OUT2_NEXT_24_port, ID_EX_RF_OUT2_NEXT_23_port, 
      ID_EX_RF_OUT2_NEXT_22_port, ID_EX_RF_OUT2_NEXT_21_port, 
      ID_EX_RF_OUT2_NEXT_20_port, ID_EX_RF_OUT2_NEXT_19_port, 
      ID_EX_RF_OUT2_NEXT_18_port, ID_EX_RF_OUT2_NEXT_17_port, 
      ID_EX_RF_OUT2_NEXT_16_port, ID_EX_RF_OUT2_NEXT_15_port, 
      ID_EX_RF_OUT2_NEXT_14_port, ID_EX_RF_OUT2_NEXT_13_port, 
      ID_EX_RF_OUT2_NEXT_12_port, ID_EX_RF_OUT2_NEXT_11_port, 
      ID_EX_RF_OUT2_NEXT_10_port, ID_EX_RF_OUT2_NEXT_9_port, 
      ID_EX_RF_OUT2_NEXT_8_port, ID_EX_RF_OUT2_NEXT_7_port, 
      ID_EX_RF_OUT2_NEXT_6_port, ID_EX_RF_OUT2_NEXT_5_port, 
      ID_EX_RF_OUT2_NEXT_4_port, ID_EX_RF_OUT2_NEXT_3_port, 
      ID_EX_RF_OUT2_NEXT_2_port, ID_EX_RF_OUT2_NEXT_1_port, 
      ID_EX_RF_OUT2_NEXT_0_port, ID_EX_IMM_NEXT_31_port, ID_EX_IMM_NEXT_30_port
      , ID_EX_IMM_NEXT_29_port, ID_EX_IMM_NEXT_28_port, ID_EX_IMM_NEXT_27_port,
      ID_EX_IMM_NEXT_26_port, ID_EX_IMM_NEXT_25_port, ID_EX_IMM_NEXT_24_port, 
      ID_EX_IMM_NEXT_23_port, ID_EX_IMM_NEXT_22_port, ID_EX_IMM_NEXT_21_port, 
      ID_EX_IMM_NEXT_20_port, ID_EX_IMM_NEXT_19_port, ID_EX_IMM_NEXT_18_port, 
      ID_EX_IMM_NEXT_17_port, ID_EX_IMM_NEXT_16_port, ID_EX_IMM_NEXT_15_port, 
      ID_EX_IMM_NEXT_14_port, ID_EX_IMM_NEXT_13_port, ID_EX_IMM_NEXT_12_port, 
      ID_EX_IMM_NEXT_11_port, ID_EX_IMM_NEXT_10_port, ID_EX_IMM_NEXT_9_port, 
      ID_EX_IMM_NEXT_8_port, ID_EX_IMM_NEXT_7_port, ID_EX_IMM_NEXT_6_port, 
      ID_EX_IMM_NEXT_5_port, ID_EX_IMM_NEXT_4_port, ID_EX_IMM_NEXT_3_port, 
      ID_EX_IMM_NEXT_2_port, ID_EX_IMM_NEXT_1_port, ID_EX_IMM_NEXT_0_port, 
      EX_MEM_ALU_OUTPUT_NEXT_31_port, EX_MEM_ALU_OUTPUT_NEXT_30_port, 
      EX_MEM_ALU_OUTPUT_NEXT_29_port, EX_MEM_ALU_OUTPUT_NEXT_28_port, 
      EX_MEM_ALU_OUTPUT_NEXT_27_port, EX_MEM_ALU_OUTPUT_NEXT_26_port, 
      EX_MEM_ALU_OUTPUT_NEXT_25_port, EX_MEM_ALU_OUTPUT_NEXT_24_port, 
      EX_MEM_ALU_OUTPUT_NEXT_23_port, EX_MEM_ALU_OUTPUT_NEXT_22_port, 
      EX_MEM_ALU_OUTPUT_NEXT_21_port, EX_MEM_ALU_OUTPUT_NEXT_20_port, 
      EX_MEM_ALU_OUTPUT_NEXT_19_port, EX_MEM_ALU_OUTPUT_NEXT_18_port, 
      EX_MEM_ALU_OUTPUT_NEXT_17_port, EX_MEM_ALU_OUTPUT_NEXT_16_port, 
      EX_MEM_ALU_OUTPUT_NEXT_15_port, EX_MEM_ALU_OUTPUT_NEXT_14_port, 
      EX_MEM_ALU_OUTPUT_NEXT_13_port, EX_MEM_ALU_OUTPUT_NEXT_12_port, 
      EX_MEM_ALU_OUTPUT_NEXT_11_port, EX_MEM_ALU_OUTPUT_NEXT_10_port, 
      EX_MEM_ALU_OUTPUT_NEXT_9_port, EX_MEM_ALU_OUTPUT_NEXT_8_port, 
      EX_MEM_ALU_OUTPUT_NEXT_7_port, EX_MEM_ALU_OUTPUT_NEXT_6_port, 
      EX_MEM_ALU_OUTPUT_NEXT_5_port, EX_MEM_ALU_OUTPUT_NEXT_4_port, 
      EX_MEM_ALU_OUTPUT_NEXT_3_port, EX_MEM_ALU_OUTPUT_NEXT_2_port, 
      EX_MEM_ALU_OUTPUT_NEXT_1_port, EX_MEM_ALU_OUTPUT_NEXT_0_port, 
      EX_MEM_BRANCH_DETECT_NEXT, MEM_WB_DRAM_OUTPUT_NEXT_31_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_30_port, MEM_WB_DRAM_OUTPUT_NEXT_29_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_28_port, MEM_WB_DRAM_OUTPUT_NEXT_27_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_26_port, MEM_WB_DRAM_OUTPUT_NEXT_25_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_24_port, MEM_WB_DRAM_OUTPUT_NEXT_23_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_22_port, MEM_WB_DRAM_OUTPUT_NEXT_21_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_20_port, MEM_WB_DRAM_OUTPUT_NEXT_19_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_18_port, MEM_WB_DRAM_OUTPUT_NEXT_17_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_16_port, MEM_WB_DRAM_OUTPUT_NEXT_15_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_14_port, MEM_WB_DRAM_OUTPUT_NEXT_13_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_12_port, MEM_WB_DRAM_OUTPUT_NEXT_11_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_10_port, MEM_WB_DRAM_OUTPUT_NEXT_9_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_8_port, MEM_WB_DRAM_OUTPUT_NEXT_7_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_6_port, MEM_WB_DRAM_OUTPUT_NEXT_5_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_4_port, MEM_WB_DRAM_OUTPUT_NEXT_3_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_2_port, MEM_WB_DRAM_OUTPUT_NEXT_1_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_0_port, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11,
      N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26
      , N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, 
      N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55
      , N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, 
      N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84
      , N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, 
      N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, 
      N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, 
      N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, 
      N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, 
      N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, 
      N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, 
      N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, 
      N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, 
      N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, 
      N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, 
      N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, 
      N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, 
      N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, 
      N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, 
      N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, 
      N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, 
      N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, 
      N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, 
      N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, 
      N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, 
      N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, 
      N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, 
      N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, 
      N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, 
      N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, 
      N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, 
      N411, N412, N413, N414, NPC_BUS_31_port, NPC_BUS_30_port, NPC_BUS_29_port
      , NPC_BUS_28_port, NPC_BUS_27_port, NPC_BUS_26_port, NPC_BUS_25_port, 
      NPC_BUS_24_port, NPC_BUS_23_port, NPC_BUS_22_port, NPC_BUS_21_port, 
      NPC_BUS_20_port, NPC_BUS_19_port, NPC_BUS_18_port, NPC_BUS_17_port, 
      NPC_BUS_16_port, NPC_BUS_15_port, NPC_BUS_14_port, NPC_BUS_13_port, 
      NPC_BUS_12_port, NPC_BUS_11_port, NPC_BUS_10_port, NPC_BUS_9_port, 
      NPC_BUS_8_port, NPC_BUS_7_port, NPC_BUS_6_port, NPC_BUS_5_port, 
      NPC_BUS_4_port, NPC_BUS_3_port, NPC_BUS_2_port, NPC_BUS_1_port, 
      NPC_BUS_0_port, ZERO_OUT, PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port,
      PC_BUS_28_port, PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, 
      PC_BUS_24_port, PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, 
      PC_BUS_20_port, PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, 
      PC_BUS_16_port, PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, 
      PC_BUS_12_port, PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, 
      PC_BUS_8_port, PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port
      , PC_BUS_3_port, PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, 
      JAL_MUX_OUT_31_port, JAL_MUX_OUT_30_port, JAL_MUX_OUT_29_port, 
      JAL_MUX_OUT_28_port, JAL_MUX_OUT_27_port, JAL_MUX_OUT_26_port, 
      JAL_MUX_OUT_25_port, JAL_MUX_OUT_24_port, JAL_MUX_OUT_23_port, 
      JAL_MUX_OUT_22_port, JAL_MUX_OUT_21_port, JAL_MUX_OUT_20_port, 
      JAL_MUX_OUT_19_port, JAL_MUX_OUT_18_port, JAL_MUX_OUT_17_port, 
      JAL_MUX_OUT_16_port, JAL_MUX_OUT_15_port, JAL_MUX_OUT_14_port, 
      JAL_MUX_OUT_13_port, JAL_MUX_OUT_12_port, JAL_MUX_OUT_11_port, 
      JAL_MUX_OUT_10_port, JAL_MUX_OUT_9_port, JAL_MUX_OUT_8_port, 
      JAL_MUX_OUT_7_port, JAL_MUX_OUT_6_port, JAL_MUX_OUT_5_port, 
      JAL_MUX_OUT_4_port, JAL_MUX_OUT_3_port, JAL_MUX_OUT_2_port, 
      JAL_MUX_OUT_1_port, JAL_MUX_OUT_0_port, RF_OUT1_31_port, RF_OUT1_30_port,
      RF_OUT1_29_port, RF_OUT1_28_port, RF_OUT1_27_port, RF_OUT1_26_port, 
      RF_OUT1_25_port, RF_OUT1_24_port, RF_OUT1_23_port, RF_OUT1_22_port, 
      RF_OUT1_21_port, RF_OUT1_20_port, RF_OUT1_19_port, RF_OUT1_18_port, 
      RF_OUT1_17_port, RF_OUT1_16_port, RF_OUT1_15_port, RF_OUT1_14_port, 
      RF_OUT1_13_port, RF_OUT1_12_port, RF_OUT1_11_port, RF_OUT1_10_port, 
      RF_OUT1_9_port, RF_OUT1_8_port, RF_OUT1_7_port, RF_OUT1_6_port, 
      RF_OUT1_5_port, RF_OUT1_4_port, RF_OUT1_3_port, RF_OUT1_2_port, 
      RF_OUT1_1_port, RF_OUT1_0_port, RF_OUT2_31_port, RF_OUT2_30_port, 
      RF_OUT2_29_port, RF_OUT2_28_port, RF_OUT2_27_port, RF_OUT2_26_port, 
      RF_OUT2_25_port, RF_OUT2_24_port, RF_OUT2_23_port, RF_OUT2_22_port, 
      RF_OUT2_21_port, RF_OUT2_20_port, RF_OUT2_19_port, RF_OUT2_18_port, 
      RF_OUT2_17_port, RF_OUT2_16_port, RF_OUT2_15_port, RF_OUT2_14_port, 
      RF_OUT2_13_port, RF_OUT2_12_port, RF_OUT2_11_port, RF_OUT2_10_port, 
      RF_OUT2_9_port, RF_OUT2_8_port, RF_OUT2_7_port, RF_OUT2_6_port, 
      RF_OUT2_5_port, RF_OUT2_4_port, RF_OUT2_3_port, RF_OUT2_2_port, 
      RF_OUT2_1_port, RF_OUT2_0_port, IMM_OUT_31_port, IMM_OUT_30_port, 
      IMM_OUT_29_port, IMM_OUT_28_port, IMM_OUT_27_port, IMM_OUT_26_port, 
      IMM_OUT_25_port, IMM_OUT_24_port, IMM_OUT_23_port, IMM_OUT_22_port, 
      IMM_OUT_21_port, IMM_OUT_20_port, IMM_OUT_19_port, IMM_OUT_18_port, 
      IMM_OUT_17_port, IMM_OUT_16_port, IMM_OUT_15_port, IMM_OUT_14_port, 
      IMM_OUT_13_port, IMM_OUT_12_port, IMM_OUT_11_port, IMM_OUT_10_port, 
      IMM_OUT_9_port, IMM_OUT_8_port, IMM_OUT_7_port, IMM_OUT_6_port, 
      IMM_OUT_5_port, IMM_OUT_4_port, IMM_OUT_3_port, IMM_OUT_2_port, 
      IMM_OUT_1_port, IMM_OUT_0_port, FORWARD_A_1_port, FORWARD_A_0_port, 
      ALU_PREOP1_31_port, ALU_PREOP1_30_port, ALU_PREOP1_29_port, 
      ALU_PREOP1_28_port, ALU_PREOP1_27_port, ALU_PREOP1_26_port, 
      ALU_PREOP1_25_port, ALU_PREOP1_24_port, ALU_PREOP1_23_port, 
      ALU_PREOP1_22_port, ALU_PREOP1_21_port, ALU_PREOP1_20_port, 
      ALU_PREOP1_19_port, ALU_PREOP1_18_port, ALU_PREOP1_17_port, 
      ALU_PREOP1_16_port, ALU_PREOP1_15_port, ALU_PREOP1_14_port, 
      ALU_PREOP1_13_port, ALU_PREOP1_12_port, ALU_PREOP1_11_port, 
      ALU_PREOP1_10_port, ALU_PREOP1_9_port, ALU_PREOP1_8_port, 
      ALU_PREOP1_7_port, ALU_PREOP1_6_port, ALU_PREOP1_5_port, 
      ALU_PREOP1_4_port, ALU_PREOP1_3_port, ALU_PREOP1_2_port, 
      ALU_PREOP1_1_port, ALU_PREOP1_0_port, FORWARD_B_1_port, FORWARD_B_0_port,
      ALU_PREOP2_31_port, ALU_PREOP2_30_port, ALU_PREOP2_29_port, 
      ALU_PREOP2_28_port, ALU_PREOP2_27_port, ALU_PREOP2_26_port, 
      ALU_PREOP2_25_port, ALU_PREOP2_24_port, ALU_PREOP2_23_port, 
      ALU_PREOP2_22_port, ALU_PREOP2_21_port, ALU_PREOP2_20_port, 
      ALU_PREOP2_19_port, ALU_PREOP2_18_port, ALU_PREOP2_17_port, 
      ALU_PREOP2_16_port, ALU_PREOP2_15_port, ALU_PREOP2_14_port, 
      ALU_PREOP2_13_port, ALU_PREOP2_12_port, ALU_PREOP2_11_port, 
      ALU_PREOP2_10_port, ALU_PREOP2_9_port, ALU_PREOP2_8_port, 
      ALU_PREOP2_7_port, ALU_PREOP2_6_port, ALU_PREOP2_5_port, 
      ALU_PREOP2_4_port, ALU_PREOP2_3_port, ALU_PREOP2_2_port, 
      ALU_PREOP2_1_port, ALU_PREOP2_0_port, ALU_OP1_31_port, ALU_OP1_30_port, 
      ALU_OP1_29_port, ALU_OP1_28_port, ALU_OP1_27_port, ALU_OP1_26_port, 
      ALU_OP1_25_port, ALU_OP1_24_port, ALU_OP1_23_port, ALU_OP1_22_port, 
      ALU_OP1_21_port, ALU_OP1_20_port, ALU_OP1_19_port, ALU_OP1_18_port, 
      ALU_OP1_17_port, ALU_OP1_16_port, ALU_OP1_15_port, ALU_OP1_14_port, 
      ALU_OP1_13_port, ALU_OP1_12_port, ALU_OP1_11_port, ALU_OP1_10_port, 
      ALU_OP1_9_port, ALU_OP1_8_port, ALU_OP1_7_port, ALU_OP1_6_port, 
      ALU_OP1_5_port, ALU_OP1_4_port, ALU_OP1_3_port, ALU_OP1_2_port, 
      ALU_OP1_1_port, ALU_OP1_0_port, ALU_OP2_31_port, ALU_OP2_30_port, 
      ALU_OP2_29_port, ALU_OP2_28_port, ALU_OP2_27_port, ALU_OP2_26_port, 
      ALU_OP2_25_port, ALU_OP2_24_port, ALU_OP2_23_port, ALU_OP2_22_port, 
      ALU_OP2_21_port, ALU_OP2_20_port, ALU_OP2_19_port, ALU_OP2_18_port, 
      ALU_OP2_17_port, ALU_OP2_16_port, ALU_OP2_15_port, ALU_OP2_14_port, 
      ALU_OP2_13_port, ALU_OP2_12_port, ALU_OP2_11_port, ALU_OP2_10_port, 
      ALU_OP2_9_port, ALU_OP2_8_port, ALU_OP2_7_port, ALU_OP2_6_port, 
      ALU_OP2_5_port, ALU_OP2_4_port, ALU_OP2_3_port, ALU_OP2_2_port, 
      ALU_OP2_1_port, ALU_OP2_0_port, ALU_OUTPUT_31_port, ALU_OUTPUT_30_port, 
      ALU_OUTPUT_29_port, ALU_OUTPUT_28_port, ALU_OUTPUT_27_port, 
      ALU_OUTPUT_26_port, ALU_OUTPUT_25_port, ALU_OUTPUT_24_port, 
      ALU_OUTPUT_23_port, ALU_OUTPUT_22_port, ALU_OUTPUT_21_port, 
      ALU_OUTPUT_20_port, ALU_OUTPUT_19_port, ALU_OUTPUT_18_port, 
      ALU_OUTPUT_17_port, ALU_OUTPUT_16_port, ALU_OUTPUT_15_port, 
      ALU_OUTPUT_14_port, ALU_OUTPUT_13_port, ALU_OUTPUT_12_port, 
      ALU_OUTPUT_11_port, ALU_OUTPUT_10_port, ALU_OUTPUT_9_port, 
      ALU_OUTPUT_8_port, ALU_OUTPUT_7_port, ALU_OUTPUT_6_port, 
      ALU_OUTPUT_5_port, ALU_OUTPUT_4_port, ALU_OUTPUT_3_port, 
      ALU_OUTPUT_2_port, ALU_OUTPUT_1_port, ALU_OUTPUT_0_port, BRANCH_DETECT, 
      WB_MUX_OUT_31_port, WB_MUX_OUT_30_port, WB_MUX_OUT_29_port, 
      WB_MUX_OUT_28_port, WB_MUX_OUT_27_port, WB_MUX_OUT_26_port, 
      WB_MUX_OUT_25_port, WB_MUX_OUT_24_port, WB_MUX_OUT_23_port, 
      WB_MUX_OUT_22_port, WB_MUX_OUT_21_port, WB_MUX_OUT_20_port, 
      WB_MUX_OUT_19_port, WB_MUX_OUT_18_port, WB_MUX_OUT_17_port, 
      WB_MUX_OUT_16_port, WB_MUX_OUT_15_port, WB_MUX_OUT_14_port, 
      WB_MUX_OUT_13_port, WB_MUX_OUT_12_port, WB_MUX_OUT_11_port, 
      WB_MUX_OUT_10_port, WB_MUX_OUT_9_port, WB_MUX_OUT_8_port, 
      WB_MUX_OUT_7_port, WB_MUX_OUT_6_port, WB_MUX_OUT_5_port, 
      WB_MUX_OUT_4_port, WB_MUX_OUT_3_port, WB_MUX_OUT_2_port, 
      WB_MUX_OUT_1_port, WB_MUX_OUT_0_port, n1, n5_port, net31024, net31028, 
      net31098, net31096, net31094, net31092, net31090, net31088, net31086, 
      net31084, net31082, net31080, net31078, net31076, net31074, net31072, 
      net31070, net31068, net31066, net31064, net31062, net31060, net31058, 
      net31056, net31054, net31046, net31044, net31260, net31258, n2_port, 
      n3_port, n4_port, n6_port, n7_port, n8_port, n9_port, n10_port, n11_port,
      n12_port, n13_port, n14_port, n15_port, n16_port, n17_port, n18_port, 
      n19_port, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313,
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, 
      n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, 
      n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, 
      n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, 
      n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, 
      n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, 
      n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, 
      n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, 
      n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, 
      n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, 
      n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, 
      n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, 
      n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, 
      n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, 
      n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, 
      n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, 
      n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, 
      n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, 
      n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, 
      n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, 
      n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, 
      n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, 
      n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, 
      n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, 
      n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, 
      n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, 
      n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, 
      n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, 
      n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, 
      n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, 
      n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, 
      n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, 
      n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, 
      n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, 
      n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, 
      n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, 
      n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, 
      n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, 
      n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, 
      n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, 
      n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, 
      n_1710, n_1711, n_1712, n_1713, n_1714, n_1715 : std_logic;

begin
   IR_OUT <= ( IR_OUT_31_port, IR_OUT_30_port, IR_OUT_29_port, IR_OUT_28_port, 
      IR_OUT_27_port, IR_OUT_26_port, IR_OUT_25_port, IR_OUT_24_port, 
      IR_OUT_23_port, IR_OUT_22_port, IR_OUT_21_port, IR_OUT_20_port, 
      IR_OUT_19_port, IR_OUT_18_port, IR_OUT_17_port, IR_OUT_16_port, 
      IR_OUT_15_port, IR_OUT_14_port, IR_OUT_13_port, IR_OUT_12_port, 
      IR_OUT_11_port, IR_OUT_10_port, IR_OUT_9_port, IR_OUT_8_port, 
      IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port, IR_OUT_4_port, IR_OUT_3_port
      , IR_OUT_2_port, IR_OUT_1_port, IR_OUT_0_port );
   PC_OUT <= ( PC_OUT_31_port, PC_OUT_30_port, PC_OUT_29_port, PC_OUT_28_port, 
      PC_OUT_27_port, PC_OUT_26_port, PC_OUT_25_port, PC_OUT_24_port, 
      PC_OUT_23_port, PC_OUT_22_port, PC_OUT_21_port, PC_OUT_20_port, 
      PC_OUT_19_port, PC_OUT_18_port, PC_OUT_17_port, PC_OUT_16_port, 
      PC_OUT_15_port, PC_OUT_14_port, PC_OUT_13_port, PC_OUT_12_port, 
      PC_OUT_11_port, PC_OUT_10_port, PC_OUT_9_port, PC_OUT_8_port, 
      PC_OUT_7_port, PC_OUT_6_port, PC_OUT_5_port, PC_OUT_4_port, PC_OUT_3_port
      , PC_OUT_2_port, PC_OUT_1_port, PC_OUT_0_port );
   ALU_OUT <= ( ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, 
      ALU_OUT_28_port, ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, 
      ALU_OUT_24_port, ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, 
      ALU_OUT_20_port, ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, 
      ALU_OUT_16_port, ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, 
      ALU_OUT_12_port, ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, 
      ALU_OUT_8_port, ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, 
      ALU_OUT_4_port, ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, 
      ALU_OUT_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n1 <= '0';
   IF_ID_IR_reg_30_inst : DFF_X1 port map( D => N64, CK => CLK, Q => 
                           IF_ID_IR_30_port, QN => n4_port);
   IF_ID_IR_reg_29_inst : DFF_X1 port map( D => N63, CK => CLK, Q => 
                           IF_ID_IR_29_port, QN => n9_port);
   IF_ID_IR_reg_27_inst : DFF_X1 port map( D => N61, CK => CLK, Q => 
                           IF_ID_IR_27_port, QN => n16_port);
   IF_ID_IR_reg_26_inst : DFF_X1 port map( D => N60, CK => CLK, Q => 
                           IF_ID_IR_26_port, QN => n14_port);
   IF_ID_IR_reg_25_inst : DFF_X1 port map( D => N59, CK => CLK, Q => 
                           IF_ID_IR_25_port, QN => n_1306);
   IF_ID_IR_reg_24_inst : DFF_X1 port map( D => N58, CK => CLK, Q => 
                           IF_ID_IR_24_port, QN => n_1307);
   IF_ID_IR_reg_23_inst : DFF_X1 port map( D => N57, CK => CLK, Q => 
                           IF_ID_IR_23_port, QN => n_1308);
   IF_ID_IR_reg_22_inst : DFF_X1 port map( D => N56, CK => CLK, Q => 
                           IF_ID_IR_22_port, QN => n_1309);
   IF_ID_IR_reg_21_inst : DFF_X1 port map( D => N55, CK => CLK, Q => 
                           IF_ID_IR_21_port, QN => n_1310);
   IF_ID_IR_reg_20_inst : DFF_X1 port map( D => N54, CK => CLK, Q => 
                           IF_ID_IR_20_port, QN => n_1311);
   IF_ID_IR_reg_19_inst : DFF_X1 port map( D => N53, CK => CLK, Q => 
                           IF_ID_IR_19_port, QN => n_1312);
   IF_ID_IR_reg_18_inst : DFF_X1 port map( D => N52, CK => CLK, Q => 
                           IF_ID_IR_18_port, QN => n_1313);
   IF_ID_IR_reg_17_inst : DFF_X1 port map( D => N51, CK => CLK, Q => 
                           IF_ID_IR_17_port, QN => n_1314);
   IF_ID_IR_reg_16_inst : DFF_X1 port map( D => N50, CK => CLK, Q => 
                           IF_ID_IR_16_port, QN => n_1315);
   IF_ID_IR_reg_15_inst : DFF_X1 port map( D => N49, CK => CLK, Q => 
                           IF_ID_IR_15_port, QN => n_1316);
   IF_ID_IR_reg_14_inst : DFF_X1 port map( D => N48, CK => CLK, Q => 
                           IF_ID_IR_14_port, QN => n_1317);
   IF_ID_IR_reg_13_inst : DFF_X1 port map( D => N47, CK => CLK, Q => 
                           IF_ID_IR_13_port, QN => n_1318);
   IF_ID_IR_reg_12_inst : DFF_X1 port map( D => N46, CK => CLK, Q => 
                           IF_ID_IR_12_port, QN => n_1319);
   IF_ID_IR_reg_11_inst : DFF_X1 port map( D => N45, CK => CLK, Q => 
                           IF_ID_IR_11_port, QN => n_1320);
   IF_ID_IR_reg_10_inst : DFF_X1 port map( D => N44, CK => CLK, Q => 
                           IF_ID_IR_10_port, QN => n_1321);
   IF_ID_IR_reg_9_inst : DFF_X1 port map( D => N43, CK => CLK, Q => 
                           IF_ID_IR_9_port, QN => n_1322);
   IF_ID_IR_reg_8_inst : DFF_X1 port map( D => N42, CK => CLK, Q => 
                           IF_ID_IR_8_port, QN => n_1323);
   IF_ID_IR_reg_7_inst : DFF_X1 port map( D => N41, CK => CLK, Q => 
                           IF_ID_IR_7_port, QN => n_1324);
   IF_ID_IR_reg_6_inst : DFF_X1 port map( D => N40, CK => CLK, Q => 
                           IF_ID_IR_6_port, QN => n_1325);
   IF_ID_IR_reg_5_inst : DFF_X1 port map( D => N39, CK => CLK, Q => 
                           IF_ID_IR_5_port, QN => n_1326);
   IF_ID_IR_reg_4_inst : DFF_X1 port map( D => N38, CK => CLK, Q => 
                           IF_ID_IR_4_port, QN => n_1327);
   IF_ID_IR_reg_3_inst : DFF_X1 port map( D => N37, CK => CLK, Q => 
                           IF_ID_IR_3_port, QN => n_1328);
   IF_ID_IR_reg_2_inst : DFF_X1 port map( D => N36, CK => CLK, Q => 
                           IF_ID_IR_2_port, QN => n_1329);
   IF_ID_IR_reg_1_inst : DFF_X1 port map( D => N35, CK => CLK, Q => 
                           IF_ID_IR_1_port, QN => n_1330);
   IF_ID_IR_reg_0_inst : DFF_X1 port map( D => N34, CK => CLK, Q => 
                           IF_ID_IR_0_port, QN => n_1331);
   ID_EX_RF_WE_reg : DFF_X1 port map( D => N98, CK => CLK, Q => ID_EX_RF_WE, QN
                           => n_1332);
   ID_EX_RS1_reg_3_inst : DFF_X1 port map( D => N102, CK => CLK, Q => 
                           ID_EX_RS1_3_port, QN => n_1333);
   ID_EX_RS1_reg_2_inst : DFF_X1 port map( D => N101, CK => CLK, Q => 
                           ID_EX_RS1_2_port, QN => n_1334);
   ID_EX_RS1_reg_1_inst : DFF_X1 port map( D => N100, CK => CLK, Q => 
                           ID_EX_RS1_1_port, QN => n_1335);
   ID_EX_RS1_reg_0_inst : DFF_X1 port map( D => N99, CK => CLK, Q => 
                           ID_EX_RS1_0_port, QN => n_1336);
   ID_EX_RD_reg_3_inst : DFF_X1 port map( D => N112, CK => CLK, Q => 
                           ID_EX_RD_3_port, QN => n_1337);
   ID_EX_RD_reg_1_inst : DFF_X1 port map( D => N110, CK => CLK, Q => 
                           ID_EX_RD_1_port, QN => n_1338);
   ID_EX_IMM_reg_31_inst : DFF_X1 port map( D => N209, CK => CLK, Q => 
                           ID_EX_IMM_31_port, QN => n_1339);
   ID_EX_IMM_reg_30_inst : DFF_X1 port map( D => N208, CK => CLK, Q => 
                           ID_EX_IMM_30_port, QN => n_1340);
   ID_EX_IMM_reg_29_inst : DFF_X1 port map( D => N207, CK => CLK, Q => 
                           ID_EX_IMM_29_port, QN => n_1341);
   ID_EX_IMM_reg_28_inst : DFF_X1 port map( D => N206, CK => CLK, Q => 
                           ID_EX_IMM_28_port, QN => n_1342);
   ID_EX_IMM_reg_27_inst : DFF_X1 port map( D => N205, CK => CLK, Q => 
                           ID_EX_IMM_27_port, QN => n_1343);
   ID_EX_IMM_reg_26_inst : DFF_X1 port map( D => N204, CK => CLK, Q => 
                           ID_EX_IMM_26_port, QN => n_1344);
   ID_EX_IMM_reg_25_inst : DFF_X1 port map( D => N203, CK => CLK, Q => 
                           ID_EX_IMM_25_port, QN => n_1345);
   ID_EX_IMM_reg_24_inst : DFF_X1 port map( D => N202, CK => CLK, Q => 
                           ID_EX_IMM_24_port, QN => n_1346);
   ID_EX_IMM_reg_23_inst : DFF_X1 port map( D => N201, CK => CLK, Q => 
                           ID_EX_IMM_23_port, QN => n_1347);
   ID_EX_IMM_reg_22_inst : DFF_X1 port map( D => N200, CK => CLK, Q => 
                           ID_EX_IMM_22_port, QN => n_1348);
   ID_EX_IMM_reg_21_inst : DFF_X1 port map( D => N199, CK => CLK, Q => 
                           ID_EX_IMM_21_port, QN => n_1349);
   ID_EX_IMM_reg_20_inst : DFF_X1 port map( D => N198, CK => CLK, Q => 
                           ID_EX_IMM_20_port, QN => n_1350);
   ID_EX_IMM_reg_19_inst : DFF_X1 port map( D => N197, CK => CLK, Q => 
                           ID_EX_IMM_19_port, QN => n_1351);
   ID_EX_IMM_reg_18_inst : DFF_X1 port map( D => N196, CK => CLK, Q => 
                           ID_EX_IMM_18_port, QN => n_1352);
   ID_EX_IMM_reg_17_inst : DFF_X1 port map( D => N195, CK => CLK, Q => 
                           ID_EX_IMM_17_port, QN => n_1353);
   ID_EX_IMM_reg_16_inst : DFF_X1 port map( D => N194, CK => CLK, Q => 
                           ID_EX_IMM_16_port, QN => n_1354);
   ID_EX_IMM_reg_15_inst : DFF_X1 port map( D => N193, CK => CLK, Q => 
                           ID_EX_IMM_15_port, QN => n_1355);
   ID_EX_IMM_reg_14_inst : DFF_X1 port map( D => N192, CK => CLK, Q => 
                           ID_EX_IMM_14_port, QN => n_1356);
   ID_EX_IMM_reg_13_inst : DFF_X1 port map( D => N191, CK => CLK, Q => 
                           ID_EX_IMM_13_port, QN => n_1357);
   ID_EX_IMM_reg_12_inst : DFF_X1 port map( D => N190, CK => CLK, Q => 
                           ID_EX_IMM_12_port, QN => n_1358);
   ID_EX_IMM_reg_11_inst : DFF_X1 port map( D => N189, CK => CLK, Q => 
                           ID_EX_IMM_11_port, QN => n_1359);
   ID_EX_IMM_reg_10_inst : DFF_X1 port map( D => N188, CK => CLK, Q => 
                           ID_EX_IMM_10_port, QN => n_1360);
   ID_EX_IMM_reg_9_inst : DFF_X1 port map( D => N187, CK => CLK, Q => 
                           ID_EX_IMM_9_port, QN => n_1361);
   ID_EX_IMM_reg_8_inst : DFF_X1 port map( D => N186, CK => CLK, Q => 
                           ID_EX_IMM_8_port, QN => n_1362);
   ID_EX_IMM_reg_7_inst : DFF_X1 port map( D => N185, CK => CLK, Q => 
                           ID_EX_IMM_7_port, QN => n_1363);
   ID_EX_IMM_reg_6_inst : DFF_X1 port map( D => N184, CK => CLK, Q => 
                           ID_EX_IMM_6_port, QN => n_1364);
   ID_EX_IMM_reg_5_inst : DFF_X1 port map( D => N183, CK => CLK, Q => 
                           ID_EX_IMM_5_port, QN => n_1365);
   ID_EX_IMM_reg_4_inst : DFF_X1 port map( D => N182, CK => CLK, Q => 
                           ID_EX_IMM_4_port, QN => n_1366);
   ID_EX_IMM_reg_3_inst : DFF_X1 port map( D => N181, CK => CLK, Q => 
                           ID_EX_IMM_3_port, QN => n_1367);
   ID_EX_IMM_reg_2_inst : DFF_X1 port map( D => N180, CK => CLK, Q => 
                           ID_EX_IMM_2_port, QN => n_1368);
   ID_EX_IMM_reg_1_inst : DFF_X1 port map( D => N179, CK => CLK, Q => 
                           ID_EX_IMM_1_port, QN => n_1369);
   ID_EX_IMM_reg_0_inst : DFF_X1 port map( D => N178, CK => CLK, Q => 
                           ID_EX_IMM_0_port, QN => n_1370);
   EX_MEM_RF_WE_reg : DFF_X1 port map( D => N242, CK => CLK, Q => EX_MEM_RF_WE,
                           QN => n_1371);
   EX_MEM_RD_reg_4_inst : DFF_X1 port map( D => N312, CK => CLK, Q => 
                           EX_MEM_RD_4_port, QN => n_1372);
   EX_MEM_RD_reg_3_inst : DFF_X1 port map( D => N311, CK => CLK, Q => 
                           EX_MEM_RD_3_port, QN => n_1373);
   EX_MEM_RD_reg_2_inst : DFF_X1 port map( D => N310, CK => CLK, Q => 
                           EX_MEM_RD_2_port, QN => n_1374);
   EX_MEM_RD_reg_1_inst : DFF_X1 port map( D => N309, CK => CLK, Q => 
                           EX_MEM_RD_1_port, QN => n_1375);
   EX_MEM_RD_reg_0_inst : DFF_X1 port map( D => N308, CK => CLK, Q => 
                           EX_MEM_RD_0_port, QN => n_1376);
   MEM_WB_RF_WE_reg : DFF_X1 port map( D => N345, CK => CLK, Q => MEM_WB_RF_WE,
                           QN => n_1377);
   MEM_WB_DRAM_OUTPUT_reg_31_inst : DFF_X1 port map( D => N409, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_31_port, QN => n_1378);
   MEM_WB_DRAM_OUTPUT_reg_30_inst : DFF_X1 port map( D => N408, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_30_port, QN => n_1379);
   MEM_WB_DRAM_OUTPUT_reg_29_inst : DFF_X1 port map( D => N407, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_29_port, QN => n_1380);
   MEM_WB_DRAM_OUTPUT_reg_28_inst : DFF_X1 port map( D => N406, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_28_port, QN => n_1381);
   MEM_WB_DRAM_OUTPUT_reg_27_inst : DFF_X1 port map( D => N405, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_27_port, QN => n_1382);
   MEM_WB_DRAM_OUTPUT_reg_26_inst : DFF_X1 port map( D => N404, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_26_port, QN => n_1383);
   MEM_WB_DRAM_OUTPUT_reg_25_inst : DFF_X1 port map( D => N403, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_25_port, QN => n_1384);
   MEM_WB_DRAM_OUTPUT_reg_24_inst : DFF_X1 port map( D => N402, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_24_port, QN => n_1385);
   MEM_WB_DRAM_OUTPUT_reg_23_inst : DFF_X1 port map( D => N401, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_23_port, QN => n_1386);
   MEM_WB_DRAM_OUTPUT_reg_22_inst : DFF_X1 port map( D => N400, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_22_port, QN => n_1387);
   MEM_WB_DRAM_OUTPUT_reg_21_inst : DFF_X1 port map( D => N399, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_21_port, QN => n_1388);
   MEM_WB_DRAM_OUTPUT_reg_20_inst : DFF_X1 port map( D => N398, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_20_port, QN => n_1389);
   MEM_WB_DRAM_OUTPUT_reg_19_inst : DFF_X1 port map( D => N397, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_19_port, QN => n_1390);
   MEM_WB_DRAM_OUTPUT_reg_18_inst : DFF_X1 port map( D => N396, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_18_port, QN => n_1391);
   MEM_WB_DRAM_OUTPUT_reg_17_inst : DFF_X1 port map( D => N395, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_17_port, QN => n_1392);
   MEM_WB_DRAM_OUTPUT_reg_16_inst : DFF_X1 port map( D => N394, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_16_port, QN => n_1393);
   MEM_WB_DRAM_OUTPUT_reg_15_inst : DFF_X1 port map( D => N393, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_15_port, QN => n_1394);
   MEM_WB_DRAM_OUTPUT_reg_14_inst : DFF_X1 port map( D => N392, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_14_port, QN => n_1395);
   MEM_WB_DRAM_OUTPUT_reg_13_inst : DFF_X1 port map( D => N391, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_13_port, QN => n_1396);
   MEM_WB_DRAM_OUTPUT_reg_12_inst : DFF_X1 port map( D => N390, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_12_port, QN => n_1397);
   MEM_WB_DRAM_OUTPUT_reg_11_inst : DFF_X1 port map( D => N389, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_11_port, QN => n_1398);
   MEM_WB_DRAM_OUTPUT_reg_10_inst : DFF_X1 port map( D => N388, CK => CLK, Q =>
                           MEM_WB_DRAM_OUTPUT_10_port, QN => n_1399);
   MEM_WB_DRAM_OUTPUT_reg_9_inst : DFF_X1 port map( D => N387, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_9_port, QN => n_1400);
   MEM_WB_DRAM_OUTPUT_reg_8_inst : DFF_X1 port map( D => N386, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_8_port, QN => n_1401);
   MEM_WB_DRAM_OUTPUT_reg_7_inst : DFF_X1 port map( D => N385, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_7_port, QN => n_1402);
   MEM_WB_DRAM_OUTPUT_reg_6_inst : DFF_X1 port map( D => N384, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_6_port, QN => n_1403);
   MEM_WB_DRAM_OUTPUT_reg_5_inst : DFF_X1 port map( D => N383, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_5_port, QN => n_1404);
   MEM_WB_DRAM_OUTPUT_reg_4_inst : DFF_X1 port map( D => N382, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_4_port, QN => n_1405);
   MEM_WB_DRAM_OUTPUT_reg_3_inst : DFF_X1 port map( D => N381, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_3_port, QN => n_1406);
   MEM_WB_DRAM_OUTPUT_reg_2_inst : DFF_X1 port map( D => N380, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_2_port, QN => n_1407);
   MEM_WB_DRAM_OUTPUT_reg_1_inst : DFF_X1 port map( D => N379, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_1_port, QN => n_1408);
   MEM_WB_DRAM_OUTPUT_reg_0_inst : DFF_X1 port map( D => N378, CK => CLK, Q => 
                           MEM_WB_DRAM_OUTPUT_0_port, QN => n_1409);
   MEM_WB_RD_reg_4_inst : DFF_X1 port map( D => N414, CK => CLK, Q => 
                           MEM_WB_RD_4_port, QN => n_1410);
   MEM_WB_RD_reg_3_inst : DFF_X1 port map( D => N413, CK => CLK, Q => 
                           MEM_WB_RD_3_port, QN => n_1411);
   MEM_WB_RD_reg_2_inst : DFF_X1 port map( D => N412, CK => CLK, Q => 
                           MEM_WB_RD_2_port, QN => n_1412);
   MEM_WB_RD_reg_1_inst : DFF_X1 port map( D => N411, CK => CLK, Q => 
                           MEM_WB_RD_1_port, QN => n_1413);
   MEM_WB_RD_reg_0_inst : DFF_X1 port map( D => N410, CK => CLK, Q => 
                           MEM_WB_RD_0_port, QN => n_1414);
   ID_EX_RF_OUT2_reg_0_inst : DFF_X1 port map( D => N146, CK => CLK, Q => 
                           ID_EX_RF_OUT2_0_port, QN => n_1415);
   EX_MEM_RF_OUT2_reg_0_inst : DFF_X1 port map( D => N243, CK => CLK, Q => 
                           DRAM_IN(0), QN => n_1416);
   ID_EX_RF_OUT2_reg_1_inst : DFF_X1 port map( D => N147, CK => CLK, Q => 
                           ID_EX_RF_OUT2_1_port, QN => n_1417);
   EX_MEM_RF_OUT2_reg_1_inst : DFF_X1 port map( D => N244, CK => CLK, Q => 
                           DRAM_IN(1), QN => n_1418);
   ID_EX_RF_OUT2_reg_2_inst : DFF_X1 port map( D => N148, CK => CLK, Q => 
                           ID_EX_RF_OUT2_2_port, QN => n_1419);
   EX_MEM_RF_OUT2_reg_2_inst : DFF_X1 port map( D => N245, CK => CLK, Q => 
                           DRAM_IN(2), QN => n_1420);
   ID_EX_RF_OUT2_reg_3_inst : DFF_X1 port map( D => N149, CK => CLK, Q => 
                           ID_EX_RF_OUT2_3_port, QN => n_1421);
   EX_MEM_RF_OUT2_reg_3_inst : DFF_X1 port map( D => N246, CK => CLK, Q => 
                           DRAM_IN(3), QN => n_1422);
   ID_EX_RF_OUT2_reg_4_inst : DFF_X1 port map( D => N150, CK => CLK, Q => 
                           ID_EX_RF_OUT2_4_port, QN => n_1423);
   EX_MEM_RF_OUT2_reg_4_inst : DFF_X1 port map( D => N247, CK => CLK, Q => 
                           DRAM_IN(4), QN => n_1424);
   ID_EX_RF_OUT2_reg_5_inst : DFF_X1 port map( D => N151, CK => CLK, Q => 
                           ID_EX_RF_OUT2_5_port, QN => n_1425);
   EX_MEM_RF_OUT2_reg_5_inst : DFF_X1 port map( D => N248, CK => CLK, Q => 
                           DRAM_IN(5), QN => n_1426);
   ID_EX_RF_OUT2_reg_6_inst : DFF_X1 port map( D => N152, CK => CLK, Q => 
                           ID_EX_RF_OUT2_6_port, QN => n_1427);
   EX_MEM_RF_OUT2_reg_6_inst : DFF_X1 port map( D => N249, CK => CLK, Q => 
                           DRAM_IN(6), QN => n_1428);
   ID_EX_RF_OUT2_reg_7_inst : DFF_X1 port map( D => N153, CK => CLK, Q => 
                           ID_EX_RF_OUT2_7_port, QN => n_1429);
   EX_MEM_RF_OUT2_reg_7_inst : DFF_X1 port map( D => N250, CK => CLK, Q => 
                           DRAM_IN(7), QN => n_1430);
   ID_EX_RF_OUT2_reg_8_inst : DFF_X1 port map( D => N154, CK => CLK, Q => 
                           ID_EX_RF_OUT2_8_port, QN => n_1431);
   EX_MEM_RF_OUT2_reg_8_inst : DFF_X1 port map( D => N251, CK => CLK, Q => 
                           DRAM_IN(8), QN => n_1432);
   ID_EX_RF_OUT2_reg_9_inst : DFF_X1 port map( D => N155, CK => CLK, Q => 
                           ID_EX_RF_OUT2_9_port, QN => n_1433);
   EX_MEM_RF_OUT2_reg_9_inst : DFF_X1 port map( D => N252, CK => CLK, Q => 
                           DRAM_IN(9), QN => n_1434);
   ID_EX_RF_OUT2_reg_10_inst : DFF_X1 port map( D => N156, CK => CLK, Q => 
                           ID_EX_RF_OUT2_10_port, QN => n_1435);
   EX_MEM_RF_OUT2_reg_10_inst : DFF_X1 port map( D => N253, CK => CLK, Q => 
                           DRAM_IN(10), QN => n_1436);
   ID_EX_RF_OUT2_reg_11_inst : DFF_X1 port map( D => N157, CK => CLK, Q => 
                           ID_EX_RF_OUT2_11_port, QN => n_1437);
   EX_MEM_RF_OUT2_reg_11_inst : DFF_X1 port map( D => N254, CK => CLK, Q => 
                           DRAM_IN(11), QN => n_1438);
   ID_EX_RF_OUT2_reg_12_inst : DFF_X1 port map( D => N158, CK => CLK, Q => 
                           ID_EX_RF_OUT2_12_port, QN => n_1439);
   EX_MEM_RF_OUT2_reg_12_inst : DFF_X1 port map( D => N255, CK => CLK, Q => 
                           DRAM_IN(12), QN => n_1440);
   ID_EX_RF_OUT2_reg_13_inst : DFF_X1 port map( D => N159, CK => CLK, Q => 
                           ID_EX_RF_OUT2_13_port, QN => n_1441);
   EX_MEM_RF_OUT2_reg_13_inst : DFF_X1 port map( D => N256, CK => CLK, Q => 
                           DRAM_IN(13), QN => n_1442);
   ID_EX_RF_OUT2_reg_14_inst : DFF_X1 port map( D => N160, CK => CLK, Q => 
                           ID_EX_RF_OUT2_14_port, QN => n_1443);
   EX_MEM_RF_OUT2_reg_14_inst : DFF_X1 port map( D => N257, CK => CLK, Q => 
                           DRAM_IN(14), QN => n_1444);
   ID_EX_RF_OUT2_reg_15_inst : DFF_X1 port map( D => N161, CK => CLK, Q => 
                           ID_EX_RF_OUT2_15_port, QN => n_1445);
   EX_MEM_RF_OUT2_reg_15_inst : DFF_X1 port map( D => N258, CK => CLK, Q => 
                           DRAM_IN(15), QN => n_1446);
   ID_EX_RF_OUT2_reg_16_inst : DFF_X1 port map( D => N162, CK => CLK, Q => 
                           ID_EX_RF_OUT2_16_port, QN => n_1447);
   EX_MEM_RF_OUT2_reg_16_inst : DFF_X1 port map( D => N259, CK => CLK, Q => 
                           DRAM_IN(16), QN => n_1448);
   ID_EX_RF_OUT2_reg_17_inst : DFF_X1 port map( D => N163, CK => CLK, Q => 
                           ID_EX_RF_OUT2_17_port, QN => n_1449);
   EX_MEM_RF_OUT2_reg_17_inst : DFF_X1 port map( D => N260, CK => CLK, Q => 
                           DRAM_IN(17), QN => n_1450);
   ID_EX_RF_OUT2_reg_18_inst : DFF_X1 port map( D => N164, CK => CLK, Q => 
                           ID_EX_RF_OUT2_18_port, QN => n_1451);
   EX_MEM_RF_OUT2_reg_18_inst : DFF_X1 port map( D => N261, CK => CLK, Q => 
                           DRAM_IN(18), QN => n_1452);
   ID_EX_RF_OUT2_reg_19_inst : DFF_X1 port map( D => N165, CK => CLK, Q => 
                           ID_EX_RF_OUT2_19_port, QN => n_1453);
   EX_MEM_RF_OUT2_reg_19_inst : DFF_X1 port map( D => N262, CK => CLK, Q => 
                           DRAM_IN(19), QN => n_1454);
   ID_EX_RF_OUT2_reg_20_inst : DFF_X1 port map( D => N166, CK => CLK, Q => 
                           ID_EX_RF_OUT2_20_port, QN => n_1455);
   EX_MEM_RF_OUT2_reg_20_inst : DFF_X1 port map( D => N263, CK => CLK, Q => 
                           DRAM_IN(20), QN => n_1456);
   ID_EX_RF_OUT2_reg_21_inst : DFF_X1 port map( D => N167, CK => CLK, Q => 
                           ID_EX_RF_OUT2_21_port, QN => n_1457);
   EX_MEM_RF_OUT2_reg_21_inst : DFF_X1 port map( D => N264, CK => CLK, Q => 
                           DRAM_IN(21), QN => n_1458);
   ID_EX_RF_OUT2_reg_22_inst : DFF_X1 port map( D => N168, CK => CLK, Q => 
                           ID_EX_RF_OUT2_22_port, QN => n_1459);
   EX_MEM_RF_OUT2_reg_22_inst : DFF_X1 port map( D => N265, CK => CLK, Q => 
                           DRAM_IN(22), QN => n_1460);
   ID_EX_RF_OUT2_reg_23_inst : DFF_X1 port map( D => N169, CK => CLK, Q => 
                           ID_EX_RF_OUT2_23_port, QN => n_1461);
   EX_MEM_RF_OUT2_reg_23_inst : DFF_X1 port map( D => N266, CK => CLK, Q => 
                           DRAM_IN(23), QN => n_1462);
   ID_EX_RF_OUT2_reg_24_inst : DFF_X1 port map( D => N170, CK => CLK, Q => 
                           ID_EX_RF_OUT2_24_port, QN => n_1463);
   EX_MEM_RF_OUT2_reg_24_inst : DFF_X1 port map( D => N267, CK => CLK, Q => 
                           DRAM_IN(24), QN => n_1464);
   ID_EX_RF_OUT2_reg_25_inst : DFF_X1 port map( D => N171, CK => CLK, Q => 
                           ID_EX_RF_OUT2_25_port, QN => n_1465);
   EX_MEM_RF_OUT2_reg_25_inst : DFF_X1 port map( D => N268, CK => CLK, Q => 
                           DRAM_IN(25), QN => n_1466);
   ID_EX_RF_OUT2_reg_26_inst : DFF_X1 port map( D => N172, CK => CLK, Q => 
                           ID_EX_RF_OUT2_26_port, QN => n_1467);
   EX_MEM_RF_OUT2_reg_26_inst : DFF_X1 port map( D => N269, CK => CLK, Q => 
                           DRAM_IN(26), QN => n_1468);
   ID_EX_RF_OUT2_reg_27_inst : DFF_X1 port map( D => N173, CK => CLK, Q => 
                           ID_EX_RF_OUT2_27_port, QN => n_1469);
   EX_MEM_RF_OUT2_reg_27_inst : DFF_X1 port map( D => N270, CK => CLK, Q => 
                           DRAM_IN(27), QN => n_1470);
   ID_EX_RF_OUT2_reg_28_inst : DFF_X1 port map( D => N174, CK => CLK, Q => 
                           ID_EX_RF_OUT2_28_port, QN => n_1471);
   EX_MEM_RF_OUT2_reg_28_inst : DFF_X1 port map( D => N271, CK => CLK, Q => 
                           DRAM_IN(28), QN => n_1472);
   ID_EX_RF_OUT2_reg_29_inst : DFF_X1 port map( D => N175, CK => CLK, Q => 
                           ID_EX_RF_OUT2_29_port, QN => n_1473);
   EX_MEM_RF_OUT2_reg_29_inst : DFF_X1 port map( D => N272, CK => CLK, Q => 
                           DRAM_IN(29), QN => n_1474);
   ID_EX_RF_OUT2_reg_30_inst : DFF_X1 port map( D => N176, CK => CLK, Q => 
                           ID_EX_RF_OUT2_30_port, QN => n_1475);
   EX_MEM_RF_OUT2_reg_30_inst : DFF_X1 port map( D => N273, CK => CLK, Q => 
                           DRAM_IN(30), QN => n_1476);
   ID_EX_RF_OUT2_reg_31_inst : DFF_X1 port map( D => N177, CK => CLK, Q => 
                           ID_EX_RF_OUT2_31_port, QN => n_1477);
   EX_MEM_RF_OUT2_reg_31_inst : DFF_X1 port map( D => N274, CK => CLK, Q => 
                           DRAM_IN(31), QN => n_1478);
   ID_EX_RF_OUT1_reg_0_inst : DFF_X1 port map( D => N114, CK => CLK, Q => 
                           ID_EX_RF_OUT1_0_port, QN => n_1479);
   ID_EX_RF_OUT1_reg_1_inst : DFF_X1 port map( D => N115, CK => CLK, Q => 
                           ID_EX_RF_OUT1_1_port, QN => n_1480);
   ID_EX_RF_OUT1_reg_2_inst : DFF_X1 port map( D => N116, CK => CLK, Q => 
                           ID_EX_RF_OUT1_2_port, QN => n_1481);
   ID_EX_RF_OUT1_reg_3_inst : DFF_X1 port map( D => N117, CK => CLK, Q => 
                           ID_EX_RF_OUT1_3_port, QN => n_1482);
   ID_EX_RF_OUT1_reg_4_inst : DFF_X1 port map( D => N118, CK => CLK, Q => 
                           ID_EX_RF_OUT1_4_port, QN => n_1483);
   ID_EX_RF_OUT1_reg_5_inst : DFF_X1 port map( D => N119, CK => CLK, Q => 
                           ID_EX_RF_OUT1_5_port, QN => n_1484);
   ID_EX_RF_OUT1_reg_6_inst : DFF_X1 port map( D => N120, CK => CLK, Q => 
                           ID_EX_RF_OUT1_6_port, QN => n_1485);
   ID_EX_RF_OUT1_reg_7_inst : DFF_X1 port map( D => N121, CK => CLK, Q => 
                           ID_EX_RF_OUT1_7_port, QN => n_1486);
   ID_EX_RF_OUT1_reg_8_inst : DFF_X1 port map( D => N122, CK => CLK, Q => 
                           ID_EX_RF_OUT1_8_port, QN => n_1487);
   ID_EX_RF_OUT1_reg_9_inst : DFF_X1 port map( D => N123, CK => CLK, Q => 
                           ID_EX_RF_OUT1_9_port, QN => n_1488);
   ID_EX_RF_OUT1_reg_10_inst : DFF_X1 port map( D => N124, CK => CLK, Q => 
                           ID_EX_RF_OUT1_10_port, QN => n_1489);
   ID_EX_RF_OUT1_reg_11_inst : DFF_X1 port map( D => N125, CK => CLK, Q => 
                           ID_EX_RF_OUT1_11_port, QN => n_1490);
   ID_EX_RF_OUT1_reg_12_inst : DFF_X1 port map( D => N126, CK => CLK, Q => 
                           ID_EX_RF_OUT1_12_port, QN => n_1491);
   ID_EX_RF_OUT1_reg_13_inst : DFF_X1 port map( D => N127, CK => CLK, Q => 
                           ID_EX_RF_OUT1_13_port, QN => n_1492);
   ID_EX_RF_OUT1_reg_14_inst : DFF_X1 port map( D => N128, CK => CLK, Q => 
                           ID_EX_RF_OUT1_14_port, QN => n_1493);
   ID_EX_RF_OUT1_reg_15_inst : DFF_X1 port map( D => N129, CK => CLK, Q => 
                           ID_EX_RF_OUT1_15_port, QN => n_1494);
   ID_EX_RF_OUT1_reg_16_inst : DFF_X1 port map( D => N130, CK => CLK, Q => 
                           ID_EX_RF_OUT1_16_port, QN => n_1495);
   ID_EX_RF_OUT1_reg_17_inst : DFF_X1 port map( D => N131, CK => CLK, Q => 
                           ID_EX_RF_OUT1_17_port, QN => n_1496);
   ID_EX_RF_OUT1_reg_18_inst : DFF_X1 port map( D => N132, CK => CLK, Q => 
                           ID_EX_RF_OUT1_18_port, QN => n_1497);
   ID_EX_RF_OUT1_reg_19_inst : DFF_X1 port map( D => N133, CK => CLK, Q => 
                           ID_EX_RF_OUT1_19_port, QN => n_1498);
   ID_EX_RF_OUT1_reg_20_inst : DFF_X1 port map( D => N134, CK => CLK, Q => 
                           ID_EX_RF_OUT1_20_port, QN => n_1499);
   ID_EX_RF_OUT1_reg_21_inst : DFF_X1 port map( D => N135, CK => CLK, Q => 
                           ID_EX_RF_OUT1_21_port, QN => n_1500);
   ID_EX_RF_OUT1_reg_22_inst : DFF_X1 port map( D => N136, CK => CLK, Q => 
                           ID_EX_RF_OUT1_22_port, QN => n_1501);
   ID_EX_RF_OUT1_reg_23_inst : DFF_X1 port map( D => N137, CK => CLK, Q => 
                           ID_EX_RF_OUT1_23_port, QN => n_1502);
   ID_EX_RF_OUT1_reg_24_inst : DFF_X1 port map( D => N138, CK => CLK, Q => 
                           ID_EX_RF_OUT1_24_port, QN => n_1503);
   ID_EX_RF_OUT1_reg_25_inst : DFF_X1 port map( D => N139, CK => CLK, Q => 
                           ID_EX_RF_OUT1_25_port, QN => n_1504);
   ID_EX_RF_OUT1_reg_26_inst : DFF_X1 port map( D => N140, CK => CLK, Q => 
                           ID_EX_RF_OUT1_26_port, QN => n_1505);
   ID_EX_RF_OUT1_reg_27_inst : DFF_X1 port map( D => N141, CK => CLK, Q => 
                           ID_EX_RF_OUT1_27_port, QN => n_1506);
   ID_EX_RF_OUT1_reg_28_inst : DFF_X1 port map( D => N142, CK => CLK, Q => 
                           ID_EX_RF_OUT1_28_port, QN => n_1507);
   ID_EX_RF_OUT1_reg_29_inst : DFF_X1 port map( D => N143, CK => CLK, Q => 
                           ID_EX_RF_OUT1_29_port, QN => n_1508);
   ID_EX_RF_OUT1_reg_30_inst : DFF_X1 port map( D => N144, CK => CLK, Q => 
                           ID_EX_RF_OUT1_30_port, QN => n_1509);
   ID_EX_RF_OUT1_reg_31_inst : DFF_X1 port map( D => N145, CK => CLK, Q => 
                           ID_EX_RF_OUT1_31_port, QN => n_1510);
   EX_MEM_BRANCH_DETECT_reg : DFF_X1 port map( D => N307, CK => CLK, Q => 
                           EX_MEM_BRANCH_DETECT, QN => n_1511);
   EX_MEM_ALU_OUTPUT_reg_0_inst : DFF_X1 port map( D => N275, CK => CLK, Q => 
                           ALU_OUT_0_port, QN => n_1512);
   MEM_WB_ALU_OUTPUT_reg_0_inst : DFF_X1 port map( D => N346, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_0_port, QN => n_1513);
   EX_MEM_ALU_OUTPUT_reg_1_inst : DFF_X1 port map( D => N276, CK => CLK, Q => 
                           ALU_OUT_1_port, QN => n_1514);
   MEM_WB_ALU_OUTPUT_reg_1_inst : DFF_X1 port map( D => N347, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_1_port, QN => n_1515);
   EX_MEM_ALU_OUTPUT_reg_2_inst : DFF_X1 port map( D => N277, CK => CLK, Q => 
                           ALU_OUT_2_port, QN => n_1516);
   MEM_WB_ALU_OUTPUT_reg_2_inst : DFF_X1 port map( D => N348, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_2_port, QN => n_1517);
   EX_MEM_ALU_OUTPUT_reg_3_inst : DFF_X1 port map( D => N278, CK => CLK, Q => 
                           ALU_OUT_3_port, QN => n_1518);
   MEM_WB_ALU_OUTPUT_reg_3_inst : DFF_X1 port map( D => N349, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_3_port, QN => n_1519);
   EX_MEM_ALU_OUTPUT_reg_4_inst : DFF_X1 port map( D => N279, CK => CLK, Q => 
                           ALU_OUT_4_port, QN => n_1520);
   MEM_WB_ALU_OUTPUT_reg_4_inst : DFF_X1 port map( D => N350, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_4_port, QN => n_1521);
   EX_MEM_ALU_OUTPUT_reg_5_inst : DFF_X1 port map( D => N280, CK => CLK, Q => 
                           ALU_OUT_5_port, QN => n_1522);
   MEM_WB_ALU_OUTPUT_reg_5_inst : DFF_X1 port map( D => N351, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_5_port, QN => n_1523);
   EX_MEM_ALU_OUTPUT_reg_6_inst : DFF_X1 port map( D => N281, CK => CLK, Q => 
                           ALU_OUT_6_port, QN => n_1524);
   MEM_WB_ALU_OUTPUT_reg_6_inst : DFF_X1 port map( D => N352, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_6_port, QN => n_1525);
   EX_MEM_ALU_OUTPUT_reg_7_inst : DFF_X1 port map( D => N282, CK => CLK, Q => 
                           ALU_OUT_7_port, QN => n_1526);
   MEM_WB_ALU_OUTPUT_reg_7_inst : DFF_X1 port map( D => N353, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_7_port, QN => n_1527);
   EX_MEM_ALU_OUTPUT_reg_8_inst : DFF_X1 port map( D => N283, CK => CLK, Q => 
                           ALU_OUT_8_port, QN => n_1528);
   MEM_WB_ALU_OUTPUT_reg_8_inst : DFF_X1 port map( D => N354, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_8_port, QN => n_1529);
   EX_MEM_ALU_OUTPUT_reg_9_inst : DFF_X1 port map( D => N284, CK => CLK, Q => 
                           ALU_OUT_9_port, QN => n_1530);
   MEM_WB_ALU_OUTPUT_reg_9_inst : DFF_X1 port map( D => N355, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_9_port, QN => n_1531);
   EX_MEM_ALU_OUTPUT_reg_10_inst : DFF_X1 port map( D => N285, CK => CLK, Q => 
                           ALU_OUT_10_port, QN => n_1532);
   MEM_WB_ALU_OUTPUT_reg_10_inst : DFF_X1 port map( D => N356, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_10_port, QN => n_1533);
   EX_MEM_ALU_OUTPUT_reg_11_inst : DFF_X1 port map( D => N286, CK => CLK, Q => 
                           ALU_OUT_11_port, QN => n_1534);
   MEM_WB_ALU_OUTPUT_reg_11_inst : DFF_X1 port map( D => N357, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_11_port, QN => n_1535);
   EX_MEM_ALU_OUTPUT_reg_12_inst : DFF_X1 port map( D => N287, CK => CLK, Q => 
                           ALU_OUT_12_port, QN => n_1536);
   MEM_WB_ALU_OUTPUT_reg_12_inst : DFF_X1 port map( D => N358, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_12_port, QN => n_1537);
   EX_MEM_ALU_OUTPUT_reg_13_inst : DFF_X1 port map( D => N288, CK => CLK, Q => 
                           ALU_OUT_13_port, QN => n_1538);
   MEM_WB_ALU_OUTPUT_reg_13_inst : DFF_X1 port map( D => N359, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_13_port, QN => n_1539);
   EX_MEM_ALU_OUTPUT_reg_14_inst : DFF_X1 port map( D => N289, CK => CLK, Q => 
                           ALU_OUT_14_port, QN => n_1540);
   MEM_WB_ALU_OUTPUT_reg_14_inst : DFF_X1 port map( D => N360, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_14_port, QN => n_1541);
   EX_MEM_ALU_OUTPUT_reg_15_inst : DFF_X1 port map( D => N290, CK => CLK, Q => 
                           ALU_OUT_15_port, QN => n_1542);
   MEM_WB_ALU_OUTPUT_reg_15_inst : DFF_X1 port map( D => N361, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_15_port, QN => n_1543);
   EX_MEM_ALU_OUTPUT_reg_16_inst : DFF_X1 port map( D => N291, CK => CLK, Q => 
                           ALU_OUT_16_port, QN => n_1544);
   MEM_WB_ALU_OUTPUT_reg_16_inst : DFF_X1 port map( D => N362, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_16_port, QN => n_1545);
   EX_MEM_ALU_OUTPUT_reg_17_inst : DFF_X1 port map( D => N292, CK => CLK, Q => 
                           ALU_OUT_17_port, QN => n_1546);
   MEM_WB_ALU_OUTPUT_reg_17_inst : DFF_X1 port map( D => N363, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_17_port, QN => n_1547);
   EX_MEM_ALU_OUTPUT_reg_18_inst : DFF_X1 port map( D => N293, CK => CLK, Q => 
                           ALU_OUT_18_port, QN => n_1548);
   MEM_WB_ALU_OUTPUT_reg_18_inst : DFF_X1 port map( D => N364, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_18_port, QN => n_1549);
   EX_MEM_ALU_OUTPUT_reg_19_inst : DFF_X1 port map( D => N294, CK => CLK, Q => 
                           ALU_OUT_19_port, QN => n_1550);
   MEM_WB_ALU_OUTPUT_reg_19_inst : DFF_X1 port map( D => N365, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_19_port, QN => n_1551);
   EX_MEM_ALU_OUTPUT_reg_20_inst : DFF_X1 port map( D => N295, CK => CLK, Q => 
                           ALU_OUT_20_port, QN => n_1552);
   MEM_WB_ALU_OUTPUT_reg_20_inst : DFF_X1 port map( D => N366, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_20_port, QN => n_1553);
   EX_MEM_ALU_OUTPUT_reg_21_inst : DFF_X1 port map( D => N296, CK => CLK, Q => 
                           ALU_OUT_21_port, QN => n_1554);
   MEM_WB_ALU_OUTPUT_reg_21_inst : DFF_X1 port map( D => N367, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_21_port, QN => n_1555);
   EX_MEM_ALU_OUTPUT_reg_22_inst : DFF_X1 port map( D => N297, CK => CLK, Q => 
                           ALU_OUT_22_port, QN => n_1556);
   MEM_WB_ALU_OUTPUT_reg_22_inst : DFF_X1 port map( D => N368, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_22_port, QN => n_1557);
   EX_MEM_ALU_OUTPUT_reg_23_inst : DFF_X1 port map( D => N298, CK => CLK, Q => 
                           ALU_OUT_23_port, QN => n_1558);
   MEM_WB_ALU_OUTPUT_reg_23_inst : DFF_X1 port map( D => N369, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_23_port, QN => n_1559);
   EX_MEM_ALU_OUTPUT_reg_24_inst : DFF_X1 port map( D => N299, CK => CLK, Q => 
                           ALU_OUT_24_port, QN => n_1560);
   MEM_WB_ALU_OUTPUT_reg_24_inst : DFF_X1 port map( D => N370, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_24_port, QN => n_1561);
   EX_MEM_ALU_OUTPUT_reg_25_inst : DFF_X1 port map( D => N300, CK => CLK, Q => 
                           ALU_OUT_25_port, QN => n_1562);
   MEM_WB_ALU_OUTPUT_reg_25_inst : DFF_X1 port map( D => N371, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_25_port, QN => n_1563);
   EX_MEM_ALU_OUTPUT_reg_26_inst : DFF_X1 port map( D => N301, CK => CLK, Q => 
                           ALU_OUT_26_port, QN => n_1564);
   MEM_WB_ALU_OUTPUT_reg_26_inst : DFF_X1 port map( D => N372, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_26_port, QN => n_1565);
   EX_MEM_ALU_OUTPUT_reg_27_inst : DFF_X1 port map( D => N302, CK => CLK, Q => 
                           ALU_OUT_27_port, QN => n_1566);
   MEM_WB_ALU_OUTPUT_reg_27_inst : DFF_X1 port map( D => N373, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_27_port, QN => n_1567);
   EX_MEM_ALU_OUTPUT_reg_28_inst : DFF_X1 port map( D => N303, CK => CLK, Q => 
                           ALU_OUT_28_port, QN => n_1568);
   MEM_WB_ALU_OUTPUT_reg_28_inst : DFF_X1 port map( D => N374, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_28_port, QN => n_1569);
   EX_MEM_ALU_OUTPUT_reg_29_inst : DFF_X1 port map( D => N304, CK => CLK, Q => 
                           ALU_OUT_29_port, QN => n_1570);
   MEM_WB_ALU_OUTPUT_reg_29_inst : DFF_X1 port map( D => N375, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_29_port, QN => n_1571);
   EX_MEM_ALU_OUTPUT_reg_30_inst : DFF_X1 port map( D => N305, CK => CLK, Q => 
                           ALU_OUT_30_port, QN => n_1572);
   MEM_WB_ALU_OUTPUT_reg_30_inst : DFF_X1 port map( D => N376, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_30_port, QN => n_1573);
   EX_MEM_ALU_OUTPUT_reg_31_inst : DFF_X1 port map( D => N306, CK => CLK, Q => 
                           ALU_OUT_31_port, QN => n_1574);
   IF_ID_NPC_reg_0_inst : DFF_X1 port map( D => N2, CK => CLK, Q => 
                           IF_ID_NPC_0_port, QN => n_1575);
   ID_EX_NPC_reg_0_inst : DFF_X1 port map( D => N66, CK => CLK, Q => 
                           ID_EX_NPC_0_port, QN => n_1576);
   EX_MEM_NPC_reg_0_inst : DFF_X1 port map( D => N210, CK => CLK, Q => 
                           EX_MEM_NPC_0_port, QN => n_1577);
   MEM_WB_NPC_reg_0_inst : DFF_X1 port map( D => N313, CK => CLK, Q => 
                           MEM_WB_NPC_0_port, QN => n_1578);
   IF_ID_NPC_reg_1_inst : DFF_X1 port map( D => N3, CK => CLK, Q => 
                           IF_ID_NPC_1_port, QN => n_1579);
   ID_EX_NPC_reg_1_inst : DFF_X1 port map( D => N67, CK => CLK, Q => 
                           ID_EX_NPC_1_port, QN => n_1580);
   EX_MEM_NPC_reg_1_inst : DFF_X1 port map( D => N211, CK => CLK, Q => 
                           EX_MEM_NPC_1_port, QN => n_1581);
   MEM_WB_NPC_reg_1_inst : DFF_X1 port map( D => N314, CK => CLK, Q => 
                           MEM_WB_NPC_1_port, QN => n_1582);
   IF_ID_NPC_reg_2_inst : DFF_X1 port map( D => N4, CK => CLK, Q => 
                           IF_ID_NPC_2_port, QN => n_1583);
   ID_EX_NPC_reg_2_inst : DFF_X1 port map( D => N68, CK => CLK, Q => 
                           ID_EX_NPC_2_port, QN => n_1584);
   EX_MEM_NPC_reg_2_inst : DFF_X1 port map( D => N212, CK => CLK, Q => 
                           EX_MEM_NPC_2_port, QN => n_1585);
   MEM_WB_NPC_reg_2_inst : DFF_X1 port map( D => N315, CK => CLK, Q => 
                           MEM_WB_NPC_2_port, QN => n_1586);
   IF_ID_NPC_reg_3_inst : DFF_X1 port map( D => N5, CK => CLK, Q => 
                           IF_ID_NPC_3_port, QN => n_1587);
   ID_EX_NPC_reg_3_inst : DFF_X1 port map( D => N69, CK => CLK, Q => 
                           ID_EX_NPC_3_port, QN => n_1588);
   EX_MEM_NPC_reg_3_inst : DFF_X1 port map( D => N213, CK => CLK, Q => 
                           EX_MEM_NPC_3_port, QN => n_1589);
   MEM_WB_NPC_reg_3_inst : DFF_X1 port map( D => N316, CK => CLK, Q => 
                           MEM_WB_NPC_3_port, QN => n_1590);
   IF_ID_NPC_reg_4_inst : DFF_X1 port map( D => N6, CK => CLK, Q => 
                           IF_ID_NPC_4_port, QN => n_1591);
   ID_EX_NPC_reg_4_inst : DFF_X1 port map( D => N70, CK => CLK, Q => 
                           ID_EX_NPC_4_port, QN => n_1592);
   EX_MEM_NPC_reg_4_inst : DFF_X1 port map( D => N214, CK => CLK, Q => 
                           EX_MEM_NPC_4_port, QN => n_1593);
   MEM_WB_NPC_reg_4_inst : DFF_X1 port map( D => N317, CK => CLK, Q => 
                           MEM_WB_NPC_4_port, QN => n_1594);
   IF_ID_NPC_reg_5_inst : DFF_X1 port map( D => N7, CK => CLK, Q => 
                           IF_ID_NPC_5_port, QN => n_1595);
   ID_EX_NPC_reg_5_inst : DFF_X1 port map( D => N71, CK => CLK, Q => 
                           ID_EX_NPC_5_port, QN => n_1596);
   EX_MEM_NPC_reg_5_inst : DFF_X1 port map( D => N215, CK => CLK, Q => 
                           EX_MEM_NPC_5_port, QN => n_1597);
   MEM_WB_NPC_reg_5_inst : DFF_X1 port map( D => N318, CK => CLK, Q => 
                           MEM_WB_NPC_5_port, QN => n_1598);
   IF_ID_NPC_reg_6_inst : DFF_X1 port map( D => N8, CK => CLK, Q => 
                           IF_ID_NPC_6_port, QN => n_1599);
   ID_EX_NPC_reg_6_inst : DFF_X1 port map( D => N72, CK => CLK, Q => 
                           ID_EX_NPC_6_port, QN => n_1600);
   EX_MEM_NPC_reg_6_inst : DFF_X1 port map( D => N216, CK => CLK, Q => 
                           EX_MEM_NPC_6_port, QN => n_1601);
   MEM_WB_NPC_reg_6_inst : DFF_X1 port map( D => N319, CK => CLK, Q => 
                           MEM_WB_NPC_6_port, QN => n_1602);
   IF_ID_NPC_reg_7_inst : DFF_X1 port map( D => N9, CK => CLK, Q => 
                           IF_ID_NPC_7_port, QN => n_1603);
   ID_EX_NPC_reg_7_inst : DFF_X1 port map( D => N73, CK => CLK, Q => 
                           ID_EX_NPC_7_port, QN => n_1604);
   EX_MEM_NPC_reg_7_inst : DFF_X1 port map( D => N217, CK => CLK, Q => 
                           EX_MEM_NPC_7_port, QN => n_1605);
   MEM_WB_NPC_reg_7_inst : DFF_X1 port map( D => N320, CK => CLK, Q => 
                           MEM_WB_NPC_7_port, QN => n_1606);
   IF_ID_NPC_reg_8_inst : DFF_X1 port map( D => N10, CK => CLK, Q => 
                           IF_ID_NPC_8_port, QN => n_1607);
   ID_EX_NPC_reg_8_inst : DFF_X1 port map( D => N74, CK => CLK, Q => 
                           ID_EX_NPC_8_port, QN => n_1608);
   EX_MEM_NPC_reg_8_inst : DFF_X1 port map( D => N218, CK => CLK, Q => 
                           EX_MEM_NPC_8_port, QN => n_1609);
   MEM_WB_NPC_reg_8_inst : DFF_X1 port map( D => N321, CK => CLK, Q => 
                           MEM_WB_NPC_8_port, QN => n_1610);
   IF_ID_NPC_reg_9_inst : DFF_X1 port map( D => N11, CK => CLK, Q => 
                           IF_ID_NPC_9_port, QN => n_1611);
   ID_EX_NPC_reg_9_inst : DFF_X1 port map( D => N75, CK => CLK, Q => 
                           ID_EX_NPC_9_port, QN => n_1612);
   EX_MEM_NPC_reg_9_inst : DFF_X1 port map( D => N219, CK => CLK, Q => 
                           EX_MEM_NPC_9_port, QN => n_1613);
   MEM_WB_NPC_reg_9_inst : DFF_X1 port map( D => N322, CK => CLK, Q => 
                           MEM_WB_NPC_9_port, QN => n_1614);
   IF_ID_NPC_reg_10_inst : DFF_X1 port map( D => N12, CK => CLK, Q => 
                           IF_ID_NPC_10_port, QN => n_1615);
   ID_EX_NPC_reg_10_inst : DFF_X1 port map( D => N76, CK => CLK, Q => 
                           ID_EX_NPC_10_port, QN => n_1616);
   EX_MEM_NPC_reg_10_inst : DFF_X1 port map( D => N220, CK => CLK, Q => 
                           EX_MEM_NPC_10_port, QN => n_1617);
   MEM_WB_NPC_reg_10_inst : DFF_X1 port map( D => N323, CK => CLK, Q => 
                           MEM_WB_NPC_10_port, QN => n_1618);
   IF_ID_NPC_reg_11_inst : DFF_X1 port map( D => N13, CK => CLK, Q => 
                           IF_ID_NPC_11_port, QN => n_1619);
   ID_EX_NPC_reg_11_inst : DFF_X1 port map( D => N77, CK => CLK, Q => 
                           ID_EX_NPC_11_port, QN => n_1620);
   EX_MEM_NPC_reg_11_inst : DFF_X1 port map( D => N221, CK => CLK, Q => 
                           EX_MEM_NPC_11_port, QN => n_1621);
   MEM_WB_NPC_reg_11_inst : DFF_X1 port map( D => N324, CK => CLK, Q => 
                           MEM_WB_NPC_11_port, QN => n_1622);
   IF_ID_NPC_reg_12_inst : DFF_X1 port map( D => N14, CK => CLK, Q => 
                           IF_ID_NPC_12_port, QN => n_1623);
   ID_EX_NPC_reg_12_inst : DFF_X1 port map( D => N78, CK => CLK, Q => 
                           ID_EX_NPC_12_port, QN => n_1624);
   EX_MEM_NPC_reg_12_inst : DFF_X1 port map( D => N222, CK => CLK, Q => 
                           EX_MEM_NPC_12_port, QN => n_1625);
   MEM_WB_NPC_reg_12_inst : DFF_X1 port map( D => N325, CK => CLK, Q => 
                           MEM_WB_NPC_12_port, QN => n_1626);
   IF_ID_NPC_reg_13_inst : DFF_X1 port map( D => N15, CK => CLK, Q => 
                           IF_ID_NPC_13_port, QN => n_1627);
   ID_EX_NPC_reg_13_inst : DFF_X1 port map( D => N79, CK => CLK, Q => 
                           ID_EX_NPC_13_port, QN => n_1628);
   EX_MEM_NPC_reg_13_inst : DFF_X1 port map( D => N223, CK => CLK, Q => 
                           EX_MEM_NPC_13_port, QN => n_1629);
   MEM_WB_NPC_reg_13_inst : DFF_X1 port map( D => N326, CK => CLK, Q => 
                           MEM_WB_NPC_13_port, QN => n_1630);
   IF_ID_NPC_reg_14_inst : DFF_X1 port map( D => N16, CK => CLK, Q => 
                           IF_ID_NPC_14_port, QN => n_1631);
   ID_EX_NPC_reg_14_inst : DFF_X1 port map( D => N80, CK => CLK, Q => 
                           ID_EX_NPC_14_port, QN => n_1632);
   EX_MEM_NPC_reg_14_inst : DFF_X1 port map( D => N224, CK => CLK, Q => 
                           EX_MEM_NPC_14_port, QN => n_1633);
   MEM_WB_NPC_reg_14_inst : DFF_X1 port map( D => N327, CK => CLK, Q => 
                           MEM_WB_NPC_14_port, QN => n_1634);
   IF_ID_NPC_reg_15_inst : DFF_X1 port map( D => N17, CK => CLK, Q => 
                           IF_ID_NPC_15_port, QN => n_1635);
   ID_EX_NPC_reg_15_inst : DFF_X1 port map( D => N81, CK => CLK, Q => 
                           ID_EX_NPC_15_port, QN => n_1636);
   EX_MEM_NPC_reg_15_inst : DFF_X1 port map( D => N225, CK => CLK, Q => 
                           EX_MEM_NPC_15_port, QN => n_1637);
   MEM_WB_NPC_reg_15_inst : DFF_X1 port map( D => N328, CK => CLK, Q => 
                           MEM_WB_NPC_15_port, QN => n_1638);
   IF_ID_NPC_reg_16_inst : DFF_X1 port map( D => N18, CK => CLK, Q => 
                           IF_ID_NPC_16_port, QN => n_1639);
   ID_EX_NPC_reg_16_inst : DFF_X1 port map( D => N82, CK => CLK, Q => 
                           ID_EX_NPC_16_port, QN => n_1640);
   EX_MEM_NPC_reg_16_inst : DFF_X1 port map( D => N226, CK => CLK, Q => 
                           EX_MEM_NPC_16_port, QN => n_1641);
   MEM_WB_NPC_reg_16_inst : DFF_X1 port map( D => N329, CK => CLK, Q => 
                           MEM_WB_NPC_16_port, QN => n_1642);
   IF_ID_NPC_reg_17_inst : DFF_X1 port map( D => N19, CK => CLK, Q => 
                           IF_ID_NPC_17_port, QN => n_1643);
   ID_EX_NPC_reg_17_inst : DFF_X1 port map( D => N83, CK => CLK, Q => 
                           ID_EX_NPC_17_port, QN => n_1644);
   EX_MEM_NPC_reg_17_inst : DFF_X1 port map( D => N227, CK => CLK, Q => 
                           EX_MEM_NPC_17_port, QN => n_1645);
   MEM_WB_NPC_reg_17_inst : DFF_X1 port map( D => N330, CK => CLK, Q => 
                           MEM_WB_NPC_17_port, QN => n_1646);
   IF_ID_NPC_reg_18_inst : DFF_X1 port map( D => N20, CK => CLK, Q => 
                           IF_ID_NPC_18_port, QN => n_1647);
   ID_EX_NPC_reg_18_inst : DFF_X1 port map( D => N84, CK => CLK, Q => 
                           ID_EX_NPC_18_port, QN => n_1648);
   EX_MEM_NPC_reg_18_inst : DFF_X1 port map( D => N228, CK => CLK, Q => 
                           EX_MEM_NPC_18_port, QN => n_1649);
   MEM_WB_NPC_reg_18_inst : DFF_X1 port map( D => N331, CK => CLK, Q => 
                           MEM_WB_NPC_18_port, QN => n_1650);
   IF_ID_NPC_reg_19_inst : DFF_X1 port map( D => N21, CK => CLK, Q => 
                           IF_ID_NPC_19_port, QN => n_1651);
   ID_EX_NPC_reg_19_inst : DFF_X1 port map( D => N85, CK => CLK, Q => 
                           ID_EX_NPC_19_port, QN => n_1652);
   EX_MEM_NPC_reg_19_inst : DFF_X1 port map( D => N229, CK => CLK, Q => 
                           EX_MEM_NPC_19_port, QN => n_1653);
   MEM_WB_NPC_reg_19_inst : DFF_X1 port map( D => N332, CK => CLK, Q => 
                           MEM_WB_NPC_19_port, QN => n_1654);
   IF_ID_NPC_reg_20_inst : DFF_X1 port map( D => N22, CK => CLK, Q => 
                           IF_ID_NPC_20_port, QN => n_1655);
   ID_EX_NPC_reg_20_inst : DFF_X1 port map( D => N86, CK => CLK, Q => 
                           ID_EX_NPC_20_port, QN => n_1656);
   EX_MEM_NPC_reg_20_inst : DFF_X1 port map( D => N230, CK => CLK, Q => 
                           EX_MEM_NPC_20_port, QN => n_1657);
   MEM_WB_NPC_reg_20_inst : DFF_X1 port map( D => N333, CK => CLK, Q => 
                           MEM_WB_NPC_20_port, QN => n_1658);
   IF_ID_NPC_reg_21_inst : DFF_X1 port map( D => N23, CK => CLK, Q => 
                           IF_ID_NPC_21_port, QN => n_1659);
   ID_EX_NPC_reg_21_inst : DFF_X1 port map( D => N87, CK => CLK, Q => 
                           ID_EX_NPC_21_port, QN => n_1660);
   EX_MEM_NPC_reg_21_inst : DFF_X1 port map( D => N231, CK => CLK, Q => 
                           EX_MEM_NPC_21_port, QN => n_1661);
   MEM_WB_NPC_reg_21_inst : DFF_X1 port map( D => N334, CK => CLK, Q => 
                           MEM_WB_NPC_21_port, QN => n_1662);
   IF_ID_NPC_reg_22_inst : DFF_X1 port map( D => N24, CK => CLK, Q => 
                           IF_ID_NPC_22_port, QN => n_1663);
   ID_EX_NPC_reg_22_inst : DFF_X1 port map( D => N88, CK => CLK, Q => 
                           ID_EX_NPC_22_port, QN => n_1664);
   EX_MEM_NPC_reg_22_inst : DFF_X1 port map( D => N232, CK => CLK, Q => 
                           EX_MEM_NPC_22_port, QN => n_1665);
   MEM_WB_NPC_reg_22_inst : DFF_X1 port map( D => N335, CK => CLK, Q => 
                           MEM_WB_NPC_22_port, QN => n_1666);
   IF_ID_NPC_reg_23_inst : DFF_X1 port map( D => N25, CK => CLK, Q => 
                           IF_ID_NPC_23_port, QN => n_1667);
   ID_EX_NPC_reg_23_inst : DFF_X1 port map( D => N89, CK => CLK, Q => 
                           ID_EX_NPC_23_port, QN => n_1668);
   EX_MEM_NPC_reg_23_inst : DFF_X1 port map( D => N233, CK => CLK, Q => 
                           EX_MEM_NPC_23_port, QN => n_1669);
   MEM_WB_NPC_reg_23_inst : DFF_X1 port map( D => N336, CK => CLK, Q => 
                           MEM_WB_NPC_23_port, QN => n_1670);
   IF_ID_NPC_reg_24_inst : DFF_X1 port map( D => N26, CK => CLK, Q => 
                           IF_ID_NPC_24_port, QN => n_1671);
   ID_EX_NPC_reg_24_inst : DFF_X1 port map( D => N90, CK => CLK, Q => 
                           ID_EX_NPC_24_port, QN => n_1672);
   EX_MEM_NPC_reg_24_inst : DFF_X1 port map( D => N234, CK => CLK, Q => 
                           EX_MEM_NPC_24_port, QN => n_1673);
   MEM_WB_NPC_reg_24_inst : DFF_X1 port map( D => N337, CK => CLK, Q => 
                           MEM_WB_NPC_24_port, QN => n_1674);
   IF_ID_NPC_reg_25_inst : DFF_X1 port map( D => N27, CK => CLK, Q => 
                           IF_ID_NPC_25_port, QN => n_1675);
   ID_EX_NPC_reg_25_inst : DFF_X1 port map( D => N91, CK => CLK, Q => 
                           ID_EX_NPC_25_port, QN => n_1676);
   EX_MEM_NPC_reg_25_inst : DFF_X1 port map( D => N235, CK => CLK, Q => 
                           EX_MEM_NPC_25_port, QN => n_1677);
   MEM_WB_NPC_reg_25_inst : DFF_X1 port map( D => N338, CK => CLK, Q => 
                           MEM_WB_NPC_25_port, QN => n_1678);
   IF_ID_NPC_reg_26_inst : DFF_X1 port map( D => N28, CK => CLK, Q => 
                           IF_ID_NPC_26_port, QN => n_1679);
   ID_EX_NPC_reg_26_inst : DFF_X1 port map( D => N92, CK => CLK, Q => 
                           ID_EX_NPC_26_port, QN => n_1680);
   EX_MEM_NPC_reg_26_inst : DFF_X1 port map( D => N236, CK => CLK, Q => 
                           EX_MEM_NPC_26_port, QN => n_1681);
   MEM_WB_NPC_reg_26_inst : DFF_X1 port map( D => N339, CK => CLK, Q => 
                           MEM_WB_NPC_26_port, QN => n_1682);
   IF_ID_NPC_reg_27_inst : DFF_X1 port map( D => N29, CK => CLK, Q => 
                           IF_ID_NPC_27_port, QN => n_1683);
   ID_EX_NPC_reg_27_inst : DFF_X1 port map( D => N93, CK => CLK, Q => 
                           ID_EX_NPC_27_port, QN => n_1684);
   EX_MEM_NPC_reg_27_inst : DFF_X1 port map( D => N237, CK => CLK, Q => 
                           EX_MEM_NPC_27_port, QN => n_1685);
   MEM_WB_NPC_reg_27_inst : DFF_X1 port map( D => N340, CK => CLK, Q => 
                           MEM_WB_NPC_27_port, QN => n_1686);
   IF_ID_NPC_reg_28_inst : DFF_X1 port map( D => N30, CK => CLK, Q => 
                           IF_ID_NPC_28_port, QN => n_1687);
   ID_EX_NPC_reg_28_inst : DFF_X1 port map( D => N94, CK => CLK, Q => 
                           ID_EX_NPC_28_port, QN => n_1688);
   EX_MEM_NPC_reg_28_inst : DFF_X1 port map( D => N238, CK => CLK, Q => 
                           EX_MEM_NPC_28_port, QN => n_1689);
   MEM_WB_NPC_reg_28_inst : DFF_X1 port map( D => N341, CK => CLK, Q => 
                           MEM_WB_NPC_28_port, QN => n_1690);
   IF_ID_NPC_reg_29_inst : DFF_X1 port map( D => N31, CK => CLK, Q => 
                           IF_ID_NPC_29_port, QN => n_1691);
   ID_EX_NPC_reg_29_inst : DFF_X1 port map( D => N95, CK => CLK, Q => 
                           ID_EX_NPC_29_port, QN => n_1692);
   EX_MEM_NPC_reg_29_inst : DFF_X1 port map( D => N239, CK => CLK, Q => 
                           EX_MEM_NPC_29_port, QN => n_1693);
   MEM_WB_NPC_reg_29_inst : DFF_X1 port map( D => N342, CK => CLK, Q => 
                           MEM_WB_NPC_29_port, QN => n_1694);
   IF_ID_NPC_reg_30_inst : DFF_X1 port map( D => N32, CK => CLK, Q => 
                           IF_ID_NPC_30_port, QN => n_1695);
   ID_EX_NPC_reg_30_inst : DFF_X1 port map( D => N96, CK => CLK, Q => 
                           ID_EX_NPC_30_port, QN => n_1696);
   EX_MEM_NPC_reg_30_inst : DFF_X1 port map( D => N240, CK => CLK, Q => 
                           EX_MEM_NPC_30_port, QN => n_1697);
   MEM_WB_NPC_reg_30_inst : DFF_X1 port map( D => N343, CK => CLK, Q => 
                           MEM_WB_NPC_30_port, QN => n_1698);
   IF_ID_NPC_reg_31_inst : DFF_X1 port map( D => N33, CK => CLK, Q => 
                           IF_ID_NPC_31_port, QN => n_1699);
   ID_EX_NPC_reg_31_inst : DFF_X1 port map( D => N97, CK => CLK, Q => 
                           ID_EX_NPC_31_port, QN => n_1700);
   EX_MEM_NPC_reg_31_inst : DFF_X1 port map( D => N241, CK => CLK, Q => 
                           EX_MEM_NPC_31_port, QN => n_1701);
   MEM_WB_NPC_reg_31_inst : DFF_X1 port map( D => N344, CK => CLK, Q => 
                           MEM_WB_NPC_31_port, QN => n_1702);
   MEM_WB_ALU_OUTPUT_reg_31_inst : DFF_X1 port map( D => N377, CK => CLK, Q => 
                           MEM_WB_ALU_OUTPUT_31_port, QN => n_1703);
   PROGRAM_COUNTER : FFDR_N32 port map( CLK => CLK, RST => net31258, EN => 
                           PC_LATCH_EN, REGIN(31) => PC_BUS_31_port, REGIN(30) 
                           => PC_BUS_30_port, REGIN(29) => PC_BUS_29_port, 
                           REGIN(28) => PC_BUS_28_port, REGIN(27) => 
                           PC_BUS_27_port, REGIN(26) => PC_BUS_26_port, 
                           REGIN(25) => PC_BUS_25_port, REGIN(24) => 
                           PC_BUS_24_port, REGIN(23) => PC_BUS_23_port, 
                           REGIN(22) => PC_BUS_22_port, REGIN(21) => 
                           PC_BUS_21_port, REGIN(20) => PC_BUS_20_port, 
                           REGIN(19) => PC_BUS_19_port, REGIN(18) => 
                           PC_BUS_18_port, REGIN(17) => PC_BUS_17_port, 
                           REGIN(16) => PC_BUS_16_port, REGIN(15) => 
                           PC_BUS_15_port, REGIN(14) => PC_BUS_14_port, 
                           REGIN(13) => PC_BUS_13_port, REGIN(12) => 
                           PC_BUS_12_port, REGIN(11) => PC_BUS_11_port, 
                           REGIN(10) => PC_BUS_10_port, REGIN(9) => 
                           PC_BUS_9_port, REGIN(8) => PC_BUS_8_port, REGIN(7) 
                           => PC_BUS_7_port, REGIN(6) => PC_BUS_6_port, 
                           REGIN(5) => PC_BUS_5_port, REGIN(4) => PC_BUS_4_port
                           , REGIN(3) => PC_BUS_3_port, REGIN(2) => 
                           PC_BUS_2_port, REGIN(1) => PC_BUS_1_port, REGIN(0) 
                           => PC_BUS_0_port, REGOUT(31) => PC_OUT_31_port, 
                           REGOUT(30) => PC_OUT_30_port, REGOUT(29) => 
                           PC_OUT_29_port, REGOUT(28) => PC_OUT_28_port, 
                           REGOUT(27) => PC_OUT_27_port, REGOUT(26) => 
                           PC_OUT_26_port, REGOUT(25) => PC_OUT_25_port, 
                           REGOUT(24) => PC_OUT_24_port, REGOUT(23) => 
                           PC_OUT_23_port, REGOUT(22) => PC_OUT_22_port, 
                           REGOUT(21) => PC_OUT_21_port, REGOUT(20) => 
                           PC_OUT_20_port, REGOUT(19) => PC_OUT_19_port, 
                           REGOUT(18) => PC_OUT_18_port, REGOUT(17) => 
                           PC_OUT_17_port, REGOUT(16) => PC_OUT_16_port, 
                           REGOUT(15) => PC_OUT_15_port, REGOUT(14) => 
                           PC_OUT_14_port, REGOUT(13) => PC_OUT_13_port, 
                           REGOUT(12) => PC_OUT_12_port, REGOUT(11) => 
                           PC_OUT_11_port, REGOUT(10) => PC_OUT_10_port, 
                           REGOUT(9) => PC_OUT_9_port, REGOUT(8) => 
                           PC_OUT_8_port, REGOUT(7) => PC_OUT_7_port, REGOUT(6)
                           => PC_OUT_6_port, REGOUT(5) => PC_OUT_5_port, 
                           REGOUT(4) => PC_OUT_4_port, REGOUT(3) => 
                           PC_OUT_3_port, REGOUT(2) => PC_OUT_2_port, REGOUT(1)
                           => PC_OUT_1_port, REGOUT(0) => PC_OUT_0_port);
   PC_MUX : MUX21_N32_4 port map( A(31) => NPC_BUS_31_port, A(30) => 
                           NPC_BUS_30_port, A(29) => NPC_BUS_29_port, A(28) => 
                           NPC_BUS_28_port, A(27) => NPC_BUS_27_port, A(26) => 
                           NPC_BUS_26_port, A(25) => NPC_BUS_25_port, A(24) => 
                           NPC_BUS_24_port, A(23) => NPC_BUS_23_port, A(22) => 
                           NPC_BUS_22_port, A(21) => NPC_BUS_21_port, A(20) => 
                           NPC_BUS_20_port, A(19) => NPC_BUS_19_port, A(18) => 
                           NPC_BUS_18_port, A(17) => NPC_BUS_17_port, A(16) => 
                           NPC_BUS_16_port, A(15) => NPC_BUS_15_port, A(14) => 
                           NPC_BUS_14_port, A(13) => NPC_BUS_13_port, A(12) => 
                           NPC_BUS_12_port, A(11) => NPC_BUS_11_port, A(10) => 
                           NPC_BUS_10_port, A(9) => NPC_BUS_9_port, A(8) => 
                           NPC_BUS_8_port, A(7) => NPC_BUS_7_port, A(6) => 
                           NPC_BUS_6_port, A(5) => NPC_BUS_5_port, A(4) => 
                           NPC_BUS_4_port, A(3) => NPC_BUS_3_port, A(2) => 
                           NPC_BUS_2_port, A(1) => NPC_BUS_1_port, A(0) => 
                           NPC_BUS_0_port, B(31) => ALU_OUT_31_port, B(30) => 
                           ALU_OUT_30_port, B(29) => ALU_OUT_29_port, B(28) => 
                           ALU_OUT_28_port, B(27) => ALU_OUT_27_port, B(26) => 
                           ALU_OUT_26_port, B(25) => ALU_OUT_25_port, B(24) => 
                           ALU_OUT_24_port, B(23) => ALU_OUT_23_port, B(22) => 
                           ALU_OUT_22_port, B(21) => ALU_OUT_21_port, B(20) => 
                           ALU_OUT_20_port, B(19) => ALU_OUT_19_port, B(18) => 
                           ALU_OUT_18_port, B(17) => ALU_OUT_17_port, B(16) => 
                           ALU_OUT_16_port, B(15) => ALU_OUT_15_port, B(14) => 
                           ALU_OUT_14_port, B(13) => ALU_OUT_13_port, B(12) => 
                           ALU_OUT_12_port, B(11) => ALU_OUT_11_port, B(10) => 
                           ALU_OUT_10_port, B(9) => ALU_OUT_9_port, B(8) => 
                           ALU_OUT_8_port, B(7) => ALU_OUT_7_port, B(6) => 
                           ALU_OUT_6_port, B(5) => ALU_OUT_5_port, B(4) => 
                           ALU_OUT_4_port, B(3) => ALU_OUT_3_port, B(2) => 
                           ALU_OUT_2_port, B(1) => ALU_OUT_1_port, B(0) => 
                           ALU_OUT_0_port, S => n19_port, Y(31) => 
                           PC_BUS_31_port, Y(30) => PC_BUS_30_port, Y(29) => 
                           PC_BUS_29_port, Y(28) => PC_BUS_28_port, Y(27) => 
                           PC_BUS_27_port, Y(26) => PC_BUS_26_port, Y(25) => 
                           PC_BUS_25_port, Y(24) => PC_BUS_24_port, Y(23) => 
                           PC_BUS_23_port, Y(22) => PC_BUS_22_port, Y(21) => 
                           PC_BUS_21_port, Y(20) => PC_BUS_20_port, Y(19) => 
                           PC_BUS_19_port, Y(18) => PC_BUS_18_port, Y(17) => 
                           PC_BUS_17_port, Y(16) => PC_BUS_16_port, Y(15) => 
                           PC_BUS_15_port, Y(14) => PC_BUS_14_port, Y(13) => 
                           PC_BUS_13_port, Y(12) => PC_BUS_12_port, Y(11) => 
                           PC_BUS_11_port, Y(10) => PC_BUS_10_port, Y(9) => 
                           PC_BUS_9_port, Y(8) => PC_BUS_8_port, Y(7) => 
                           PC_BUS_7_port, Y(6) => PC_BUS_6_port, Y(5) => 
                           PC_BUS_5_port, Y(4) => PC_BUS_4_port, Y(3) => 
                           PC_BUS_3_port, Y(2) => PC_BUS_2_port, Y(1) => 
                           PC_BUS_1_port, Y(0) => PC_BUS_0_port);
   NEXT_PROGRAM_COUNTER : LDR_N32_6 port map( RST => net31258, EN => 
                           NPC_LATCH_EN, REGIN(31) => PC_BUS_31_port, REGIN(30)
                           => PC_BUS_30_port, REGIN(29) => PC_BUS_29_port, 
                           REGIN(28) => PC_BUS_28_port, REGIN(27) => 
                           PC_BUS_27_port, REGIN(26) => PC_BUS_26_port, 
                           REGIN(25) => PC_BUS_25_port, REGIN(24) => 
                           PC_BUS_24_port, REGIN(23) => PC_BUS_23_port, 
                           REGIN(22) => PC_BUS_22_port, REGIN(21) => 
                           PC_BUS_21_port, REGIN(20) => PC_BUS_20_port, 
                           REGIN(19) => PC_BUS_19_port, REGIN(18) => 
                           PC_BUS_18_port, REGIN(17) => PC_BUS_17_port, 
                           REGIN(16) => PC_BUS_16_port, REGIN(15) => 
                           PC_BUS_15_port, REGIN(14) => PC_BUS_14_port, 
                           REGIN(13) => PC_BUS_13_port, REGIN(12) => 
                           PC_BUS_12_port, REGIN(11) => PC_BUS_11_port, 
                           REGIN(10) => PC_BUS_10_port, REGIN(9) => 
                           PC_BUS_9_port, REGIN(8) => PC_BUS_8_port, REGIN(7) 
                           => PC_BUS_7_port, REGIN(6) => PC_BUS_6_port, 
                           REGIN(5) => PC_BUS_5_port, REGIN(4) => PC_BUS_4_port
                           , REGIN(3) => PC_BUS_3_port, REGIN(2) => 
                           PC_BUS_2_port, REGIN(1) => PC_BUS_1_port, REGIN(0) 
                           => PC_BUS_0_port, REGOUT(31) => 
                           IF_ID_NPC_NEXT_31_port, REGOUT(30) => 
                           IF_ID_NPC_NEXT_30_port, REGOUT(29) => 
                           IF_ID_NPC_NEXT_29_port, REGOUT(28) => 
                           IF_ID_NPC_NEXT_28_port, REGOUT(27) => 
                           IF_ID_NPC_NEXT_27_port, REGOUT(26) => 
                           IF_ID_NPC_NEXT_26_port, REGOUT(25) => 
                           IF_ID_NPC_NEXT_25_port, REGOUT(24) => 
                           IF_ID_NPC_NEXT_24_port, REGOUT(23) => 
                           IF_ID_NPC_NEXT_23_port, REGOUT(22) => 
                           IF_ID_NPC_NEXT_22_port, REGOUT(21) => 
                           IF_ID_NPC_NEXT_21_port, REGOUT(20) => 
                           IF_ID_NPC_NEXT_20_port, REGOUT(19) => 
                           IF_ID_NPC_NEXT_19_port, REGOUT(18) => 
                           IF_ID_NPC_NEXT_18_port, REGOUT(17) => 
                           IF_ID_NPC_NEXT_17_port, REGOUT(16) => 
                           IF_ID_NPC_NEXT_16_port, REGOUT(15) => 
                           IF_ID_NPC_NEXT_15_port, REGOUT(14) => 
                           IF_ID_NPC_NEXT_14_port, REGOUT(13) => 
                           IF_ID_NPC_NEXT_13_port, REGOUT(12) => 
                           IF_ID_NPC_NEXT_12_port, REGOUT(11) => 
                           IF_ID_NPC_NEXT_11_port, REGOUT(10) => 
                           IF_ID_NPC_NEXT_10_port, REGOUT(9) => 
                           IF_ID_NPC_NEXT_9_port, REGOUT(8) => 
                           IF_ID_NPC_NEXT_8_port, REGOUT(7) => 
                           IF_ID_NPC_NEXT_7_port, REGOUT(6) => 
                           IF_ID_NPC_NEXT_6_port, REGOUT(5) => 
                           IF_ID_NPC_NEXT_5_port, REGOUT(4) => 
                           IF_ID_NPC_NEXT_4_port, REGOUT(3) => 
                           IF_ID_NPC_NEXT_3_port, REGOUT(2) => 
                           IF_ID_NPC_NEXT_2_port, REGOUT(1) => 
                           IF_ID_NPC_NEXT_1_port, REGOUT(0) => 
                           IF_ID_NPC_NEXT_0_port);
   INSTRUCTION_REGISTER : LDR_N32_5 port map( RST => net31258, EN => 
                           IR_LATCH_EN, REGIN(31) => IR_IN(31), REGIN(30) => 
                           IR_IN(30), REGIN(29) => IR_IN(29), REGIN(28) => 
                           IR_IN(28), REGIN(27) => IR_IN(27), REGIN(26) => 
                           IR_IN(26), REGIN(25) => IR_IN(25), REGIN(24) => 
                           IR_IN(24), REGIN(23) => IR_IN(23), REGIN(22) => 
                           IR_IN(22), REGIN(21) => IR_IN(21), REGIN(20) => 
                           IR_IN(20), REGIN(19) => IR_IN(19), REGIN(18) => 
                           IR_IN(18), REGIN(17) => IR_IN(17), REGIN(16) => 
                           IR_IN(16), REGIN(15) => IR_IN(15), REGIN(14) => 
                           IR_IN(14), REGIN(13) => IR_IN(13), REGIN(12) => 
                           IR_IN(12), REGIN(11) => IR_IN(11), REGIN(10) => 
                           IR_IN(10), REGIN(9) => IR_IN(9), REGIN(8) => 
                           IR_IN(8), REGIN(7) => IR_IN(7), REGIN(6) => IR_IN(6)
                           , REGIN(5) => IR_IN(5), REGIN(4) => IR_IN(4), 
                           REGIN(3) => IR_IN(3), REGIN(2) => IR_IN(2), REGIN(1)
                           => IR_IN(1), REGIN(0) => IR_IN(0), REGOUT(31) => 
                           IR_OUT_31_port, REGOUT(30) => IR_OUT_30_port, 
                           REGOUT(29) => IR_OUT_29_port, REGOUT(28) => 
                           IR_OUT_28_port, REGOUT(27) => IR_OUT_27_port, 
                           REGOUT(26) => IR_OUT_26_port, REGOUT(25) => 
                           IR_OUT_25_port, REGOUT(24) => IR_OUT_24_port, 
                           REGOUT(23) => IR_OUT_23_port, REGOUT(22) => 
                           IR_OUT_22_port, REGOUT(21) => IR_OUT_21_port, 
                           REGOUT(20) => IR_OUT_20_port, REGOUT(19) => 
                           IR_OUT_19_port, REGOUT(18) => IR_OUT_18_port, 
                           REGOUT(17) => IR_OUT_17_port, REGOUT(16) => 
                           IR_OUT_16_port, REGOUT(15) => IR_OUT_15_port, 
                           REGOUT(14) => IR_OUT_14_port, REGOUT(13) => 
                           IR_OUT_13_port, REGOUT(12) => IR_OUT_12_port, 
                           REGOUT(11) => IR_OUT_11_port, REGOUT(10) => 
                           IR_OUT_10_port, REGOUT(9) => IR_OUT_9_port, 
                           REGOUT(8) => IR_OUT_8_port, REGOUT(7) => 
                           IR_OUT_7_port, REGOUT(6) => IR_OUT_6_port, REGOUT(5)
                           => IR_OUT_5_port, REGOUT(4) => IR_OUT_4_port, 
                           REGOUT(3) => IR_OUT_3_port, REGOUT(2) => 
                           IR_OUT_2_port, REGOUT(1) => IR_OUT_1_port, REGOUT(0)
                           => IR_OUT_0_port);
   REGISTER_FILE : RF_N32_NA5 port map( RST => net31258, EN => X_Logic1_port, 
                           EN_RD1 => X_Logic1_port, EN_RD2 => X_Logic1_port, 
                           EN_WR => MEM_WB_RF_WE, ADD_RD1(4) => n3_port, 
                           ADD_RD1(3) => ID_EX_RS1_NEXT_3_port, ADD_RD1(2) => 
                           ID_EX_RS1_NEXT_2_port, ADD_RD1(1) => 
                           ID_EX_RS1_NEXT_1_port, ADD_RD1(0) => n2_port, 
                           ADD_RD2(4) => n13_port, ADD_RD2(3) => net31024, 
                           ADD_RD2(2) => net31028, ADD_RD2(1) => n12_port, 
                           ADD_RD2(0) => n11_port, ADD_WR(4) => 
                           MEM_WB_RD_4_port, ADD_WR(3) => MEM_WB_RD_3_port, 
                           ADD_WR(2) => MEM_WB_RD_2_port, ADD_WR(1) => 
                           MEM_WB_RD_1_port, ADD_WR(0) => MEM_WB_RD_0_port, 
                           DATAIN(31) => JAL_MUX_OUT_31_port, DATAIN(30) => 
                           JAL_MUX_OUT_30_port, DATAIN(29) => 
                           JAL_MUX_OUT_29_port, DATAIN(28) => 
                           JAL_MUX_OUT_28_port, DATAIN(27) => 
                           JAL_MUX_OUT_27_port, DATAIN(26) => 
                           JAL_MUX_OUT_26_port, DATAIN(25) => 
                           JAL_MUX_OUT_25_port, DATAIN(24) => 
                           JAL_MUX_OUT_24_port, DATAIN(23) => 
                           JAL_MUX_OUT_23_port, DATAIN(22) => 
                           JAL_MUX_OUT_22_port, DATAIN(21) => 
                           JAL_MUX_OUT_21_port, DATAIN(20) => 
                           JAL_MUX_OUT_20_port, DATAIN(19) => 
                           JAL_MUX_OUT_19_port, DATAIN(18) => 
                           JAL_MUX_OUT_18_port, DATAIN(17) => 
                           JAL_MUX_OUT_17_port, DATAIN(16) => 
                           JAL_MUX_OUT_16_port, DATAIN(15) => 
                           JAL_MUX_OUT_15_port, DATAIN(14) => 
                           JAL_MUX_OUT_14_port, DATAIN(13) => 
                           JAL_MUX_OUT_13_port, DATAIN(12) => 
                           JAL_MUX_OUT_12_port, DATAIN(11) => 
                           JAL_MUX_OUT_11_port, DATAIN(10) => 
                           JAL_MUX_OUT_10_port, DATAIN(9) => JAL_MUX_OUT_9_port
                           , DATAIN(8) => JAL_MUX_OUT_8_port, DATAIN(7) => 
                           JAL_MUX_OUT_7_port, DATAIN(6) => JAL_MUX_OUT_6_port,
                           DATAIN(5) => JAL_MUX_OUT_5_port, DATAIN(4) => 
                           JAL_MUX_OUT_4_port, DATAIN(3) => JAL_MUX_OUT_3_port,
                           DATAIN(2) => JAL_MUX_OUT_2_port, DATAIN(1) => 
                           JAL_MUX_OUT_1_port, DATAIN(0) => JAL_MUX_OUT_0_port,
                           OUT1(31) => RF_OUT1_31_port, OUT1(30) => 
                           RF_OUT1_30_port, OUT1(29) => RF_OUT1_29_port, 
                           OUT1(28) => RF_OUT1_28_port, OUT1(27) => 
                           RF_OUT1_27_port, OUT1(26) => RF_OUT1_26_port, 
                           OUT1(25) => RF_OUT1_25_port, OUT1(24) => 
                           RF_OUT1_24_port, OUT1(23) => RF_OUT1_23_port, 
                           OUT1(22) => RF_OUT1_22_port, OUT1(21) => 
                           RF_OUT1_21_port, OUT1(20) => RF_OUT1_20_port, 
                           OUT1(19) => RF_OUT1_19_port, OUT1(18) => 
                           RF_OUT1_18_port, OUT1(17) => RF_OUT1_17_port, 
                           OUT1(16) => RF_OUT1_16_port, OUT1(15) => 
                           RF_OUT1_15_port, OUT1(14) => RF_OUT1_14_port, 
                           OUT1(13) => RF_OUT1_13_port, OUT1(12) => 
                           RF_OUT1_12_port, OUT1(11) => RF_OUT1_11_port, 
                           OUT1(10) => RF_OUT1_10_port, OUT1(9) => 
                           RF_OUT1_9_port, OUT1(8) => RF_OUT1_8_port, OUT1(7) 
                           => RF_OUT1_7_port, OUT1(6) => RF_OUT1_6_port, 
                           OUT1(5) => RF_OUT1_5_port, OUT1(4) => RF_OUT1_4_port
                           , OUT1(3) => RF_OUT1_3_port, OUT1(2) => 
                           RF_OUT1_2_port, OUT1(1) => RF_OUT1_1_port, OUT1(0) 
                           => RF_OUT1_0_port, OUT2(31) => RF_OUT2_31_port, 
                           OUT2(30) => RF_OUT2_30_port, OUT2(29) => 
                           RF_OUT2_29_port, OUT2(28) => RF_OUT2_28_port, 
                           OUT2(27) => RF_OUT2_27_port, OUT2(26) => 
                           RF_OUT2_26_port, OUT2(25) => RF_OUT2_25_port, 
                           OUT2(24) => RF_OUT2_24_port, OUT2(23) => 
                           RF_OUT2_23_port, OUT2(22) => RF_OUT2_22_port, 
                           OUT2(21) => RF_OUT2_21_port, OUT2(20) => 
                           RF_OUT2_20_port, OUT2(19) => RF_OUT2_19_port, 
                           OUT2(18) => RF_OUT2_18_port, OUT2(17) => 
                           RF_OUT2_17_port, OUT2(16) => RF_OUT2_16_port, 
                           OUT2(15) => RF_OUT2_15_port, OUT2(14) => 
                           RF_OUT2_14_port, OUT2(13) => RF_OUT2_13_port, 
                           OUT2(12) => RF_OUT2_12_port, OUT2(11) => 
                           RF_OUT2_11_port, OUT2(10) => RF_OUT2_10_port, 
                           OUT2(9) => RF_OUT2_9_port, OUT2(8) => RF_OUT2_8_port
                           , OUT2(7) => RF_OUT2_7_port, OUT2(6) => 
                           RF_OUT2_6_port, OUT2(5) => RF_OUT2_5_port, OUT2(4) 
                           => RF_OUT2_4_port, OUT2(3) => RF_OUT2_3_port, 
                           OUT2(2) => RF_OUT2_2_port, OUT2(1) => RF_OUT2_1_port
                           , OUT2(0) => RF_OUT2_0_port);
   SIGN_EXTEND : SIGNEX_N32_OPC6_REG5 port map( INSTR(31) => n8_port, INSTR(30)
                           => n6_port, INSTR(29) => n10_port, INSTR(28) => 
                           IF_ID_IR_28_port, INSTR(27) => n17_port, INSTR(26) 
                           => n15_port, INSTR(25) => IF_ID_IR_25_port, 
                           INSTR(24) => IF_ID_IR_24_port, INSTR(23) => 
                           IF_ID_IR_23_port, INSTR(22) => IF_ID_IR_22_port, 
                           INSTR(21) => IF_ID_IR_21_port, INSTR(20) => 
                           IF_ID_IR_20_port, INSTR(19) => IF_ID_IR_19_port, 
                           INSTR(18) => IF_ID_IR_18_port, INSTR(17) => 
                           IF_ID_IR_17_port, INSTR(16) => IF_ID_IR_16_port, 
                           INSTR(15) => IF_ID_IR_15_port, INSTR(14) => 
                           IF_ID_IR_14_port, INSTR(13) => IF_ID_IR_13_port, 
                           INSTR(12) => IF_ID_IR_12_port, INSTR(11) => 
                           IF_ID_IR_11_port, INSTR(10) => IF_ID_IR_10_port, 
                           INSTR(9) => IF_ID_IR_9_port, INSTR(8) => 
                           IF_ID_IR_8_port, INSTR(7) => IF_ID_IR_7_port, 
                           INSTR(6) => IF_ID_IR_6_port, INSTR(5) => 
                           IF_ID_IR_5_port, INSTR(4) => IF_ID_IR_4_port, 
                           INSTR(3) => IF_ID_IR_3_port, INSTR(2) => 
                           IF_ID_IR_2_port, INSTR(1) => IF_ID_IR_1_port, 
                           INSTR(0) => IF_ID_IR_0_port, IMM(31) => 
                           IMM_OUT_31_port, IMM(30) => IMM_OUT_30_port, IMM(29)
                           => IMM_OUT_29_port, IMM(28) => IMM_OUT_28_port, 
                           IMM(27) => IMM_OUT_27_port, IMM(26) => 
                           IMM_OUT_26_port, IMM(25) => IMM_OUT_25_port, IMM(24)
                           => IMM_OUT_24_port, IMM(23) => IMM_OUT_23_port, 
                           IMM(22) => IMM_OUT_22_port, IMM(21) => 
                           IMM_OUT_21_port, IMM(20) => IMM_OUT_20_port, IMM(19)
                           => IMM_OUT_19_port, IMM(18) => IMM_OUT_18_port, 
                           IMM(17) => IMM_OUT_17_port, IMM(16) => 
                           IMM_OUT_16_port, IMM(15) => IMM_OUT_15_port, IMM(14)
                           => IMM_OUT_14_port, IMM(13) => IMM_OUT_13_port, 
                           IMM(12) => IMM_OUT_12_port, IMM(11) => 
                           IMM_OUT_11_port, IMM(10) => IMM_OUT_10_port, IMM(9) 
                           => IMM_OUT_9_port, IMM(8) => IMM_OUT_8_port, IMM(7) 
                           => IMM_OUT_7_port, IMM(6) => IMM_OUT_6_port, IMM(5) 
                           => IMM_OUT_5_port, IMM(4) => IMM_OUT_4_port, IMM(3) 
                           => IMM_OUT_3_port, IMM(2) => IMM_OUT_2_port, IMM(1) 
                           => IMM_OUT_1_port, IMM(0) => IMM_OUT_0_port);
   REGISTER_ADDRESSER : REGADDR_N32_OPC6_REG5 port map( INSTR(31) => 
                           IF_ID_IR_31_port, INSTR(30) => IF_ID_IR_30_port, 
                           INSTR(29) => IF_ID_IR_29_port, INSTR(28) => 
                           IF_ID_IR_28_port, INSTR(27) => IF_ID_IR_27_port, 
                           INSTR(26) => IF_ID_IR_26_port, INSTR(25) => 
                           IF_ID_IR_25_port, INSTR(24) => IF_ID_IR_24_port, 
                           INSTR(23) => IF_ID_IR_23_port, INSTR(22) => 
                           IF_ID_IR_22_port, INSTR(21) => IF_ID_IR_21_port, 
                           INSTR(20) => IF_ID_IR_20_port, INSTR(19) => 
                           IF_ID_IR_19_port, INSTR(18) => IF_ID_IR_18_port, 
                           INSTR(17) => IF_ID_IR_17_port, INSTR(16) => 
                           IF_ID_IR_16_port, INSTR(15) => IF_ID_IR_15_port, 
                           INSTR(14) => IF_ID_IR_14_port, INSTR(13) => 
                           IF_ID_IR_13_port, INSTR(12) => IF_ID_IR_12_port, 
                           INSTR(11) => IF_ID_IR_11_port, INSTR(10) => 
                           IF_ID_IR_10_port, INSTR(9) => IF_ID_IR_9_port, 
                           INSTR(8) => IF_ID_IR_8_port, INSTR(7) => 
                           IF_ID_IR_7_port, INSTR(6) => IF_ID_IR_6_port, 
                           INSTR(5) => IF_ID_IR_5_port, INSTR(4) => 
                           IF_ID_IR_4_port, INSTR(3) => IF_ID_IR_3_port, 
                           INSTR(2) => IF_ID_IR_2_port, INSTR(1) => 
                           IF_ID_IR_1_port, INSTR(0) => IF_ID_IR_0_port, RS1(4)
                           => ID_EX_RS1_NEXT_4_port, RS1(3) => 
                           ID_EX_RS1_NEXT_3_port, RS1(2) => 
                           ID_EX_RS1_NEXT_2_port, RS1(1) => 
                           ID_EX_RS1_NEXT_1_port, RS1(0) => 
                           ID_EX_RS1_NEXT_0_port, RS2(4) => 
                           ID_EX_RS2_NEXT_4_port, RS2(3) => 
                           ID_EX_RS2_NEXT_3_port, RS2(2) => 
                           ID_EX_RS2_NEXT_2_port, RS2(1) => 
                           ID_EX_RS2_NEXT_1_port, RS2(0) => 
                           ID_EX_RS2_NEXT_0_port, RD(4) => ID_EX_RD_NEXT_4_port
                           , RD(3) => ID_EX_RD_NEXT_3_port, RD(2) => 
                           ID_EX_RD_NEXT_2_port, RD(1) => ID_EX_RD_NEXT_1_port,
                           RD(0) => ID_EX_RD_NEXT_0_port);
   LATCH_RF1 : LDR_N32_4 port map( RST => net31258, EN => RegA_LATCH_EN, 
                           REGIN(31) => RF_OUT1_31_port, REGIN(30) => 
                           RF_OUT1_30_port, REGIN(29) => RF_OUT1_29_port, 
                           REGIN(28) => RF_OUT1_28_port, REGIN(27) => 
                           RF_OUT1_27_port, REGIN(26) => RF_OUT1_26_port, 
                           REGIN(25) => RF_OUT1_25_port, REGIN(24) => 
                           RF_OUT1_24_port, REGIN(23) => RF_OUT1_23_port, 
                           REGIN(22) => RF_OUT1_22_port, REGIN(21) => 
                           RF_OUT1_21_port, REGIN(20) => RF_OUT1_20_port, 
                           REGIN(19) => RF_OUT1_19_port, REGIN(18) => 
                           RF_OUT1_18_port, REGIN(17) => RF_OUT1_17_port, 
                           REGIN(16) => RF_OUT1_16_port, REGIN(15) => 
                           RF_OUT1_15_port, REGIN(14) => RF_OUT1_14_port, 
                           REGIN(13) => RF_OUT1_13_port, REGIN(12) => 
                           RF_OUT1_12_port, REGIN(11) => RF_OUT1_11_port, 
                           REGIN(10) => RF_OUT1_10_port, REGIN(9) => 
                           RF_OUT1_9_port, REGIN(8) => RF_OUT1_8_port, REGIN(7)
                           => RF_OUT1_7_port, REGIN(6) => RF_OUT1_6_port, 
                           REGIN(5) => RF_OUT1_5_port, REGIN(4) => 
                           RF_OUT1_4_port, REGIN(3) => RF_OUT1_3_port, REGIN(2)
                           => RF_OUT1_2_port, REGIN(1) => RF_OUT1_1_port, 
                           REGIN(0) => RF_OUT1_0_port, REGOUT(31) => 
                           ID_EX_RF_OUT1_NEXT_31_port, REGOUT(30) => 
                           ID_EX_RF_OUT1_NEXT_30_port, REGOUT(29) => 
                           ID_EX_RF_OUT1_NEXT_29_port, REGOUT(28) => 
                           ID_EX_RF_OUT1_NEXT_28_port, REGOUT(27) => 
                           ID_EX_RF_OUT1_NEXT_27_port, REGOUT(26) => 
                           ID_EX_RF_OUT1_NEXT_26_port, REGOUT(25) => 
                           ID_EX_RF_OUT1_NEXT_25_port, REGOUT(24) => 
                           ID_EX_RF_OUT1_NEXT_24_port, REGOUT(23) => 
                           ID_EX_RF_OUT1_NEXT_23_port, REGOUT(22) => 
                           ID_EX_RF_OUT1_NEXT_22_port, REGOUT(21) => 
                           ID_EX_RF_OUT1_NEXT_21_port, REGOUT(20) => 
                           ID_EX_RF_OUT1_NEXT_20_port, REGOUT(19) => 
                           ID_EX_RF_OUT1_NEXT_19_port, REGOUT(18) => 
                           ID_EX_RF_OUT1_NEXT_18_port, REGOUT(17) => 
                           ID_EX_RF_OUT1_NEXT_17_port, REGOUT(16) => 
                           ID_EX_RF_OUT1_NEXT_16_port, REGOUT(15) => 
                           ID_EX_RF_OUT1_NEXT_15_port, REGOUT(14) => 
                           ID_EX_RF_OUT1_NEXT_14_port, REGOUT(13) => 
                           ID_EX_RF_OUT1_NEXT_13_port, REGOUT(12) => 
                           ID_EX_RF_OUT1_NEXT_12_port, REGOUT(11) => 
                           ID_EX_RF_OUT1_NEXT_11_port, REGOUT(10) => 
                           ID_EX_RF_OUT1_NEXT_10_port, REGOUT(9) => 
                           ID_EX_RF_OUT1_NEXT_9_port, REGOUT(8) => 
                           ID_EX_RF_OUT1_NEXT_8_port, REGOUT(7) => 
                           ID_EX_RF_OUT1_NEXT_7_port, REGOUT(6) => 
                           ID_EX_RF_OUT1_NEXT_6_port, REGOUT(5) => 
                           ID_EX_RF_OUT1_NEXT_5_port, REGOUT(4) => 
                           ID_EX_RF_OUT1_NEXT_4_port, REGOUT(3) => 
                           ID_EX_RF_OUT1_NEXT_3_port, REGOUT(2) => 
                           ID_EX_RF_OUT1_NEXT_2_port, REGOUT(1) => 
                           ID_EX_RF_OUT1_NEXT_1_port, REGOUT(0) => 
                           ID_EX_RF_OUT1_NEXT_0_port);
   LATCH_RF2 : LDR_N32_3 port map( RST => net31258, EN => RegB_LATCH_EN, 
                           REGIN(31) => RF_OUT2_31_port, REGIN(30) => 
                           RF_OUT2_30_port, REGIN(29) => RF_OUT2_29_port, 
                           REGIN(28) => RF_OUT2_28_port, REGIN(27) => 
                           RF_OUT2_27_port, REGIN(26) => RF_OUT2_26_port, 
                           REGIN(25) => RF_OUT2_25_port, REGIN(24) => 
                           RF_OUT2_24_port, REGIN(23) => RF_OUT2_23_port, 
                           REGIN(22) => RF_OUT2_22_port, REGIN(21) => 
                           RF_OUT2_21_port, REGIN(20) => RF_OUT2_20_port, 
                           REGIN(19) => RF_OUT2_19_port, REGIN(18) => 
                           RF_OUT2_18_port, REGIN(17) => RF_OUT2_17_port, 
                           REGIN(16) => RF_OUT2_16_port, REGIN(15) => 
                           RF_OUT2_15_port, REGIN(14) => RF_OUT2_14_port, 
                           REGIN(13) => RF_OUT2_13_port, REGIN(12) => 
                           RF_OUT2_12_port, REGIN(11) => RF_OUT2_11_port, 
                           REGIN(10) => RF_OUT2_10_port, REGIN(9) => 
                           RF_OUT2_9_port, REGIN(8) => RF_OUT2_8_port, REGIN(7)
                           => RF_OUT2_7_port, REGIN(6) => RF_OUT2_6_port, 
                           REGIN(5) => RF_OUT2_5_port, REGIN(4) => 
                           RF_OUT2_4_port, REGIN(3) => RF_OUT2_3_port, REGIN(2)
                           => RF_OUT2_2_port, REGIN(1) => RF_OUT2_1_port, 
                           REGIN(0) => RF_OUT2_0_port, REGOUT(31) => 
                           ID_EX_RF_OUT2_NEXT_31_port, REGOUT(30) => 
                           ID_EX_RF_OUT2_NEXT_30_port, REGOUT(29) => 
                           ID_EX_RF_OUT2_NEXT_29_port, REGOUT(28) => 
                           ID_EX_RF_OUT2_NEXT_28_port, REGOUT(27) => 
                           ID_EX_RF_OUT2_NEXT_27_port, REGOUT(26) => 
                           ID_EX_RF_OUT2_NEXT_26_port, REGOUT(25) => 
                           ID_EX_RF_OUT2_NEXT_25_port, REGOUT(24) => 
                           ID_EX_RF_OUT2_NEXT_24_port, REGOUT(23) => 
                           ID_EX_RF_OUT2_NEXT_23_port, REGOUT(22) => 
                           ID_EX_RF_OUT2_NEXT_22_port, REGOUT(21) => 
                           ID_EX_RF_OUT2_NEXT_21_port, REGOUT(20) => 
                           ID_EX_RF_OUT2_NEXT_20_port, REGOUT(19) => 
                           ID_EX_RF_OUT2_NEXT_19_port, REGOUT(18) => 
                           ID_EX_RF_OUT2_NEXT_18_port, REGOUT(17) => 
                           ID_EX_RF_OUT2_NEXT_17_port, REGOUT(16) => 
                           ID_EX_RF_OUT2_NEXT_16_port, REGOUT(15) => 
                           ID_EX_RF_OUT2_NEXT_15_port, REGOUT(14) => 
                           ID_EX_RF_OUT2_NEXT_14_port, REGOUT(13) => 
                           ID_EX_RF_OUT2_NEXT_13_port, REGOUT(12) => 
                           ID_EX_RF_OUT2_NEXT_12_port, REGOUT(11) => 
                           ID_EX_RF_OUT2_NEXT_11_port, REGOUT(10) => 
                           ID_EX_RF_OUT2_NEXT_10_port, REGOUT(9) => 
                           ID_EX_RF_OUT2_NEXT_9_port, REGOUT(8) => 
                           ID_EX_RF_OUT2_NEXT_8_port, REGOUT(7) => 
                           ID_EX_RF_OUT2_NEXT_7_port, REGOUT(6) => 
                           ID_EX_RF_OUT2_NEXT_6_port, REGOUT(5) => 
                           ID_EX_RF_OUT2_NEXT_5_port, REGOUT(4) => 
                           ID_EX_RF_OUT2_NEXT_4_port, REGOUT(3) => 
                           ID_EX_RF_OUT2_NEXT_3_port, REGOUT(2) => 
                           ID_EX_RF_OUT2_NEXT_2_port, REGOUT(1) => 
                           ID_EX_RF_OUT2_NEXT_1_port, REGOUT(0) => 
                           ID_EX_RF_OUT2_NEXT_0_port);
   LATCH_IMM : LDR_N32_2 port map( RST => net31258, EN => RegIMM_LATCH_EN, 
                           REGIN(31) => IMM_OUT_31_port, REGIN(30) => 
                           IMM_OUT_30_port, REGIN(29) => IMM_OUT_29_port, 
                           REGIN(28) => IMM_OUT_28_port, REGIN(27) => 
                           IMM_OUT_27_port, REGIN(26) => IMM_OUT_26_port, 
                           REGIN(25) => IMM_OUT_25_port, REGIN(24) => 
                           IMM_OUT_24_port, REGIN(23) => IMM_OUT_23_port, 
                           REGIN(22) => IMM_OUT_22_port, REGIN(21) => 
                           IMM_OUT_21_port, REGIN(20) => IMM_OUT_20_port, 
                           REGIN(19) => IMM_OUT_19_port, REGIN(18) => 
                           IMM_OUT_18_port, REGIN(17) => IMM_OUT_17_port, 
                           REGIN(16) => IMM_OUT_16_port, REGIN(15) => 
                           IMM_OUT_15_port, REGIN(14) => IMM_OUT_14_port, 
                           REGIN(13) => IMM_OUT_13_port, REGIN(12) => 
                           IMM_OUT_12_port, REGIN(11) => IMM_OUT_11_port, 
                           REGIN(10) => IMM_OUT_10_port, REGIN(9) => 
                           IMM_OUT_9_port, REGIN(8) => IMM_OUT_8_port, REGIN(7)
                           => IMM_OUT_7_port, REGIN(6) => IMM_OUT_6_port, 
                           REGIN(5) => IMM_OUT_5_port, REGIN(4) => 
                           IMM_OUT_4_port, REGIN(3) => IMM_OUT_3_port, REGIN(2)
                           => IMM_OUT_2_port, REGIN(1) => IMM_OUT_1_port, 
                           REGIN(0) => IMM_OUT_0_port, REGOUT(31) => 
                           ID_EX_IMM_NEXT_31_port, REGOUT(30) => 
                           ID_EX_IMM_NEXT_30_port, REGOUT(29) => 
                           ID_EX_IMM_NEXT_29_port, REGOUT(28) => 
                           ID_EX_IMM_NEXT_28_port, REGOUT(27) => 
                           ID_EX_IMM_NEXT_27_port, REGOUT(26) => 
                           ID_EX_IMM_NEXT_26_port, REGOUT(25) => 
                           ID_EX_IMM_NEXT_25_port, REGOUT(24) => 
                           ID_EX_IMM_NEXT_24_port, REGOUT(23) => 
                           ID_EX_IMM_NEXT_23_port, REGOUT(22) => 
                           ID_EX_IMM_NEXT_22_port, REGOUT(21) => 
                           ID_EX_IMM_NEXT_21_port, REGOUT(20) => 
                           ID_EX_IMM_NEXT_20_port, REGOUT(19) => 
                           ID_EX_IMM_NEXT_19_port, REGOUT(18) => 
                           ID_EX_IMM_NEXT_18_port, REGOUT(17) => 
                           ID_EX_IMM_NEXT_17_port, REGOUT(16) => 
                           ID_EX_IMM_NEXT_16_port, REGOUT(15) => 
                           ID_EX_IMM_NEXT_15_port, REGOUT(14) => 
                           ID_EX_IMM_NEXT_14_port, REGOUT(13) => 
                           ID_EX_IMM_NEXT_13_port, REGOUT(12) => 
                           ID_EX_IMM_NEXT_12_port, REGOUT(11) => 
                           ID_EX_IMM_NEXT_11_port, REGOUT(10) => 
                           ID_EX_IMM_NEXT_10_port, REGOUT(9) => 
                           ID_EX_IMM_NEXT_9_port, REGOUT(8) => 
                           ID_EX_IMM_NEXT_8_port, REGOUT(7) => 
                           ID_EX_IMM_NEXT_7_port, REGOUT(6) => 
                           ID_EX_IMM_NEXT_6_port, REGOUT(5) => 
                           ID_EX_IMM_NEXT_5_port, REGOUT(4) => 
                           ID_EX_IMM_NEXT_4_port, REGOUT(3) => 
                           ID_EX_IMM_NEXT_3_port, REGOUT(2) => 
                           ID_EX_IMM_NEXT_2_port, REGOUT(1) => 
                           ID_EX_IMM_NEXT_1_port, REGOUT(0) => 
                           ID_EX_IMM_NEXT_0_port);
   ALU_PRE_MUX1 : MUX41_N32_1 port map( A(31) => ID_EX_RF_OUT1_31_port, A(30) 
                           => ID_EX_RF_OUT1_30_port, A(29) => 
                           ID_EX_RF_OUT1_29_port, A(28) => 
                           ID_EX_RF_OUT1_28_port, A(27) => 
                           ID_EX_RF_OUT1_27_port, A(26) => 
                           ID_EX_RF_OUT1_26_port, A(25) => 
                           ID_EX_RF_OUT1_25_port, A(24) => 
                           ID_EX_RF_OUT1_24_port, A(23) => 
                           ID_EX_RF_OUT1_23_port, A(22) => 
                           ID_EX_RF_OUT1_22_port, A(21) => 
                           ID_EX_RF_OUT1_21_port, A(20) => 
                           ID_EX_RF_OUT1_20_port, A(19) => 
                           ID_EX_RF_OUT1_19_port, A(18) => 
                           ID_EX_RF_OUT1_18_port, A(17) => 
                           ID_EX_RF_OUT1_17_port, A(16) => 
                           ID_EX_RF_OUT1_16_port, A(15) => 
                           ID_EX_RF_OUT1_15_port, A(14) => 
                           ID_EX_RF_OUT1_14_port, A(13) => 
                           ID_EX_RF_OUT1_13_port, A(12) => 
                           ID_EX_RF_OUT1_12_port, A(11) => 
                           ID_EX_RF_OUT1_11_port, A(10) => 
                           ID_EX_RF_OUT1_10_port, A(9) => ID_EX_RF_OUT1_9_port,
                           A(8) => ID_EX_RF_OUT1_8_port, A(7) => 
                           ID_EX_RF_OUT1_7_port, A(6) => ID_EX_RF_OUT1_6_port, 
                           A(5) => ID_EX_RF_OUT1_5_port, A(4) => 
                           ID_EX_RF_OUT1_4_port, A(3) => ID_EX_RF_OUT1_3_port, 
                           A(2) => ID_EX_RF_OUT1_2_port, A(1) => 
                           ID_EX_RF_OUT1_1_port, A(0) => ID_EX_RF_OUT1_0_port, 
                           B(31) => ALU_OUT_31_port, B(30) => ALU_OUT_30_port, 
                           B(29) => ALU_OUT_29_port, B(28) => ALU_OUT_28_port, 
                           B(27) => ALU_OUT_27_port, B(26) => ALU_OUT_26_port, 
                           B(25) => ALU_OUT_25_port, B(24) => ALU_OUT_24_port, 
                           B(23) => ALU_OUT_23_port, B(22) => ALU_OUT_22_port, 
                           B(21) => ALU_OUT_21_port, B(20) => ALU_OUT_20_port, 
                           B(19) => ALU_OUT_19_port, B(18) => ALU_OUT_18_port, 
                           B(17) => ALU_OUT_17_port, B(16) => ALU_OUT_16_port, 
                           B(15) => ALU_OUT_15_port, B(14) => ALU_OUT_14_port, 
                           B(13) => ALU_OUT_13_port, B(12) => ALU_OUT_12_port, 
                           B(11) => ALU_OUT_11_port, B(10) => ALU_OUT_10_port, 
                           B(9) => ALU_OUT_9_port, B(8) => ALU_OUT_8_port, B(7)
                           => ALU_OUT_7_port, B(6) => ALU_OUT_6_port, B(5) => 
                           ALU_OUT_5_port, B(4) => ALU_OUT_4_port, B(3) => 
                           ALU_OUT_3_port, B(2) => ALU_OUT_2_port, B(1) => 
                           ALU_OUT_1_port, B(0) => ALU_OUT_0_port, C(31) => 
                           JAL_MUX_OUT_31_port, C(30) => JAL_MUX_OUT_30_port, 
                           C(29) => JAL_MUX_OUT_29_port, C(28) => 
                           JAL_MUX_OUT_28_port, C(27) => JAL_MUX_OUT_27_port, 
                           C(26) => JAL_MUX_OUT_26_port, C(25) => 
                           JAL_MUX_OUT_25_port, C(24) => JAL_MUX_OUT_24_port, 
                           C(23) => JAL_MUX_OUT_23_port, C(22) => 
                           JAL_MUX_OUT_22_port, C(21) => JAL_MUX_OUT_21_port, 
                           C(20) => JAL_MUX_OUT_20_port, C(19) => 
                           JAL_MUX_OUT_19_port, C(18) => JAL_MUX_OUT_18_port, 
                           C(17) => JAL_MUX_OUT_17_port, C(16) => 
                           JAL_MUX_OUT_16_port, C(15) => JAL_MUX_OUT_15_port, 
                           C(14) => JAL_MUX_OUT_14_port, C(13) => 
                           JAL_MUX_OUT_13_port, C(12) => JAL_MUX_OUT_12_port, 
                           C(11) => JAL_MUX_OUT_11_port, C(10) => 
                           JAL_MUX_OUT_10_port, C(9) => JAL_MUX_OUT_9_port, 
                           C(8) => JAL_MUX_OUT_8_port, C(7) => 
                           JAL_MUX_OUT_7_port, C(6) => JAL_MUX_OUT_6_port, C(5)
                           => JAL_MUX_OUT_5_port, C(4) => JAL_MUX_OUT_4_port, 
                           C(3) => JAL_MUX_OUT_3_port, C(2) => 
                           JAL_MUX_OUT_2_port, C(1) => JAL_MUX_OUT_1_port, C(0)
                           => JAL_MUX_OUT_0_port, D(31) => X_Logic0_port, D(30)
                           => X_Logic0_port, D(29) => X_Logic0_port, D(28) => 
                           X_Logic0_port, D(27) => X_Logic0_port, D(26) => 
                           X_Logic0_port, D(25) => X_Logic0_port, D(24) => 
                           X_Logic0_port, D(23) => X_Logic0_port, D(22) => 
                           X_Logic0_port, D(21) => X_Logic0_port, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, S(1) => FORWARD_A_1_port, S(0) => 
                           FORWARD_A_0_port, Y(31) => ALU_PREOP1_31_port, Y(30)
                           => ALU_PREOP1_30_port, Y(29) => ALU_PREOP1_29_port, 
                           Y(28) => ALU_PREOP1_28_port, Y(27) => 
                           ALU_PREOP1_27_port, Y(26) => ALU_PREOP1_26_port, 
                           Y(25) => ALU_PREOP1_25_port, Y(24) => 
                           ALU_PREOP1_24_port, Y(23) => ALU_PREOP1_23_port, 
                           Y(22) => ALU_PREOP1_22_port, Y(21) => 
                           ALU_PREOP1_21_port, Y(20) => ALU_PREOP1_20_port, 
                           Y(19) => ALU_PREOP1_19_port, Y(18) => 
                           ALU_PREOP1_18_port, Y(17) => ALU_PREOP1_17_port, 
                           Y(16) => ALU_PREOP1_16_port, Y(15) => 
                           ALU_PREOP1_15_port, Y(14) => ALU_PREOP1_14_port, 
                           Y(13) => ALU_PREOP1_13_port, Y(12) => 
                           ALU_PREOP1_12_port, Y(11) => ALU_PREOP1_11_port, 
                           Y(10) => ALU_PREOP1_10_port, Y(9) => 
                           ALU_PREOP1_9_port, Y(8) => ALU_PREOP1_8_port, Y(7) 
                           => ALU_PREOP1_7_port, Y(6) => ALU_PREOP1_6_port, 
                           Y(5) => ALU_PREOP1_5_port, Y(4) => ALU_PREOP1_4_port
                           , Y(3) => ALU_PREOP1_3_port, Y(2) => 
                           ALU_PREOP1_2_port, Y(1) => ALU_PREOP1_1_port, Y(0) 
                           => ALU_PREOP1_0_port);
   ALU_PRE_MUX2 : MUX41_N32_0 port map( A(31) => ID_EX_RF_OUT2_31_port, A(30) 
                           => ID_EX_RF_OUT2_30_port, A(29) => 
                           ID_EX_RF_OUT2_29_port, A(28) => 
                           ID_EX_RF_OUT2_28_port, A(27) => 
                           ID_EX_RF_OUT2_27_port, A(26) => 
                           ID_EX_RF_OUT2_26_port, A(25) => 
                           ID_EX_RF_OUT2_25_port, A(24) => 
                           ID_EX_RF_OUT2_24_port, A(23) => 
                           ID_EX_RF_OUT2_23_port, A(22) => 
                           ID_EX_RF_OUT2_22_port, A(21) => 
                           ID_EX_RF_OUT2_21_port, A(20) => 
                           ID_EX_RF_OUT2_20_port, A(19) => 
                           ID_EX_RF_OUT2_19_port, A(18) => 
                           ID_EX_RF_OUT2_18_port, A(17) => 
                           ID_EX_RF_OUT2_17_port, A(16) => 
                           ID_EX_RF_OUT2_16_port, A(15) => 
                           ID_EX_RF_OUT2_15_port, A(14) => 
                           ID_EX_RF_OUT2_14_port, A(13) => 
                           ID_EX_RF_OUT2_13_port, A(12) => 
                           ID_EX_RF_OUT2_12_port, A(11) => 
                           ID_EX_RF_OUT2_11_port, A(10) => 
                           ID_EX_RF_OUT2_10_port, A(9) => ID_EX_RF_OUT2_9_port,
                           A(8) => ID_EX_RF_OUT2_8_port, A(7) => 
                           ID_EX_RF_OUT2_7_port, A(6) => ID_EX_RF_OUT2_6_port, 
                           A(5) => ID_EX_RF_OUT2_5_port, A(4) => 
                           ID_EX_RF_OUT2_4_port, A(3) => ID_EX_RF_OUT2_3_port, 
                           A(2) => ID_EX_RF_OUT2_2_port, A(1) => 
                           ID_EX_RF_OUT2_1_port, A(0) => ID_EX_RF_OUT2_0_port, 
                           B(31) => ALU_OUT_31_port, B(30) => ALU_OUT_30_port, 
                           B(29) => ALU_OUT_29_port, B(28) => ALU_OUT_28_port, 
                           B(27) => ALU_OUT_27_port, B(26) => ALU_OUT_26_port, 
                           B(25) => ALU_OUT_25_port, B(24) => ALU_OUT_24_port, 
                           B(23) => ALU_OUT_23_port, B(22) => ALU_OUT_22_port, 
                           B(21) => ALU_OUT_21_port, B(20) => ALU_OUT_20_port, 
                           B(19) => ALU_OUT_19_port, B(18) => ALU_OUT_18_port, 
                           B(17) => ALU_OUT_17_port, B(16) => ALU_OUT_16_port, 
                           B(15) => ALU_OUT_15_port, B(14) => ALU_OUT_14_port, 
                           B(13) => ALU_OUT_13_port, B(12) => ALU_OUT_12_port, 
                           B(11) => ALU_OUT_11_port, B(10) => ALU_OUT_10_port, 
                           B(9) => ALU_OUT_9_port, B(8) => ALU_OUT_8_port, B(7)
                           => ALU_OUT_7_port, B(6) => ALU_OUT_6_port, B(5) => 
                           ALU_OUT_5_port, B(4) => ALU_OUT_4_port, B(3) => 
                           ALU_OUT_3_port, B(2) => ALU_OUT_2_port, B(1) => 
                           ALU_OUT_1_port, B(0) => ALU_OUT_0_port, C(31) => 
                           JAL_MUX_OUT_31_port, C(30) => JAL_MUX_OUT_30_port, 
                           C(29) => JAL_MUX_OUT_29_port, C(28) => 
                           JAL_MUX_OUT_28_port, C(27) => JAL_MUX_OUT_27_port, 
                           C(26) => JAL_MUX_OUT_26_port, C(25) => 
                           JAL_MUX_OUT_25_port, C(24) => JAL_MUX_OUT_24_port, 
                           C(23) => JAL_MUX_OUT_23_port, C(22) => 
                           JAL_MUX_OUT_22_port, C(21) => JAL_MUX_OUT_21_port, 
                           C(20) => JAL_MUX_OUT_20_port, C(19) => 
                           JAL_MUX_OUT_19_port, C(18) => JAL_MUX_OUT_18_port, 
                           C(17) => JAL_MUX_OUT_17_port, C(16) => 
                           JAL_MUX_OUT_16_port, C(15) => JAL_MUX_OUT_15_port, 
                           C(14) => JAL_MUX_OUT_14_port, C(13) => 
                           JAL_MUX_OUT_13_port, C(12) => JAL_MUX_OUT_12_port, 
                           C(11) => JAL_MUX_OUT_11_port, C(10) => 
                           JAL_MUX_OUT_10_port, C(9) => JAL_MUX_OUT_9_port, 
                           C(8) => JAL_MUX_OUT_8_port, C(7) => 
                           JAL_MUX_OUT_7_port, C(6) => JAL_MUX_OUT_6_port, C(5)
                           => JAL_MUX_OUT_5_port, C(4) => JAL_MUX_OUT_4_port, 
                           C(3) => JAL_MUX_OUT_3_port, C(2) => 
                           JAL_MUX_OUT_2_port, C(1) => JAL_MUX_OUT_1_port, C(0)
                           => JAL_MUX_OUT_0_port, D(31) => X_Logic0_port, D(30)
                           => X_Logic0_port, D(29) => X_Logic0_port, D(28) => 
                           X_Logic0_port, D(27) => X_Logic0_port, D(26) => 
                           X_Logic0_port, D(25) => X_Logic0_port, D(24) => 
                           X_Logic0_port, D(23) => X_Logic0_port, D(22) => 
                           X_Logic0_port, D(21) => X_Logic0_port, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, S(1) => FORWARD_B_1_port, S(0) => 
                           FORWARD_B_0_port, Y(31) => ALU_PREOP2_31_port, Y(30)
                           => ALU_PREOP2_30_port, Y(29) => ALU_PREOP2_29_port, 
                           Y(28) => ALU_PREOP2_28_port, Y(27) => 
                           ALU_PREOP2_27_port, Y(26) => ALU_PREOP2_26_port, 
                           Y(25) => ALU_PREOP2_25_port, Y(24) => 
                           ALU_PREOP2_24_port, Y(23) => ALU_PREOP2_23_port, 
                           Y(22) => ALU_PREOP2_22_port, Y(21) => 
                           ALU_PREOP2_21_port, Y(20) => ALU_PREOP2_20_port, 
                           Y(19) => ALU_PREOP2_19_port, Y(18) => 
                           ALU_PREOP2_18_port, Y(17) => ALU_PREOP2_17_port, 
                           Y(16) => ALU_PREOP2_16_port, Y(15) => 
                           ALU_PREOP2_15_port, Y(14) => ALU_PREOP2_14_port, 
                           Y(13) => ALU_PREOP2_13_port, Y(12) => 
                           ALU_PREOP2_12_port, Y(11) => ALU_PREOP2_11_port, 
                           Y(10) => ALU_PREOP2_10_port, Y(9) => 
                           ALU_PREOP2_9_port, Y(8) => ALU_PREOP2_8_port, Y(7) 
                           => ALU_PREOP2_7_port, Y(6) => ALU_PREOP2_6_port, 
                           Y(5) => ALU_PREOP2_5_port, Y(4) => ALU_PREOP2_4_port
                           , Y(3) => ALU_PREOP2_3_port, Y(2) => 
                           ALU_PREOP2_2_port, Y(1) => ALU_PREOP2_1_port, Y(0) 
                           => ALU_PREOP2_0_port);
   ALU_MUX1 : MUX21_N32_3 port map( A(31) => ALU_PREOP1_31_port, A(30) => 
                           ALU_PREOP1_30_port, A(29) => ALU_PREOP1_29_port, 
                           A(28) => ALU_PREOP1_28_port, A(27) => 
                           ALU_PREOP1_27_port, A(26) => ALU_PREOP1_26_port, 
                           A(25) => ALU_PREOP1_25_port, A(24) => 
                           ALU_PREOP1_24_port, A(23) => ALU_PREOP1_23_port, 
                           A(22) => ALU_PREOP1_22_port, A(21) => 
                           ALU_PREOP1_21_port, A(20) => ALU_PREOP1_20_port, 
                           A(19) => ALU_PREOP1_19_port, A(18) => 
                           ALU_PREOP1_18_port, A(17) => ALU_PREOP1_17_port, 
                           A(16) => ALU_PREOP1_16_port, A(15) => 
                           ALU_PREOP1_15_port, A(14) => ALU_PREOP1_14_port, 
                           A(13) => ALU_PREOP1_13_port, A(12) => 
                           ALU_PREOP1_12_port, A(11) => ALU_PREOP1_11_port, 
                           A(10) => ALU_PREOP1_10_port, A(9) => 
                           ALU_PREOP1_9_port, A(8) => ALU_PREOP1_8_port, A(7) 
                           => ALU_PREOP1_7_port, A(6) => ALU_PREOP1_6_port, 
                           A(5) => ALU_PREOP1_5_port, A(4) => ALU_PREOP1_4_port
                           , A(3) => ALU_PREOP1_3_port, A(2) => 
                           ALU_PREOP1_2_port, A(1) => ALU_PREOP1_1_port, A(0) 
                           => ALU_PREOP1_0_port, B(31) => ID_EX_NPC_31_port, 
                           B(30) => ID_EX_NPC_30_port, B(29) => 
                           ID_EX_NPC_29_port, B(28) => ID_EX_NPC_28_port, B(27)
                           => ID_EX_NPC_27_port, B(26) => ID_EX_NPC_26_port, 
                           B(25) => ID_EX_NPC_25_port, B(24) => 
                           ID_EX_NPC_24_port, B(23) => ID_EX_NPC_23_port, B(22)
                           => ID_EX_NPC_22_port, B(21) => ID_EX_NPC_21_port, 
                           B(20) => ID_EX_NPC_20_port, B(19) => 
                           ID_EX_NPC_19_port, B(18) => ID_EX_NPC_18_port, B(17)
                           => ID_EX_NPC_17_port, B(16) => ID_EX_NPC_16_port, 
                           B(15) => ID_EX_NPC_15_port, B(14) => 
                           ID_EX_NPC_14_port, B(13) => ID_EX_NPC_13_port, B(12)
                           => ID_EX_NPC_12_port, B(11) => ID_EX_NPC_11_port, 
                           B(10) => ID_EX_NPC_10_port, B(9) => ID_EX_NPC_9_port
                           , B(8) => ID_EX_NPC_8_port, B(7) => ID_EX_NPC_7_port
                           , B(6) => ID_EX_NPC_6_port, B(5) => ID_EX_NPC_5_port
                           , B(4) => ID_EX_NPC_4_port, B(3) => ID_EX_NPC_3_port
                           , B(2) => ID_EX_NPC_2_port, B(1) => ID_EX_NPC_1_port
                           , B(0) => ID_EX_NPC_0_port, S => MUXA_SEL, Y(31) => 
                           ALU_OP1_31_port, Y(30) => ALU_OP1_30_port, Y(29) => 
                           ALU_OP1_29_port, Y(28) => ALU_OP1_28_port, Y(27) => 
                           ALU_OP1_27_port, Y(26) => ALU_OP1_26_port, Y(25) => 
                           ALU_OP1_25_port, Y(24) => ALU_OP1_24_port, Y(23) => 
                           ALU_OP1_23_port, Y(22) => ALU_OP1_22_port, Y(21) => 
                           ALU_OP1_21_port, Y(20) => ALU_OP1_20_port, Y(19) => 
                           ALU_OP1_19_port, Y(18) => ALU_OP1_18_port, Y(17) => 
                           ALU_OP1_17_port, Y(16) => ALU_OP1_16_port, Y(15) => 
                           ALU_OP1_15_port, Y(14) => ALU_OP1_14_port, Y(13) => 
                           ALU_OP1_13_port, Y(12) => ALU_OP1_12_port, Y(11) => 
                           ALU_OP1_11_port, Y(10) => ALU_OP1_10_port, Y(9) => 
                           ALU_OP1_9_port, Y(8) => ALU_OP1_8_port, Y(7) => 
                           ALU_OP1_7_port, Y(6) => ALU_OP1_6_port, Y(5) => 
                           ALU_OP1_5_port, Y(4) => ALU_OP1_4_port, Y(3) => 
                           ALU_OP1_3_port, Y(2) => ALU_OP1_2_port, Y(1) => 
                           ALU_OP1_1_port, Y(0) => ALU_OP1_0_port);
   ALU_MUX2 : MUX21_N32_2 port map( A(31) => ALU_PREOP2_31_port, A(30) => 
                           ALU_PREOP2_30_port, A(29) => ALU_PREOP2_29_port, 
                           A(28) => ALU_PREOP2_28_port, A(27) => 
                           ALU_PREOP2_27_port, A(26) => ALU_PREOP2_26_port, 
                           A(25) => ALU_PREOP2_25_port, A(24) => 
                           ALU_PREOP2_24_port, A(23) => ALU_PREOP2_23_port, 
                           A(22) => ALU_PREOP2_22_port, A(21) => 
                           ALU_PREOP2_21_port, A(20) => ALU_PREOP2_20_port, 
                           A(19) => ALU_PREOP2_19_port, A(18) => 
                           ALU_PREOP2_18_port, A(17) => ALU_PREOP2_17_port, 
                           A(16) => ALU_PREOP2_16_port, A(15) => 
                           ALU_PREOP2_15_port, A(14) => ALU_PREOP2_14_port, 
                           A(13) => ALU_PREOP2_13_port, A(12) => 
                           ALU_PREOP2_12_port, A(11) => ALU_PREOP2_11_port, 
                           A(10) => ALU_PREOP2_10_port, A(9) => 
                           ALU_PREOP2_9_port, A(8) => ALU_PREOP2_8_port, A(7) 
                           => ALU_PREOP2_7_port, A(6) => ALU_PREOP2_6_port, 
                           A(5) => ALU_PREOP2_5_port, A(4) => ALU_PREOP2_4_port
                           , A(3) => ALU_PREOP2_3_port, A(2) => 
                           ALU_PREOP2_2_port, A(1) => ALU_PREOP2_1_port, A(0) 
                           => ALU_PREOP2_0_port, B(31) => ID_EX_IMM_31_port, 
                           B(30) => ID_EX_IMM_30_port, B(29) => 
                           ID_EX_IMM_29_port, B(28) => ID_EX_IMM_28_port, B(27)
                           => ID_EX_IMM_27_port, B(26) => ID_EX_IMM_26_port, 
                           B(25) => ID_EX_IMM_25_port, B(24) => 
                           ID_EX_IMM_24_port, B(23) => ID_EX_IMM_23_port, B(22)
                           => ID_EX_IMM_22_port, B(21) => ID_EX_IMM_21_port, 
                           B(20) => ID_EX_IMM_20_port, B(19) => 
                           ID_EX_IMM_19_port, B(18) => ID_EX_IMM_18_port, B(17)
                           => ID_EX_IMM_17_port, B(16) => ID_EX_IMM_16_port, 
                           B(15) => ID_EX_IMM_15_port, B(14) => 
                           ID_EX_IMM_14_port, B(13) => ID_EX_IMM_13_port, B(12)
                           => ID_EX_IMM_12_port, B(11) => ID_EX_IMM_11_port, 
                           B(10) => ID_EX_IMM_10_port, B(9) => ID_EX_IMM_9_port
                           , B(8) => ID_EX_IMM_8_port, B(7) => ID_EX_IMM_7_port
                           , B(6) => ID_EX_IMM_6_port, B(5) => ID_EX_IMM_5_port
                           , B(4) => ID_EX_IMM_4_port, B(3) => ID_EX_IMM_3_port
                           , B(2) => ID_EX_IMM_2_port, B(1) => ID_EX_IMM_1_port
                           , B(0) => ID_EX_IMM_0_port, S => MUXB_SEL, Y(31) => 
                           ALU_OP2_31_port, Y(30) => ALU_OP2_30_port, Y(29) => 
                           ALU_OP2_29_port, Y(28) => ALU_OP2_28_port, Y(27) => 
                           ALU_OP2_27_port, Y(26) => ALU_OP2_26_port, Y(25) => 
                           ALU_OP2_25_port, Y(24) => ALU_OP2_24_port, Y(23) => 
                           ALU_OP2_23_port, Y(22) => ALU_OP2_22_port, Y(21) => 
                           ALU_OP2_21_port, Y(20) => ALU_OP2_20_port, Y(19) => 
                           ALU_OP2_19_port, Y(18) => ALU_OP2_18_port, Y(17) => 
                           ALU_OP2_17_port, Y(16) => ALU_OP2_16_port, Y(15) => 
                           ALU_OP2_15_port, Y(14) => ALU_OP2_14_port, Y(13) => 
                           ALU_OP2_13_port, Y(12) => ALU_OP2_12_port, Y(11) => 
                           ALU_OP2_11_port, Y(10) => ALU_OP2_10_port, Y(9) => 
                           ALU_OP2_9_port, Y(8) => ALU_OP2_8_port, Y(7) => 
                           ALU_OP2_7_port, Y(6) => ALU_OP2_6_port, Y(5) => 
                           ALU_OP2_5_port, Y(4) => ALU_OP2_4_port, Y(3) => 
                           ALU_OP2_3_port, Y(2) => ALU_OP2_2_port, Y(1) => 
                           ALU_OP2_1_port, Y(0) => ALU_OP2_0_port);
   ARITHMETIC_LOGIC_UNIT : ALU_N32_NB8 port map( OP1(31) => ALU_OP1_31_port, 
                           OP1(30) => ALU_OP1_30_port, OP1(29) => 
                           ALU_OP1_29_port, OP1(28) => ALU_OP1_28_port, OP1(27)
                           => ALU_OP1_27_port, OP1(26) => ALU_OP1_26_port, 
                           OP1(25) => ALU_OP1_25_port, OP1(24) => 
                           ALU_OP1_24_port, OP1(23) => ALU_OP1_23_port, OP1(22)
                           => ALU_OP1_22_port, OP1(21) => ALU_OP1_21_port, 
                           OP1(20) => ALU_OP1_20_port, OP1(19) => 
                           ALU_OP1_19_port, OP1(18) => ALU_OP1_18_port, OP1(17)
                           => ALU_OP1_17_port, OP1(16) => ALU_OP1_16_port, 
                           OP1(15) => ALU_OP1_15_port, OP1(14) => 
                           ALU_OP1_14_port, OP1(13) => ALU_OP1_13_port, OP1(12)
                           => ALU_OP1_12_port, OP1(11) => ALU_OP1_11_port, 
                           OP1(10) => ALU_OP1_10_port, OP1(9) => ALU_OP1_9_port
                           , OP1(8) => ALU_OP1_8_port, OP1(7) => ALU_OP1_7_port
                           , OP1(6) => ALU_OP1_6_port, OP1(5) => ALU_OP1_5_port
                           , OP1(4) => ALU_OP1_4_port, OP1(3) => ALU_OP1_3_port
                           , OP1(2) => ALU_OP1_2_port, OP1(1) => ALU_OP1_1_port
                           , OP1(0) => ALU_OP1_0_port, OP2(31) => 
                           ALU_OP2_31_port, OP2(30) => ALU_OP2_30_port, OP2(29)
                           => ALU_OP2_29_port, OP2(28) => ALU_OP2_28_port, 
                           OP2(27) => ALU_OP2_27_port, OP2(26) => 
                           ALU_OP2_26_port, OP2(25) => ALU_OP2_25_port, OP2(24)
                           => ALU_OP2_24_port, OP2(23) => ALU_OP2_23_port, 
                           OP2(22) => ALU_OP2_22_port, OP2(21) => 
                           ALU_OP2_21_port, OP2(20) => ALU_OP2_20_port, OP2(19)
                           => ALU_OP2_19_port, OP2(18) => ALU_OP2_18_port, 
                           OP2(17) => ALU_OP2_17_port, OP2(16) => 
                           ALU_OP2_16_port, OP2(15) => ALU_OP2_15_port, OP2(14)
                           => ALU_OP2_14_port, OP2(13) => ALU_OP2_13_port, 
                           OP2(12) => ALU_OP2_12_port, OP2(11) => 
                           ALU_OP2_11_port, OP2(10) => ALU_OP2_10_port, OP2(9) 
                           => ALU_OP2_9_port, OP2(8) => ALU_OP2_8_port, OP2(7) 
                           => ALU_OP2_7_port, OP2(6) => ALU_OP2_6_port, OP2(5) 
                           => ALU_OP2_5_port, OP2(4) => ALU_OP2_4_port, OP2(3) 
                           => ALU_OP2_3_port, OP2(2) => ALU_OP2_2_port, OP2(1) 
                           => ALU_OP2_1_port, OP2(0) => ALU_OP2_0_port, OPC(0) 
                           => ALU_OPCODE(0), OPC(1) => ALU_OPCODE(1), OPC(2) =>
                           ALU_OPCODE(2), OPC(3) => ALU_OPCODE(3), OPC(4) => 
                           ALU_OPCODE(4), OPC(5) => ALU_OPCODE(5), OPC(6) => 
                           ALU_OPCODE(6), Y(31) => ALU_OUTPUT_31_port, Y(30) =>
                           ALU_OUTPUT_30_port, Y(29) => ALU_OUTPUT_29_port, 
                           Y(28) => ALU_OUTPUT_28_port, Y(27) => 
                           ALU_OUTPUT_27_port, Y(26) => ALU_OUTPUT_26_port, 
                           Y(25) => ALU_OUTPUT_25_port, Y(24) => 
                           ALU_OUTPUT_24_port, Y(23) => ALU_OUTPUT_23_port, 
                           Y(22) => ALU_OUTPUT_22_port, Y(21) => 
                           ALU_OUTPUT_21_port, Y(20) => ALU_OUTPUT_20_port, 
                           Y(19) => ALU_OUTPUT_19_port, Y(18) => 
                           ALU_OUTPUT_18_port, Y(17) => ALU_OUTPUT_17_port, 
                           Y(16) => ALU_OUTPUT_16_port, Y(15) => 
                           ALU_OUTPUT_15_port, Y(14) => ALU_OUTPUT_14_port, 
                           Y(13) => ALU_OUTPUT_13_port, Y(12) => 
                           ALU_OUTPUT_12_port, Y(11) => ALU_OUTPUT_11_port, 
                           Y(10) => ALU_OUTPUT_10_port, Y(9) => 
                           ALU_OUTPUT_9_port, Y(8) => ALU_OUTPUT_8_port, Y(7) 
                           => ALU_OUTPUT_7_port, Y(6) => ALU_OUTPUT_6_port, 
                           Y(5) => ALU_OUTPUT_5_port, Y(4) => ALU_OUTPUT_4_port
                           , Y(3) => ALU_OUTPUT_3_port, Y(2) => 
                           ALU_OUTPUT_2_port, Y(1) => ALU_OUTPUT_1_port, Y(0) 
                           => ALU_OUTPUT_0_port, Z => n_1704);
   BRANCH_MUX : MUX21_L_320 port map( A => ZERO_OUT, B => n18_port, S => 
                           EQ_COND, Y => BRANCH_DETECT);
   Z_DETECTOR : ZERO_DETECTOR_N32_1 port map( A(31) => ALU_PREOP1_31_port, 
                           A(30) => ALU_PREOP1_30_port, A(29) => 
                           ALU_PREOP1_29_port, A(28) => ALU_PREOP1_28_port, 
                           A(27) => ALU_PREOP1_27_port, A(26) => 
                           ALU_PREOP1_26_port, A(25) => ALU_PREOP1_25_port, 
                           A(24) => ALU_PREOP1_24_port, A(23) => 
                           ALU_PREOP1_23_port, A(22) => ALU_PREOP1_22_port, 
                           A(21) => ALU_PREOP1_21_port, A(20) => 
                           ALU_PREOP1_20_port, A(19) => ALU_PREOP1_19_port, 
                           A(18) => ALU_PREOP1_18_port, A(17) => 
                           ALU_PREOP1_17_port, A(16) => ALU_PREOP1_16_port, 
                           A(15) => ALU_PREOP1_15_port, A(14) => 
                           ALU_PREOP1_14_port, A(13) => ALU_PREOP1_13_port, 
                           A(12) => ALU_PREOP1_12_port, A(11) => 
                           ALU_PREOP1_11_port, A(10) => ALU_PREOP1_10_port, 
                           A(9) => ALU_PREOP1_9_port, A(8) => ALU_PREOP1_8_port
                           , A(7) => ALU_PREOP1_7_port, A(6) => 
                           ALU_PREOP1_6_port, A(5) => ALU_PREOP1_5_port, A(4) 
                           => ALU_PREOP1_4_port, A(3) => ALU_PREOP1_3_port, 
                           A(2) => ALU_PREOP1_2_port, A(1) => ALU_PREOP1_1_port
                           , A(0) => ALU_PREOP1_0_port, Y => ZERO_OUT);
   FORWARDING_UNIT : FU_N5 port map( RS1(4) => ID_EX_RS1_4_port, RS1(3) => 
                           ID_EX_RS1_3_port, RS1(2) => ID_EX_RS1_2_port, RS1(1)
                           => ID_EX_RS1_1_port, RS1(0) => ID_EX_RS1_0_port, 
                           RS2(4) => ID_EX_RS2_4_port, RS2(3) => 
                           ID_EX_RS2_3_port, RS2(2) => ID_EX_RS2_2_port, RS2(1)
                           => ID_EX_RS2_1_port, RS2(0) => ID_EX_RS2_0_port, 
                           RD_MEM(4) => EX_MEM_RD_4_port, RD_MEM(3) => 
                           EX_MEM_RD_3_port, RD_MEM(2) => EX_MEM_RD_2_port, 
                           RD_MEM(1) => EX_MEM_RD_1_port, RD_MEM(0) => 
                           EX_MEM_RD_0_port, RD_WB(4) => MEM_WB_RD_4_port, 
                           RD_WB(3) => MEM_WB_RD_3_port, RD_WB(2) => 
                           MEM_WB_RD_2_port, RD_WB(1) => MEM_WB_RD_1_port, 
                           RD_WB(0) => MEM_WB_RD_0_port, RF_WE_MEM => 
                           EX_MEM_RF_WE, RF_WE_WB => MEM_WB_RF_WE, FORWARD_A(1)
                           => FORWARD_A_1_port, FORWARD_A(0) => 
                           FORWARD_A_0_port, FORWARD_B(1) => FORWARD_B_1_port, 
                           FORWARD_B(0) => FORWARD_B_0_port);
   LATCH_ALUOUT : LDR_N32_1 port map( RST => net31258, EN => ALU_OUTREG_EN, 
                           REGIN(31) => ALU_OUTPUT_31_port, REGIN(30) => 
                           ALU_OUTPUT_30_port, REGIN(29) => ALU_OUTPUT_29_port,
                           REGIN(28) => ALU_OUTPUT_28_port, REGIN(27) => 
                           ALU_OUTPUT_27_port, REGIN(26) => ALU_OUTPUT_26_port,
                           REGIN(25) => ALU_OUTPUT_25_port, REGIN(24) => 
                           ALU_OUTPUT_24_port, REGIN(23) => ALU_OUTPUT_23_port,
                           REGIN(22) => ALU_OUTPUT_22_port, REGIN(21) => 
                           ALU_OUTPUT_21_port, REGIN(20) => ALU_OUTPUT_20_port,
                           REGIN(19) => ALU_OUTPUT_19_port, REGIN(18) => 
                           ALU_OUTPUT_18_port, REGIN(17) => ALU_OUTPUT_17_port,
                           REGIN(16) => ALU_OUTPUT_16_port, REGIN(15) => 
                           ALU_OUTPUT_15_port, REGIN(14) => ALU_OUTPUT_14_port,
                           REGIN(13) => ALU_OUTPUT_13_port, REGIN(12) => 
                           ALU_OUTPUT_12_port, REGIN(11) => ALU_OUTPUT_11_port,
                           REGIN(10) => ALU_OUTPUT_10_port, REGIN(9) => 
                           ALU_OUTPUT_9_port, REGIN(8) => ALU_OUTPUT_8_port, 
                           REGIN(7) => ALU_OUTPUT_7_port, REGIN(6) => 
                           ALU_OUTPUT_6_port, REGIN(5) => ALU_OUTPUT_5_port, 
                           REGIN(4) => ALU_OUTPUT_4_port, REGIN(3) => 
                           ALU_OUTPUT_3_port, REGIN(2) => ALU_OUTPUT_2_port, 
                           REGIN(1) => ALU_OUTPUT_1_port, REGIN(0) => 
                           ALU_OUTPUT_0_port, REGOUT(31) => 
                           EX_MEM_ALU_OUTPUT_NEXT_31_port, REGOUT(30) => 
                           EX_MEM_ALU_OUTPUT_NEXT_30_port, REGOUT(29) => 
                           EX_MEM_ALU_OUTPUT_NEXT_29_port, REGOUT(28) => 
                           EX_MEM_ALU_OUTPUT_NEXT_28_port, REGOUT(27) => 
                           EX_MEM_ALU_OUTPUT_NEXT_27_port, REGOUT(26) => 
                           EX_MEM_ALU_OUTPUT_NEXT_26_port, REGOUT(25) => 
                           EX_MEM_ALU_OUTPUT_NEXT_25_port, REGOUT(24) => 
                           EX_MEM_ALU_OUTPUT_NEXT_24_port, REGOUT(23) => 
                           EX_MEM_ALU_OUTPUT_NEXT_23_port, REGOUT(22) => 
                           EX_MEM_ALU_OUTPUT_NEXT_22_port, REGOUT(21) => 
                           EX_MEM_ALU_OUTPUT_NEXT_21_port, REGOUT(20) => 
                           EX_MEM_ALU_OUTPUT_NEXT_20_port, REGOUT(19) => 
                           EX_MEM_ALU_OUTPUT_NEXT_19_port, REGOUT(18) => 
                           EX_MEM_ALU_OUTPUT_NEXT_18_port, REGOUT(17) => 
                           EX_MEM_ALU_OUTPUT_NEXT_17_port, REGOUT(16) => 
                           EX_MEM_ALU_OUTPUT_NEXT_16_port, REGOUT(15) => 
                           EX_MEM_ALU_OUTPUT_NEXT_15_port, REGOUT(14) => 
                           EX_MEM_ALU_OUTPUT_NEXT_14_port, REGOUT(13) => 
                           EX_MEM_ALU_OUTPUT_NEXT_13_port, REGOUT(12) => 
                           EX_MEM_ALU_OUTPUT_NEXT_12_port, REGOUT(11) => 
                           EX_MEM_ALU_OUTPUT_NEXT_11_port, REGOUT(10) => 
                           EX_MEM_ALU_OUTPUT_NEXT_10_port, REGOUT(9) => 
                           EX_MEM_ALU_OUTPUT_NEXT_9_port, REGOUT(8) => 
                           EX_MEM_ALU_OUTPUT_NEXT_8_port, REGOUT(7) => 
                           EX_MEM_ALU_OUTPUT_NEXT_7_port, REGOUT(6) => 
                           EX_MEM_ALU_OUTPUT_NEXT_6_port, REGOUT(5) => 
                           EX_MEM_ALU_OUTPUT_NEXT_5_port, REGOUT(4) => 
                           EX_MEM_ALU_OUTPUT_NEXT_4_port, REGOUT(3) => 
                           EX_MEM_ALU_OUTPUT_NEXT_3_port, REGOUT(2) => 
                           EX_MEM_ALU_OUTPUT_NEXT_2_port, REGOUT(1) => 
                           EX_MEM_ALU_OUTPUT_NEXT_1_port, REGOUT(0) => 
                           EX_MEM_ALU_OUTPUT_NEXT_0_port);
   LATCH_BRANCH : LD_224 port map( RST => net31258, EN => ALU_OUTREG_EN, D => 
                           BRANCH_DETECT, Q => EX_MEM_BRANCH_DETECT_NEXT);
   LATCH_LMD : LDR_N32_0 port map( RST => net31258, EN => LMD_LATCH_EN, 
                           REGIN(31) => DRAM_OUT(31), REGIN(30) => DRAM_OUT(30)
                           , REGIN(29) => DRAM_OUT(29), REGIN(28) => 
                           DRAM_OUT(28), REGIN(27) => DRAM_OUT(27), REGIN(26) 
                           => DRAM_OUT(26), REGIN(25) => DRAM_OUT(25), 
                           REGIN(24) => DRAM_OUT(24), REGIN(23) => DRAM_OUT(23)
                           , REGIN(22) => DRAM_OUT(22), REGIN(21) => 
                           DRAM_OUT(21), REGIN(20) => DRAM_OUT(20), REGIN(19) 
                           => DRAM_OUT(19), REGIN(18) => DRAM_OUT(18), 
                           REGIN(17) => DRAM_OUT(17), REGIN(16) => DRAM_OUT(16)
                           , REGIN(15) => DRAM_OUT(15), REGIN(14) => 
                           DRAM_OUT(14), REGIN(13) => DRAM_OUT(13), REGIN(12) 
                           => DRAM_OUT(12), REGIN(11) => DRAM_OUT(11), 
                           REGIN(10) => DRAM_OUT(10), REGIN(9) => DRAM_OUT(9), 
                           REGIN(8) => DRAM_OUT(8), REGIN(7) => DRAM_OUT(7), 
                           REGIN(6) => DRAM_OUT(6), REGIN(5) => DRAM_OUT(5), 
                           REGIN(4) => DRAM_OUT(4), REGIN(3) => DRAM_OUT(3), 
                           REGIN(2) => DRAM_OUT(2), REGIN(1) => DRAM_OUT(1), 
                           REGIN(0) => DRAM_OUT(0), REGOUT(31) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_31_port, REGOUT(30) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_30_port, REGOUT(29) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_29_port, REGOUT(28) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_28_port, REGOUT(27) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_27_port, REGOUT(26) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_26_port, REGOUT(25) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_25_port, REGOUT(24) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_24_port, REGOUT(23) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_23_port, REGOUT(22) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_22_port, REGOUT(21) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_21_port, REGOUT(20) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_20_port, REGOUT(19) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_19_port, REGOUT(18) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_18_port, REGOUT(17) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_17_port, REGOUT(16) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_16_port, REGOUT(15) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_15_port, REGOUT(14) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_14_port, REGOUT(13) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_13_port, REGOUT(12) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_12_port, REGOUT(11) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_11_port, REGOUT(10) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_10_port, REGOUT(9) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_9_port, REGOUT(8) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_8_port, REGOUT(7) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_7_port, REGOUT(6) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_6_port, REGOUT(5) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_5_port, REGOUT(4) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_4_port, REGOUT(3) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_3_port, REGOUT(2) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_2_port, REGOUT(1) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_1_port, REGOUT(0) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_0_port);
   WB_MUX : MUX21_N32_1 port map( A(31) => MEM_WB_DRAM_OUTPUT_31_port, A(30) =>
                           MEM_WB_DRAM_OUTPUT_30_port, A(29) => 
                           MEM_WB_DRAM_OUTPUT_29_port, A(28) => 
                           MEM_WB_DRAM_OUTPUT_28_port, A(27) => 
                           MEM_WB_DRAM_OUTPUT_27_port, A(26) => 
                           MEM_WB_DRAM_OUTPUT_26_port, A(25) => 
                           MEM_WB_DRAM_OUTPUT_25_port, A(24) => 
                           MEM_WB_DRAM_OUTPUT_24_port, A(23) => 
                           MEM_WB_DRAM_OUTPUT_23_port, A(22) => 
                           MEM_WB_DRAM_OUTPUT_22_port, A(21) => 
                           MEM_WB_DRAM_OUTPUT_21_port, A(20) => 
                           MEM_WB_DRAM_OUTPUT_20_port, A(19) => 
                           MEM_WB_DRAM_OUTPUT_19_port, A(18) => 
                           MEM_WB_DRAM_OUTPUT_18_port, A(17) => 
                           MEM_WB_DRAM_OUTPUT_17_port, A(16) => 
                           MEM_WB_DRAM_OUTPUT_16_port, A(15) => 
                           MEM_WB_DRAM_OUTPUT_15_port, A(14) => 
                           MEM_WB_DRAM_OUTPUT_14_port, A(13) => 
                           MEM_WB_DRAM_OUTPUT_13_port, A(12) => 
                           MEM_WB_DRAM_OUTPUT_12_port, A(11) => 
                           MEM_WB_DRAM_OUTPUT_11_port, A(10) => 
                           MEM_WB_DRAM_OUTPUT_10_port, A(9) => 
                           MEM_WB_DRAM_OUTPUT_9_port, A(8) => 
                           MEM_WB_DRAM_OUTPUT_8_port, A(7) => 
                           MEM_WB_DRAM_OUTPUT_7_port, A(6) => 
                           MEM_WB_DRAM_OUTPUT_6_port, A(5) => 
                           MEM_WB_DRAM_OUTPUT_5_port, A(4) => 
                           MEM_WB_DRAM_OUTPUT_4_port, A(3) => 
                           MEM_WB_DRAM_OUTPUT_3_port, A(2) => 
                           MEM_WB_DRAM_OUTPUT_2_port, A(1) => 
                           MEM_WB_DRAM_OUTPUT_1_port, A(0) => 
                           MEM_WB_DRAM_OUTPUT_0_port, B(31) => 
                           MEM_WB_ALU_OUTPUT_31_port, B(30) => 
                           MEM_WB_ALU_OUTPUT_30_port, B(29) => 
                           MEM_WB_ALU_OUTPUT_29_port, B(28) => 
                           MEM_WB_ALU_OUTPUT_28_port, B(27) => 
                           MEM_WB_ALU_OUTPUT_27_port, B(26) => 
                           MEM_WB_ALU_OUTPUT_26_port, B(25) => 
                           MEM_WB_ALU_OUTPUT_25_port, B(24) => 
                           MEM_WB_ALU_OUTPUT_24_port, B(23) => 
                           MEM_WB_ALU_OUTPUT_23_port, B(22) => 
                           MEM_WB_ALU_OUTPUT_22_port, B(21) => 
                           MEM_WB_ALU_OUTPUT_21_port, B(20) => 
                           MEM_WB_ALU_OUTPUT_20_port, B(19) => 
                           MEM_WB_ALU_OUTPUT_19_port, B(18) => 
                           MEM_WB_ALU_OUTPUT_18_port, B(17) => 
                           MEM_WB_ALU_OUTPUT_17_port, B(16) => 
                           MEM_WB_ALU_OUTPUT_16_port, B(15) => 
                           MEM_WB_ALU_OUTPUT_15_port, B(14) => 
                           MEM_WB_ALU_OUTPUT_14_port, B(13) => 
                           MEM_WB_ALU_OUTPUT_13_port, B(12) => 
                           MEM_WB_ALU_OUTPUT_12_port, B(11) => 
                           MEM_WB_ALU_OUTPUT_11_port, B(10) => 
                           MEM_WB_ALU_OUTPUT_10_port, B(9) => 
                           MEM_WB_ALU_OUTPUT_9_port, B(8) => 
                           MEM_WB_ALU_OUTPUT_8_port, B(7) => 
                           MEM_WB_ALU_OUTPUT_7_port, B(6) => 
                           MEM_WB_ALU_OUTPUT_6_port, B(5) => 
                           MEM_WB_ALU_OUTPUT_5_port, B(4) => 
                           MEM_WB_ALU_OUTPUT_4_port, B(3) => 
                           MEM_WB_ALU_OUTPUT_3_port, B(2) => 
                           MEM_WB_ALU_OUTPUT_2_port, B(1) => 
                           MEM_WB_ALU_OUTPUT_1_port, B(0) => 
                           MEM_WB_ALU_OUTPUT_0_port, S => WB_MUX_SEL, Y(31) => 
                           WB_MUX_OUT_31_port, Y(30) => WB_MUX_OUT_30_port, 
                           Y(29) => WB_MUX_OUT_29_port, Y(28) => 
                           WB_MUX_OUT_28_port, Y(27) => WB_MUX_OUT_27_port, 
                           Y(26) => WB_MUX_OUT_26_port, Y(25) => 
                           WB_MUX_OUT_25_port, Y(24) => WB_MUX_OUT_24_port, 
                           Y(23) => WB_MUX_OUT_23_port, Y(22) => 
                           WB_MUX_OUT_22_port, Y(21) => WB_MUX_OUT_21_port, 
                           Y(20) => WB_MUX_OUT_20_port, Y(19) => 
                           WB_MUX_OUT_19_port, Y(18) => WB_MUX_OUT_18_port, 
                           Y(17) => WB_MUX_OUT_17_port, Y(16) => 
                           WB_MUX_OUT_16_port, Y(15) => WB_MUX_OUT_15_port, 
                           Y(14) => WB_MUX_OUT_14_port, Y(13) => 
                           WB_MUX_OUT_13_port, Y(12) => WB_MUX_OUT_12_port, 
                           Y(11) => WB_MUX_OUT_11_port, Y(10) => 
                           WB_MUX_OUT_10_port, Y(9) => WB_MUX_OUT_9_port, Y(8) 
                           => WB_MUX_OUT_8_port, Y(7) => WB_MUX_OUT_7_port, 
                           Y(6) => WB_MUX_OUT_6_port, Y(5) => WB_MUX_OUT_5_port
                           , Y(4) => WB_MUX_OUT_4_port, Y(3) => 
                           WB_MUX_OUT_3_port, Y(2) => WB_MUX_OUT_2_port, Y(1) 
                           => WB_MUX_OUT_1_port, Y(0) => WB_MUX_OUT_0_port);
   JAL_MUX : MUX21_N32_0 port map( A(31) => WB_MUX_OUT_31_port, A(30) => 
                           WB_MUX_OUT_30_port, A(29) => WB_MUX_OUT_29_port, 
                           A(28) => WB_MUX_OUT_28_port, A(27) => 
                           WB_MUX_OUT_27_port, A(26) => WB_MUX_OUT_26_port, 
                           A(25) => WB_MUX_OUT_25_port, A(24) => 
                           WB_MUX_OUT_24_port, A(23) => WB_MUX_OUT_23_port, 
                           A(22) => WB_MUX_OUT_22_port, A(21) => 
                           WB_MUX_OUT_21_port, A(20) => WB_MUX_OUT_20_port, 
                           A(19) => WB_MUX_OUT_19_port, A(18) => 
                           WB_MUX_OUT_18_port, A(17) => WB_MUX_OUT_17_port, 
                           A(16) => WB_MUX_OUT_16_port, A(15) => 
                           WB_MUX_OUT_15_port, A(14) => WB_MUX_OUT_14_port, 
                           A(13) => WB_MUX_OUT_13_port, A(12) => 
                           WB_MUX_OUT_12_port, A(11) => WB_MUX_OUT_11_port, 
                           A(10) => WB_MUX_OUT_10_port, A(9) => 
                           WB_MUX_OUT_9_port, A(8) => WB_MUX_OUT_8_port, A(7) 
                           => WB_MUX_OUT_7_port, A(6) => WB_MUX_OUT_6_port, 
                           A(5) => WB_MUX_OUT_5_port, A(4) => WB_MUX_OUT_4_port
                           , A(3) => WB_MUX_OUT_3_port, A(2) => 
                           WB_MUX_OUT_2_port, A(1) => WB_MUX_OUT_1_port, A(0) 
                           => WB_MUX_OUT_0_port, B(31) => MEM_WB_NPC_31_port, 
                           B(30) => MEM_WB_NPC_30_port, B(29) => 
                           MEM_WB_NPC_29_port, B(28) => MEM_WB_NPC_28_port, 
                           B(27) => MEM_WB_NPC_27_port, B(26) => 
                           MEM_WB_NPC_26_port, B(25) => MEM_WB_NPC_25_port, 
                           B(24) => MEM_WB_NPC_24_port, B(23) => 
                           MEM_WB_NPC_23_port, B(22) => MEM_WB_NPC_22_port, 
                           B(21) => MEM_WB_NPC_21_port, B(20) => 
                           MEM_WB_NPC_20_port, B(19) => MEM_WB_NPC_19_port, 
                           B(18) => MEM_WB_NPC_18_port, B(17) => 
                           MEM_WB_NPC_17_port, B(16) => MEM_WB_NPC_16_port, 
                           B(15) => MEM_WB_NPC_15_port, B(14) => 
                           MEM_WB_NPC_14_port, B(13) => MEM_WB_NPC_13_port, 
                           B(12) => MEM_WB_NPC_12_port, B(11) => 
                           MEM_WB_NPC_11_port, B(10) => MEM_WB_NPC_10_port, 
                           B(9) => MEM_WB_NPC_9_port, B(8) => MEM_WB_NPC_8_port
                           , B(7) => MEM_WB_NPC_7_port, B(6) => 
                           MEM_WB_NPC_6_port, B(5) => MEM_WB_NPC_5_port, B(4) 
                           => MEM_WB_NPC_4_port, B(3) => MEM_WB_NPC_3_port, 
                           B(2) => MEM_WB_NPC_2_port, B(1) => MEM_WB_NPC_1_port
                           , B(0) => MEM_WB_NPC_0_port, S => JAL_MUX_SEL, Y(31)
                           => JAL_MUX_OUT_31_port, Y(30) => JAL_MUX_OUT_30_port
                           , Y(29) => JAL_MUX_OUT_29_port, Y(28) => 
                           JAL_MUX_OUT_28_port, Y(27) => JAL_MUX_OUT_27_port, 
                           Y(26) => JAL_MUX_OUT_26_port, Y(25) => 
                           JAL_MUX_OUT_25_port, Y(24) => JAL_MUX_OUT_24_port, 
                           Y(23) => JAL_MUX_OUT_23_port, Y(22) => 
                           JAL_MUX_OUT_22_port, Y(21) => JAL_MUX_OUT_21_port, 
                           Y(20) => JAL_MUX_OUT_20_port, Y(19) => 
                           JAL_MUX_OUT_19_port, Y(18) => JAL_MUX_OUT_18_port, 
                           Y(17) => JAL_MUX_OUT_17_port, Y(16) => 
                           JAL_MUX_OUT_16_port, Y(15) => JAL_MUX_OUT_15_port, 
                           Y(14) => JAL_MUX_OUT_14_port, Y(13) => 
                           JAL_MUX_OUT_13_port, Y(12) => JAL_MUX_OUT_12_port, 
                           Y(11) => JAL_MUX_OUT_11_port, Y(10) => 
                           JAL_MUX_OUT_10_port, Y(9) => JAL_MUX_OUT_9_port, 
                           Y(8) => JAL_MUX_OUT_8_port, Y(7) => 
                           JAL_MUX_OUT_7_port, Y(6) => JAL_MUX_OUT_6_port, Y(5)
                           => JAL_MUX_OUT_5_port, Y(4) => JAL_MUX_OUT_4_port, 
                           Y(3) => JAL_MUX_OUT_3_port, Y(2) => 
                           JAL_MUX_OUT_2_port, Y(1) => JAL_MUX_OUT_1_port, Y(0)
                           => JAL_MUX_OUT_0_port);
   add_630 : 
                           DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0 
                           port map( A(31) => PC_OUT_31_port, A(30) => 
                           PC_OUT_30_port, A(29) => PC_OUT_29_port, A(28) => 
                           PC_OUT_28_port, A(27) => PC_OUT_27_port, A(26) => 
                           PC_OUT_26_port, A(25) => PC_OUT_25_port, A(24) => 
                           PC_OUT_24_port, A(23) => PC_OUT_23_port, A(22) => 
                           PC_OUT_22_port, A(21) => PC_OUT_21_port, A(20) => 
                           PC_OUT_20_port, A(19) => PC_OUT_19_port, A(18) => 
                           PC_OUT_18_port, A(17) => PC_OUT_17_port, A(16) => 
                           PC_OUT_16_port, A(15) => PC_OUT_15_port, A(14) => 
                           PC_OUT_14_port, A(13) => PC_OUT_13_port, A(12) => 
                           PC_OUT_12_port, A(11) => PC_OUT_11_port, A(10) => 
                           PC_OUT_10_port, A(9) => PC_OUT_9_port, A(8) => 
                           PC_OUT_8_port, A(7) => PC_OUT_7_port, A(6) => 
                           PC_OUT_6_port, A(5) => PC_OUT_5_port, A(4) => 
                           PC_OUT_4_port, A(3) => PC_OUT_3_port, A(2) => 
                           PC_OUT_2_port, A(1) => PC_OUT_1_port, A(0) => 
                           PC_OUT_0_port, B(31) => n1, B(30) => n1, B(29) => n1
                           , B(28) => n1, B(27) => n1, B(26) => n1, B(25) => n1
                           , B(24) => n1, B(23) => n1, B(22) => n1, B(21) => n1
                           , B(20) => n1, B(19) => n1, B(18) => n1, B(17) => n1
                           , B(16) => n1, B(15) => n1, B(14) => n1, B(13) => n1
                           , B(12) => n1, B(11) => n1, B(10) => n1, B(9) => n1,
                           B(8) => n1, B(7) => n1, B(6) => n1, B(5) => n1, B(4)
                           => n1, B(3) => n1, B(2) => X_Logic1_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, CI => n1, 
                           SUM(31) => NPC_BUS_31_port, SUM(30) => 
                           NPC_BUS_30_port, SUM(29) => NPC_BUS_29_port, SUM(28)
                           => NPC_BUS_28_port, SUM(27) => NPC_BUS_27_port, 
                           SUM(26) => NPC_BUS_26_port, SUM(25) => 
                           NPC_BUS_25_port, SUM(24) => NPC_BUS_24_port, SUM(23)
                           => NPC_BUS_23_port, SUM(22) => NPC_BUS_22_port, 
                           SUM(21) => NPC_BUS_21_port, SUM(20) => 
                           NPC_BUS_20_port, SUM(19) => NPC_BUS_19_port, SUM(18)
                           => NPC_BUS_18_port, SUM(17) => NPC_BUS_17_port, 
                           SUM(16) => NPC_BUS_16_port, SUM(15) => 
                           NPC_BUS_15_port, SUM(14) => NPC_BUS_14_port, SUM(13)
                           => NPC_BUS_13_port, SUM(12) => NPC_BUS_12_port, 
                           SUM(11) => NPC_BUS_11_port, SUM(10) => 
                           NPC_BUS_10_port, SUM(9) => NPC_BUS_9_port, SUM(8) =>
                           NPC_BUS_8_port, SUM(7) => NPC_BUS_7_port, SUM(6) => 
                           NPC_BUS_6_port, SUM(5) => NPC_BUS_5_port, SUM(4) => 
                           NPC_BUS_4_port, SUM(3) => NPC_BUS_3_port, SUM(2) => 
                           NPC_BUS_2_port, SUM(1) => NPC_BUS_1_port, SUM(0) => 
                           NPC_BUS_0_port, CO => n_1705);
   IF_ID_IR_reg_31_inst : DFF_X1 port map( D => N65, CK => CLK, Q => 
                           IF_ID_IR_31_port, QN => n7_port);
   IF_ID_IR_reg_28_inst : DFF_X1 port map( D => N62, CK => CLK, Q => 
                           IF_ID_IR_28_port, QN => n_1706);
   ID_EX_RS2_reg_3_inst : DFF_X2 port map( D => N107, CK => CLK, Q => 
                           ID_EX_RS2_3_port, QN => n_1707);
   ID_EX_RS2_reg_2_inst : DFF_X2 port map( D => N106, CK => CLK, Q => 
                           ID_EX_RS2_2_port, QN => n_1708);
   ID_EX_RS1_reg_4_inst : DFF_X1 port map( D => N103, CK => CLK, Q => 
                           ID_EX_RS1_4_port, QN => n_1709);
   ID_EX_RS2_reg_4_inst : DFF_X2 port map( D => N108, CK => CLK, Q => 
                           ID_EX_RS2_4_port, QN => n_1710);
   ID_EX_RS2_reg_0_inst : DFF_X2 port map( D => N104, CK => CLK, Q => 
                           ID_EX_RS2_0_port, QN => n_1711);
   ID_EX_RS2_reg_1_inst : DFF_X2 port map( D => N105, CK => CLK, Q => 
                           ID_EX_RS2_1_port, QN => n_1712);
   ID_EX_RD_reg_2_inst : DFF_X1 port map( D => N111, CK => CLK, Q => 
                           ID_EX_RD_2_port, QN => n_1713);
   ID_EX_RD_reg_0_inst : DFF_X1 port map( D => N109, CK => CLK, Q => 
                           ID_EX_RD_0_port, QN => n_1714);
   ID_EX_RD_reg_4_inst : DFF_X1 port map( D => N113, CK => CLK, Q => 
                           ID_EX_RD_4_port, QN => n_1715);
   U3 : CLKBUF_X1 port map( A => ID_EX_RS1_NEXT_0_port, Z => n2_port);
   U5 : CLKBUF_X1 port map( A => ID_EX_RS1_NEXT_4_port, Z => n3_port);
   U6 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_3_port, A2 => RST, ZN => N107);
   U7 : CLKBUF_X1 port map( A => ID_EX_RS2_NEXT_3_port, Z => net31024);
   U8 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_2_port, A2 => RST, ZN => N106);
   U9 : CLKBUF_X1 port map( A => ID_EX_RS2_NEXT_2_port, Z => net31028);
   U10 : INV_X1 port map( A => n4_port, ZN => n6_port);
   U11 : INV_X1 port map( A => n7_port, ZN => n8_port);
   U12 : INV_X1 port map( A => n9_port, ZN => n10_port);
   U13 : BUF_X1 port map( A => RST, Z => net31092);
   U14 : BUF_X1 port map( A => RST, Z => net31090);
   U15 : BUF_X1 port map( A => RST, Z => net31098);
   U16 : BUF_X1 port map( A => RST, Z => net31094);
   U17 : BUF_X1 port map( A => RST, Z => net31096);
   U18 : BUF_X2 port map( A => RST, Z => net31258);
   U19 : BUF_X1 port map( A => net31098, Z => net31062);
   U20 : BUF_X1 port map( A => net31098, Z => net31064);
   U21 : BUF_X1 port map( A => net31098, Z => net31060);
   U22 : BUF_X1 port map( A => RST, Z => net31054);
   U23 : BUF_X1 port map( A => net31092, Z => net31082);
   U24 : BUF_X1 port map( A => RST, Z => net31056);
   U25 : BUF_X1 port map( A => net31090, Z => net31084);
   U26 : BUF_X1 port map( A => RST, Z => net31058);
   U27 : BUF_X1 port map( A => net31092, Z => net31080);
   U28 : BUF_X1 port map( A => net31092, Z => net31078);
   U29 : BUF_X1 port map( A => net31090, Z => net31086);
   U30 : BUF_X1 port map( A => net31094, Z => net31076);
   U31 : BUF_X1 port map( A => net31094, Z => net31074);
   U32 : BUF_X1 port map( A => net31094, Z => net31072);
   U33 : BUF_X1 port map( A => net31096, Z => net31070);
   U34 : BUF_X1 port map( A => net31096, Z => net31068);
   U35 : BUF_X1 port map( A => net31096, Z => net31066);
   U36 : BUF_X1 port map( A => RST, Z => net31046);
   U37 : BUF_X1 port map( A => RST, Z => net31044);
   U38 : BUF_X1 port map( A => net31090, Z => net31088);
   U39 : BUF_X4 port map( A => RST, Z => net31260);
   U40 : INV_X1 port map( A => ZERO_OUT, ZN => n18_port);
   U41 : AND2_X1 port map( A1 => RST, A2 => ID_EX_RS1_NEXT_0_port, ZN => N99);
   U42 : AND2_X1 port map( A1 => ID_EX_RS1_NEXT_4_port, A2 => RST, ZN => N103);
   U43 : AND2_X1 port map( A1 => ID_EX_RS1_NEXT_2_port, A2 => RST, ZN => N101);
   U44 : AND2_X1 port map( A1 => ID_EX_RS1_NEXT_1_port, A2 => RST, ZN => N100);
   U45 : AND2_X1 port map( A1 => ID_EX_RS1_NEXT_3_port, A2 => RST, ZN => N102);
   U46 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_0_port, A2 => RST, ZN => N109);
   U47 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_1_port, A2 => RST, ZN => N110);
   U48 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_2_port, A2 => RST, ZN => N111);
   U49 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_3_port, A2 => RST, ZN => N112);
   U50 : AND2_X1 port map( A1 => ALU_OUT_9_port, A2 => net31260, ZN => N355);
   U51 : AND2_X1 port map( A1 => ALU_OUT_31_port, A2 => net31260, ZN => N377);
   U52 : AND2_X1 port map( A1 => ALU_OUT_30_port, A2 => net31260, ZN => N376);
   U53 : AND2_X1 port map( A1 => ALU_OUT_29_port, A2 => net31260, ZN => N375);
   U54 : AND2_X1 port map( A1 => ALU_OUT_28_port, A2 => net31260, ZN => N374);
   U55 : AND2_X1 port map( A1 => ALU_OUT_27_port, A2 => net31260, ZN => N373);
   U56 : AND2_X1 port map( A1 => ALU_OUT_26_port, A2 => net31260, ZN => N372);
   U57 : AND2_X1 port map( A1 => ALU_OUT_25_port, A2 => net31260, ZN => N371);
   U58 : AND2_X1 port map( A1 => ALU_OUT_24_port, A2 => net31260, ZN => N370);
   U59 : AND2_X1 port map( A1 => ALU_OUT_23_port, A2 => net31260, ZN => N369);
   U60 : AND2_X1 port map( A1 => ALU_OUT_22_port, A2 => net31260, ZN => N368);
   U61 : AND2_X1 port map( A1 => ALU_OUT_21_port, A2 => net31260, ZN => N367);
   U62 : AND2_X1 port map( A1 => ALU_OUT_20_port, A2 => net31260, ZN => N366);
   U63 : AND2_X1 port map( A1 => ALU_OUT_19_port, A2 => net31260, ZN => N365);
   U64 : AND2_X1 port map( A1 => ALU_OUT_18_port, A2 => net31260, ZN => N364);
   U65 : AND2_X1 port map( A1 => ALU_OUT_17_port, A2 => net31260, ZN => N363);
   U66 : AND2_X1 port map( A1 => ALU_OUT_16_port, A2 => net31260, ZN => N362);
   U67 : AND2_X1 port map( A1 => ALU_OUT_15_port, A2 => net31260, ZN => N361);
   U68 : AND2_X1 port map( A1 => ALU_OUT_14_port, A2 => net31260, ZN => N360);
   U69 : AND2_X1 port map( A1 => ALU_OUT_13_port, A2 => net31260, ZN => N359);
   U70 : AND2_X1 port map( A1 => ALU_OUT_12_port, A2 => net31260, ZN => N358);
   U71 : AND2_X1 port map( A1 => ALU_OUT_11_port, A2 => net31260, ZN => N357);
   U72 : AND2_X1 port map( A1 => ALU_OUT_10_port, A2 => net31260, ZN => N356);
   U73 : AND2_X1 port map( A1 => ALU_OUT_8_port, A2 => net31260, ZN => N354);
   U74 : AND2_X1 port map( A1 => ALU_OUT_7_port, A2 => net31260, ZN => N353);
   U75 : AND2_X1 port map( A1 => ALU_OUT_6_port, A2 => net31260, ZN => N352);
   U76 : AND2_X1 port map( A1 => ALU_OUT_5_port, A2 => net31260, ZN => N351);
   U77 : AND2_X1 port map( A1 => ALU_OUT_4_port, A2 => net31260, ZN => N350);
   U78 : AND2_X1 port map( A1 => ALU_OUT_3_port, A2 => net31260, ZN => N349);
   U79 : AND2_X1 port map( A1 => ALU_OUT_2_port, A2 => net31260, ZN => N348);
   U80 : AND2_X1 port map( A1 => ALU_OUT_1_port, A2 => net31260, ZN => N347);
   U81 : AND2_X1 port map( A1 => ALU_OUT_0_port, A2 => net31260, ZN => N346);
   U82 : AND2_X1 port map( A1 => EX_MEM_RD_0_port, A2 => net31070, ZN => N410);
   U83 : AND2_X1 port map( A1 => EX_MEM_RD_1_port, A2 => net31070, ZN => N411);
   U84 : AND2_X1 port map( A1 => EX_MEM_RD_2_port, A2 => net31070, ZN => N412);
   U85 : AND2_X1 port map( A1 => EX_MEM_RD_3_port, A2 => net31070, ZN => N413);
   U86 : AND2_X1 port map( A1 => EX_MEM_RD_4_port, A2 => net31070, ZN => N414);
   U87 : AND2_X1 port map( A1 => ID_EX_NPC_9_port, A2 => net31064, ZN => N219);
   U88 : AND2_X1 port map( A1 => ID_EX_NPC_31_port, A2 => net31058, ZN => N241)
                           ;
   U89 : AND2_X1 port map( A1 => ID_EX_NPC_30_port, A2 => net31058, ZN => N240)
                           ;
   U90 : AND2_X1 port map( A1 => ID_EX_NPC_29_port, A2 => net31060, ZN => N239)
                           ;
   U91 : AND2_X1 port map( A1 => ID_EX_NPC_28_port, A2 => net31060, ZN => N238)
                           ;
   U92 : AND2_X1 port map( A1 => ID_EX_NPC_27_port, A2 => net31060, ZN => N237)
                           ;
   U93 : AND2_X1 port map( A1 => ID_EX_NPC_26_port, A2 => net31060, ZN => N236)
                           ;
   U94 : AND2_X1 port map( A1 => ID_EX_NPC_25_port, A2 => net31060, ZN => N235)
                           ;
   U95 : AND2_X1 port map( A1 => ID_EX_NPC_24_port, A2 => net31060, ZN => N234)
                           ;
   U96 : AND2_X1 port map( A1 => ID_EX_NPC_23_port, A2 => net31060, ZN => N233)
                           ;
   U97 : AND2_X1 port map( A1 => ID_EX_NPC_22_port, A2 => net31060, ZN => N232)
                           ;
   U98 : AND2_X1 port map( A1 => ID_EX_NPC_21_port, A2 => net31060, ZN => N231)
                           ;
   U99 : AND2_X1 port map( A1 => ID_EX_NPC_20_port, A2 => net31062, ZN => N230)
                           ;
   U100 : AND2_X1 port map( A1 => ID_EX_NPC_19_port, A2 => net31062, ZN => N229
                           );
   U101 : AND2_X1 port map( A1 => ID_EX_NPC_18_port, A2 => net31062, ZN => N228
                           );
   U102 : AND2_X1 port map( A1 => ID_EX_NPC_17_port, A2 => net31062, ZN => N227
                           );
   U103 : AND2_X1 port map( A1 => ID_EX_NPC_16_port, A2 => net31062, ZN => N226
                           );
   U104 : AND2_X1 port map( A1 => ID_EX_NPC_15_port, A2 => net31062, ZN => N225
                           );
   U105 : AND2_X1 port map( A1 => ID_EX_NPC_14_port, A2 => net31062, ZN => N224
                           );
   U106 : AND2_X1 port map( A1 => ID_EX_NPC_13_port, A2 => net31062, ZN => N223
                           );
   U107 : AND2_X1 port map( A1 => ID_EX_NPC_12_port, A2 => net31062, ZN => N222
                           );
   U108 : AND2_X1 port map( A1 => ID_EX_NPC_11_port, A2 => net31062, ZN => N221
                           );
   U109 : AND2_X1 port map( A1 => ID_EX_NPC_10_port, A2 => net31064, ZN => N220
                           );
   U110 : AND2_X1 port map( A1 => ID_EX_NPC_8_port, A2 => net31064, ZN => N218)
                           ;
   U111 : AND2_X1 port map( A1 => ID_EX_NPC_7_port, A2 => net31064, ZN => N217)
                           ;
   U112 : AND2_X1 port map( A1 => ID_EX_NPC_6_port, A2 => net31064, ZN => N216)
                           ;
   U113 : AND2_X1 port map( A1 => ID_EX_NPC_5_port, A2 => net31064, ZN => N215)
                           ;
   U114 : AND2_X1 port map( A1 => ID_EX_NPC_4_port, A2 => net31064, ZN => N214)
                           ;
   U115 : AND2_X1 port map( A1 => ID_EX_NPC_3_port, A2 => net31064, ZN => N213)
                           ;
   U116 : AND2_X1 port map( A1 => ID_EX_NPC_2_port, A2 => net31064, ZN => N212)
                           ;
   U117 : AND2_X1 port map( A1 => ID_EX_NPC_1_port, A2 => net31064, ZN => N211)
                           ;
   U118 : AND2_X1 port map( A1 => ID_EX_NPC_0_port, A2 => net31066, ZN => N210)
                           ;
   U119 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_31_port, A2 => RST, ZN => N274)
                           ;
   U120 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_30_port, A2 => RST, ZN => N273)
                           ;
   U121 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_29_port, A2 => RST, ZN => N272)
                           ;
   U122 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_28_port, A2 => RST, ZN => N271)
                           ;
   U123 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_27_port, A2 => RST, ZN => N270)
                           ;
   U124 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_26_port, A2 => net31054, ZN => 
                           N269);
   U125 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_25_port, A2 => net31054, ZN => 
                           N268);
   U126 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_24_port, A2 => net31054, ZN => 
                           N267);
   U127 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_23_port, A2 => net31054, ZN => 
                           N266);
   U128 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_22_port, A2 => net31054, ZN => 
                           N265);
   U129 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_21_port, A2 => net31054, ZN => 
                           N264);
   U130 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_20_port, A2 => net31054, ZN => 
                           N263);
   U131 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_19_port, A2 => net31054, ZN => 
                           N262);
   U132 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_18_port, A2 => net31054, ZN => 
                           N261);
   U133 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_17_port, A2 => net31054, ZN => 
                           N260);
   U134 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_16_port, A2 => net31056, ZN => 
                           N259);
   U135 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_15_port, A2 => net31056, ZN => 
                           N258);
   U136 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_14_port, A2 => net31056, ZN => 
                           N257);
   U137 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_13_port, A2 => net31056, ZN => 
                           N256);
   U138 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_12_port, A2 => net31056, ZN => 
                           N255);
   U139 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_11_port, A2 => net31056, ZN => 
                           N254);
   U140 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_10_port, A2 => net31056, ZN => 
                           N253);
   U141 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_9_port, A2 => net31056, ZN => 
                           N252);
   U142 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_8_port, A2 => net31056, ZN => 
                           N251);
   U143 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_7_port, A2 => net31056, ZN => 
                           N250);
   U144 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_6_port, A2 => net31058, ZN => 
                           N249);
   U145 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_5_port, A2 => net31058, ZN => 
                           N248);
   U146 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_4_port, A2 => net31058, ZN => 
                           N247);
   U147 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_3_port, A2 => net31058, ZN => 
                           N246);
   U148 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_2_port, A2 => net31058, ZN => 
                           N245);
   U149 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_1_port, A2 => net31058, ZN => 
                           N244);
   U150 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_0_port, A2 => net31058, ZN => 
                           N243);
   U151 : AND2_X1 port map( A1 => EX_MEM_RF_WE, A2 => net31260, ZN => N345);
   U152 : AND2_X1 port map( A1 => IF_ID_NPC_20_port, A2 => net31258, ZN => N86)
                           ;
   U153 : AND2_X1 port map( A1 => IF_ID_NPC_19_port, A2 => net31258, ZN => N85)
                           ;
   U154 : AND2_X1 port map( A1 => IF_ID_NPC_18_port, A2 => net31258, ZN => N84)
                           ;
   U155 : AND2_X1 port map( A1 => IF_ID_NPC_17_port, A2 => net31258, ZN => N83)
                           ;
   U156 : AND2_X1 port map( A1 => IF_ID_NPC_16_port, A2 => net31258, ZN => N82)
                           ;
   U157 : AND2_X1 port map( A1 => IF_ID_NPC_15_port, A2 => net31258, ZN => N81)
                           ;
   U158 : AND2_X1 port map( A1 => IF_ID_NPC_14_port, A2 => net31258, ZN => N80)
                           ;
   U159 : AND2_X1 port map( A1 => IF_ID_NPC_13_port, A2 => net31258, ZN => N79)
                           ;
   U160 : AND2_X1 port map( A1 => IF_ID_NPC_12_port, A2 => net31258, ZN => N78)
                           ;
   U161 : AND2_X1 port map( A1 => IF_ID_NPC_11_port, A2 => net31258, ZN => N77)
                           ;
   U162 : AND2_X1 port map( A1 => IF_ID_NPC_10_port, A2 => net31258, ZN => N76)
                           ;
   U163 : AND2_X1 port map( A1 => IF_ID_NPC_9_port, A2 => net31258, ZN => N75);
   U164 : AND2_X1 port map( A1 => IF_ID_NPC_8_port, A2 => net31258, ZN => N74);
   U165 : AND2_X1 port map( A1 => IF_ID_NPC_7_port, A2 => net31258, ZN => N73);
   U166 : AND2_X1 port map( A1 => IF_ID_NPC_6_port, A2 => net31258, ZN => N72);
   U167 : AND2_X1 port map( A1 => IF_ID_NPC_5_port, A2 => net31258, ZN => N71);
   U168 : AND2_X1 port map( A1 => IF_ID_NPC_4_port, A2 => net31258, ZN => N70);
   U169 : AND2_X1 port map( A1 => IF_ID_NPC_3_port, A2 => net31258, ZN => N69);
   U170 : AND2_X1 port map( A1 => IF_ID_NPC_2_port, A2 => net31258, ZN => N68);
   U171 : AND2_X1 port map( A1 => IF_ID_NPC_1_port, A2 => net31258, ZN => N67);
   U172 : AND2_X1 port map( A1 => IF_ID_NPC_0_port, A2 => net31258, ZN => N66);
   U173 : AND2_X1 port map( A1 => EX_MEM_NPC_31_port, A2 => net31260, ZN => 
                           N344);
   U174 : AND2_X1 port map( A1 => IF_ID_NPC_31_port, A2 => net31260, ZN => N97)
                           ;
   U175 : AND2_X1 port map( A1 => EX_MEM_NPC_30_port, A2 => net31260, ZN => 
                           N343);
   U176 : AND2_X1 port map( A1 => IF_ID_NPC_30_port, A2 => net31260, ZN => N96)
                           ;
   U177 : AND2_X1 port map( A1 => EX_MEM_NPC_29_port, A2 => net31260, ZN => 
                           N342);
   U178 : AND2_X1 port map( A1 => IF_ID_NPC_29_port, A2 => net31260, ZN => N95)
                           ;
   U179 : AND2_X1 port map( A1 => EX_MEM_NPC_28_port, A2 => net31260, ZN => 
                           N341);
   U180 : AND2_X1 port map( A1 => IF_ID_NPC_28_port, A2 => net31260, ZN => N94)
                           ;
   U181 : AND2_X1 port map( A1 => EX_MEM_NPC_27_port, A2 => net31260, ZN => 
                           N340);
   U182 : AND2_X1 port map( A1 => IF_ID_NPC_27_port, A2 => net31260, ZN => N93)
                           ;
   U183 : AND2_X1 port map( A1 => EX_MEM_NPC_26_port, A2 => net31260, ZN => 
                           N339);
   U184 : AND2_X1 port map( A1 => IF_ID_NPC_26_port, A2 => net31260, ZN => N92)
                           ;
   U185 : AND2_X1 port map( A1 => EX_MEM_NPC_25_port, A2 => net31260, ZN => 
                           N338);
   U186 : AND2_X1 port map( A1 => IF_ID_NPC_25_port, A2 => net31260, ZN => N91)
                           ;
   U187 : AND2_X1 port map( A1 => EX_MEM_NPC_24_port, A2 => net31260, ZN => 
                           N337);
   U188 : AND2_X1 port map( A1 => IF_ID_NPC_24_port, A2 => net31260, ZN => N90)
                           ;
   U189 : AND2_X1 port map( A1 => EX_MEM_NPC_23_port, A2 => net31260, ZN => 
                           N336);
   U190 : AND2_X1 port map( A1 => IF_ID_NPC_23_port, A2 => net31260, ZN => N89)
                           ;
   U191 : AND2_X1 port map( A1 => EX_MEM_NPC_22_port, A2 => net31260, ZN => 
                           N335);
   U192 : AND2_X1 port map( A1 => IF_ID_NPC_22_port, A2 => net31260, ZN => N88)
                           ;
   U193 : AND2_X1 port map( A1 => EX_MEM_NPC_21_port, A2 => net31260, ZN => 
                           N334);
   U194 : AND2_X1 port map( A1 => IF_ID_NPC_21_port, A2 => net31260, ZN => N87)
                           ;
   U195 : AND2_X1 port map( A1 => EX_MEM_NPC_20_port, A2 => net31260, ZN => 
                           N333);
   U196 : AND2_X1 port map( A1 => EX_MEM_NPC_19_port, A2 => net31260, ZN => 
                           N332);
   U197 : AND2_X1 port map( A1 => EX_MEM_NPC_18_port, A2 => net31260, ZN => 
                           N331);
   U198 : AND2_X1 port map( A1 => EX_MEM_NPC_17_port, A2 => net31260, ZN => 
                           N330);
   U199 : AND2_X1 port map( A1 => EX_MEM_NPC_16_port, A2 => net31260, ZN => 
                           N329);
   U200 : AND2_X1 port map( A1 => EX_MEM_NPC_15_port, A2 => net31260, ZN => 
                           N328);
   U201 : AND2_X1 port map( A1 => EX_MEM_NPC_14_port, A2 => net31260, ZN => 
                           N327);
   U202 : AND2_X1 port map( A1 => EX_MEM_NPC_13_port, A2 => net31260, ZN => 
                           N326);
   U203 : AND2_X1 port map( A1 => EX_MEM_NPC_12_port, A2 => net31260, ZN => 
                           N325);
   U204 : AND2_X1 port map( A1 => EX_MEM_NPC_11_port, A2 => net31260, ZN => 
                           N324);
   U205 : AND2_X1 port map( A1 => EX_MEM_NPC_10_port, A2 => net31260, ZN => 
                           N323);
   U206 : AND2_X1 port map( A1 => EX_MEM_NPC_9_port, A2 => net31260, ZN => N322
                           );
   U207 : AND2_X1 port map( A1 => EX_MEM_NPC_8_port, A2 => net31260, ZN => N321
                           );
   U208 : AND2_X1 port map( A1 => EX_MEM_NPC_7_port, A2 => net31260, ZN => N320
                           );
   U209 : AND2_X1 port map( A1 => EX_MEM_NPC_6_port, A2 => net31260, ZN => N319
                           );
   U210 : AND2_X1 port map( A1 => EX_MEM_NPC_5_port, A2 => net31260, ZN => N318
                           );
   U211 : AND2_X1 port map( A1 => EX_MEM_NPC_4_port, A2 => net31260, ZN => N317
                           );
   U212 : AND2_X1 port map( A1 => EX_MEM_NPC_3_port, A2 => net31260, ZN => N316
                           );
   U213 : AND2_X1 port map( A1 => EX_MEM_NPC_2_port, A2 => net31260, ZN => N315
                           );
   U214 : AND2_X1 port map( A1 => EX_MEM_NPC_1_port, A2 => net31260, ZN => N314
                           );
   U215 : AND2_X1 port map( A1 => EX_MEM_NPC_0_port, A2 => net31260, ZN => N313
                           );
   U216 : AND2_X1 port map( A1 => ID_EX_RD_0_port, A2 => net31260, ZN => N308);
   U217 : AND2_X1 port map( A1 => ID_EX_RD_1_port, A2 => net31260, ZN => N309);
   U218 : AND2_X1 port map( A1 => ID_EX_RD_2_port, A2 => net31260, ZN => N310);
   U219 : AND2_X1 port map( A1 => ID_EX_RD_3_port, A2 => net31260, ZN => N311);
   U220 : AND2_X1 port map( A1 => ID_EX_RD_4_port, A2 => net31260, ZN => N312);
   U221 : AND2_X1 port map( A1 => ID_EX_RF_WE, A2 => net31058, ZN => N242);
   U222 : AND2_X1 port map( A1 => IR_OUT_0_port, A2 => net31260, ZN => N34);
   U223 : AND2_X1 port map( A1 => IR_OUT_3_port, A2 => net31260, ZN => N37);
   U224 : INV_X1 port map( A => n5_port, ZN => n19_port);
   U225 : AOI21_X1 port map( B1 => JUMP_EN, B2 => EX_MEM_BRANCH_DETECT, A => 
                           JUMP_COND, ZN => n5_port);
   U226 : AND2_X1 port map( A1 => IR_OUT_1_port, A2 => net31260, ZN => N35);
   U227 : AND2_X1 port map( A1 => IR_OUT_31_port, A2 => net31258, ZN => N65);
   U228 : AND2_X1 port map( A1 => IR_OUT_29_port, A2 => net31258, ZN => N63);
   U229 : AND2_X1 port map( A1 => IR_OUT_2_port, A2 => net31260, ZN => N36);
   U230 : AND2_X1 port map( A1 => IR_OUT_27_port, A2 => net31066, ZN => N61);
   U231 : AND2_X1 port map( A1 => IR_OUT_30_port, A2 => net31258, ZN => N64);
   U232 : AND2_X1 port map( A1 => IR_OUT_26_port, A2 => net31044, ZN => N60);
   U233 : AND2_X1 port map( A1 => IR_OUT_28_port, A2 => net31258, ZN => N62);
   U234 : AND2_X1 port map( A1 => IR_OUT_4_port, A2 => net31076, ZN => N38);
   U235 : AND2_X1 port map( A1 => IR_OUT_5_port, A2 => net31074, ZN => N39);
   U236 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_8_port, A2 => net31258, ZN => 
                           N10);
   U237 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_6_port, A2 => net31258, ZN => 
                           N8);
   U238 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_5_port, A2 => net31258, ZN => 
                           N7);
   U239 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_31_port, A2 => net31260, ZN =>
                           N33);
   U240 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_30_port, A2 => net31260, ZN =>
                           N32);
   U241 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_29_port, A2 => net31260, ZN =>
                           N31);
   U242 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_28_port, A2 => net31260, ZN =>
                           N30);
   U243 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_27_port, A2 => net31260, ZN =>
                           N29);
   U244 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_7_port, A2 => net31260, ZN => 
                           N9);
   U245 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_1_port, A2 => net31260, ZN => 
                           N3);
   U246 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_31_port, A2 => 
                           net31260, ZN => N306);
   U247 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_30_port, A2 => 
                           net31260, ZN => N305);
   U248 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_29_port, A2 => 
                           net31260, ZN => N304);
   U249 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_28_port, A2 => 
                           net31260, ZN => N303);
   U250 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_27_port, A2 => 
                           net31260, ZN => N302);
   U251 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_26_port, A2 => 
                           net31260, ZN => N301);
   U252 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_25_port, A2 => 
                           net31260, ZN => N300);
   U253 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_24_port, A2 => 
                           net31260, ZN => N299);
   U254 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_23_port, A2 => 
                           net31260, ZN => N298);
   U255 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_22_port, A2 => 
                           net31260, ZN => N297);
   U256 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_21_port, A2 => 
                           net31260, ZN => N296);
   U257 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_20_port, A2 => 
                           net31260, ZN => N295);
   U258 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_19_port, A2 => 
                           net31260, ZN => N294);
   U259 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_18_port, A2 => 
                           net31260, ZN => N293);
   U260 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_17_port, A2 => 
                           net31260, ZN => N292);
   U261 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_16_port, A2 => 
                           net31260, ZN => N291);
   U262 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_15_port, A2 => 
                           net31260, ZN => N290);
   U263 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_14_port, A2 => 
                           net31260, ZN => N289);
   U264 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_13_port, A2 => 
                           net31260, ZN => N288);
   U265 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_12_port, A2 => 
                           net31260, ZN => N287);
   U266 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_11_port, A2 => 
                           net31260, ZN => N286);
   U267 : AND2_X1 port map( A1 => EX_MEM_BRANCH_DETECT_NEXT, A2 => net31260, ZN
                           => N307);
   U268 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_1_port, A2 => 
                           net31260, ZN => N379);
   U269 : AND2_X1 port map( A1 => IR_OUT_10_port, A2 => net31068, ZN => N44);
   U270 : AND2_X1 port map( A1 => IR_OUT_6_port, A2 => net31072, ZN => N40);
   U271 : AND2_X1 port map( A1 => IR_OUT_7_port, A2 => net31070, ZN => N41);
   U272 : AND2_X1 port map( A1 => IR_OUT_8_port, A2 => net31070, ZN => N42);
   U273 : AND2_X1 port map( A1 => IR_OUT_9_port, A2 => net31070, ZN => N43);
   U274 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_26_port, A2 => RST, ZN => N28)
                           ;
   U275 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_25_port, A2 => RST, ZN => N27)
                           ;
   U276 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_24_port, A2 => net31056, ZN =>
                           N26);
   U277 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_23_port, A2 => net31058, ZN =>
                           N25);
   U278 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_22_port, A2 => net31060, ZN =>
                           N24);
   U279 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_21_port, A2 => net31062, ZN =>
                           N23);
   U280 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_20_port, A2 => net31064, ZN =>
                           N22);
   U281 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_19_port, A2 => net31066, ZN =>
                           N21);
   U282 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_18_port, A2 => RST, ZN => N20)
                           ;
   U283 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_17_port, A2 => net31078, ZN =>
                           N19);
   U284 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_16_port, A2 => net31080, ZN =>
                           N18);
   U285 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_15_port, A2 => net31082, ZN =>
                           N17);
   U286 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_14_port, A2 => net31084, ZN =>
                           N16);
   U287 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_13_port, A2 => net31086, ZN =>
                           N15);
   U288 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_12_port, A2 => net31088, ZN =>
                           N14);
   U289 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_11_port, A2 => net31044, ZN =>
                           N13);
   U290 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_10_port, A2 => net31046, ZN =>
                           N12);
   U291 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_9_port, A2 => RST, ZN => N11);
   U292 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_4_port, A2 => net31076, ZN => 
                           N6);
   U293 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_3_port, A2 => net31068, ZN => 
                           N5);
   U294 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_2_port, A2 => net31072, ZN => 
                           N4);
   U295 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_0_port, A2 => RST, ZN => N2);
   U296 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_10_port, A2 => 
                           net31060, ZN => N285);
   U297 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_9_port, A2 => RST, ZN 
                           => N284);
   U298 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_8_port, A2 => RST, ZN 
                           => N283);
   U299 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_7_port, A2 => RST, ZN 
                           => N282);
   U300 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_6_port, A2 => RST, ZN 
                           => N281);
   U301 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_5_port, A2 => RST, ZN 
                           => N280);
   U302 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_4_port, A2 => RST, ZN 
                           => N279);
   U303 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_3_port, A2 => RST, ZN 
                           => N278);
   U304 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_2_port, A2 => RST, ZN 
                           => N277);
   U305 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_1_port, A2 => RST, ZN 
                           => N276);
   U306 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_0_port, A2 => RST, ZN 
                           => N275);
   U307 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_31_port, A2 => net31086, 
                           ZN => N145);
   U308 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_30_port, A2 => net31086, 
                           ZN => N144);
   U309 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_29_port, A2 => net31088, 
                           ZN => N143);
   U310 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_28_port, A2 => net31088, 
                           ZN => N142);
   U311 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_27_port, A2 => net31088, 
                           ZN => N141);
   U312 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_26_port, A2 => net31088, 
                           ZN => N140);
   U313 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_25_port, A2 => net31088, 
                           ZN => N139);
   U314 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_24_port, A2 => net31088, 
                           ZN => N138);
   U315 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_23_port, A2 => net31054, 
                           ZN => N137);
   U316 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_22_port, A2 => net31044, 
                           ZN => N136);
   U317 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_21_port, A2 => net31044, 
                           ZN => N135);
   U318 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_20_port, A2 => net31044, 
                           ZN => N134);
   U319 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_19_port, A2 => net31044, 
                           ZN => N133);
   U320 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_18_port, A2 => net31044, 
                           ZN => N132);
   U321 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_17_port, A2 => net31044, 
                           ZN => N131);
   U322 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_16_port, A2 => net31044, 
                           ZN => N130);
   U323 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_15_port, A2 => net31044, 
                           ZN => N129);
   U324 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_14_port, A2 => net31044, 
                           ZN => N128);
   U325 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_13_port, A2 => net31046, 
                           ZN => N127);
   U326 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_12_port, A2 => net31046, 
                           ZN => N126);
   U327 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_11_port, A2 => net31046, 
                           ZN => N125);
   U328 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_10_port, A2 => net31046, 
                           ZN => N124);
   U329 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_9_port, A2 => net31046, ZN
                           => N123);
   U330 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_8_port, A2 => net31046, ZN
                           => N122);
   U331 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_7_port, A2 => net31046, ZN
                           => N121);
   U332 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_6_port, A2 => net31046, ZN
                           => N120);
   U333 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_5_port, A2 => net31046, ZN
                           => N119);
   U334 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_4_port, A2 => net31046, ZN
                           => N118);
   U335 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_3_port, A2 => RST, ZN => 
                           N117);
   U336 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_2_port, A2 => RST, ZN => 
                           N116);
   U337 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_1_port, A2 => RST, ZN => 
                           N115);
   U338 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_0_port, A2 => RST, ZN => 
                           N114);
   U339 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_31_port, A2 => net31080, 
                           ZN => N177);
   U340 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_30_port, A2 => net31080, 
                           ZN => N176);
   U341 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_29_port, A2 => net31080, 
                           ZN => N175);
   U342 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_28_port, A2 => net31080, 
                           ZN => N174);
   U343 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_27_port, A2 => net31080, 
                           ZN => N173);
   U344 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_26_port, A2 => net31082, 
                           ZN => N172);
   U345 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_25_port, A2 => net31082, 
                           ZN => N171);
   U346 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_24_port, A2 => net31082, 
                           ZN => N170);
   U347 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_23_port, A2 => net31082, 
                           ZN => N169);
   U348 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_22_port, A2 => net31082, 
                           ZN => N168);
   U349 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_21_port, A2 => net31082, 
                           ZN => N167);
   U350 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_20_port, A2 => net31082, 
                           ZN => N166);
   U351 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_19_port, A2 => net31082, 
                           ZN => N165);
   U352 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_18_port, A2 => net31082, 
                           ZN => N164);
   U353 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_17_port, A2 => net31082, 
                           ZN => N163);
   U354 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_16_port, A2 => net31084, 
                           ZN => N162);
   U355 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_15_port, A2 => net31084, 
                           ZN => N161);
   U356 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_14_port, A2 => net31084, 
                           ZN => N160);
   U357 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_13_port, A2 => net31084, 
                           ZN => N159);
   U358 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_12_port, A2 => net31084, 
                           ZN => N158);
   U359 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_11_port, A2 => net31084, 
                           ZN => N157);
   U360 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_10_port, A2 => net31084, 
                           ZN => N156);
   U361 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_9_port, A2 => net31084, ZN
                           => N155);
   U362 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_8_port, A2 => net31084, ZN
                           => N154);
   U363 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_7_port, A2 => net31084, ZN
                           => N153);
   U364 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_6_port, A2 => net31086, ZN
                           => N152);
   U365 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_5_port, A2 => net31086, ZN
                           => N151);
   U366 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_4_port, A2 => net31086, ZN
                           => N150);
   U367 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_3_port, A2 => net31086, ZN
                           => N149);
   U368 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_2_port, A2 => net31086, ZN
                           => N148);
   U369 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_1_port, A2 => net31086, ZN
                           => N147);
   U370 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_0_port, A2 => net31086, ZN
                           => N146);
   U371 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_0_port, A2 => 
                           net31076, ZN => N378);
   U372 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_2_port, A2 => 
                           net31076, ZN => N380);
   U373 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_3_port, A2 => 
                           net31076, ZN => N381);
   U374 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_4_port, A2 => 
                           net31076, ZN => N382);
   U375 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_5_port, A2 => 
                           net31076, ZN => N383);
   U376 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_6_port, A2 => 
                           net31076, ZN => N384);
   U377 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_7_port, A2 => 
                           net31076, ZN => N385);
   U378 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_8_port, A2 => 
                           net31076, ZN => N386);
   U379 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_9_port, A2 => 
                           net31076, ZN => N387);
   U380 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_10_port, A2 => 
                           net31074, ZN => N388);
   U381 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_11_port, A2 => 
                           net31074, ZN => N389);
   U382 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_12_port, A2 => 
                           net31074, ZN => N390);
   U383 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_13_port, A2 => 
                           net31074, ZN => N391);
   U384 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_14_port, A2 => 
                           net31074, ZN => N392);
   U385 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_15_port, A2 => 
                           net31074, ZN => N393);
   U386 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_16_port, A2 => 
                           net31074, ZN => N394);
   U387 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_17_port, A2 => 
                           net31074, ZN => N395);
   U388 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_18_port, A2 => 
                           net31074, ZN => N396);
   U389 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_19_port, A2 => 
                           net31074, ZN => N397);
   U390 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_20_port, A2 => 
                           net31072, ZN => N398);
   U391 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_21_port, A2 => 
                           net31072, ZN => N399);
   U392 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_22_port, A2 => 
                           net31072, ZN => N400);
   U393 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_23_port, A2 => 
                           net31072, ZN => N401);
   U394 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_24_port, A2 => 
                           net31072, ZN => N402);
   U395 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_25_port, A2 => 
                           net31072, ZN => N403);
   U396 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_26_port, A2 => 
                           net31072, ZN => N404);
   U397 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_27_port, A2 => 
                           net31072, ZN => N405);
   U398 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_28_port, A2 => 
                           net31072, ZN => N406);
   U399 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_29_port, A2 => 
                           net31070, ZN => N407);
   U400 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_30_port, A2 => 
                           net31070, ZN => N408);
   U401 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_31_port, A2 => 
                           net31070, ZN => N409);
   U402 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_0_port, A2 => net31080, ZN => 
                           N178);
   U403 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_1_port, A2 => net31080, ZN => 
                           N179);
   U404 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_2_port, A2 => net31080, ZN => 
                           N180);
   U405 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_3_port, A2 => net31080, ZN => 
                           N181);
   U406 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_4_port, A2 => net31080, ZN => 
                           N182);
   U407 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_5_port, A2 => net31078, ZN => 
                           N183);
   U408 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_6_port, A2 => net31078, ZN => 
                           N184);
   U409 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_7_port, A2 => net31078, ZN => 
                           N185);
   U410 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_8_port, A2 => net31078, ZN => 
                           N186);
   U411 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_9_port, A2 => net31078, ZN => 
                           N187);
   U412 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_10_port, A2 => net31078, ZN =>
                           N188);
   U413 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_11_port, A2 => net31078, ZN =>
                           N189);
   U414 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_12_port, A2 => net31078, ZN =>
                           N190);
   U415 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_13_port, A2 => net31078, ZN =>
                           N191);
   U416 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_14_port, A2 => net31078, ZN =>
                           N192);
   U417 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_15_port, A2 => net31086, ZN =>
                           N193);
   U418 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_16_port, A2 => RST, ZN => N194
                           );
   U419 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_17_port, A2 => RST, ZN => N195
                           );
   U420 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_18_port, A2 => RST, ZN => N196
                           );
   U421 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_19_port, A2 => RST, ZN => N197
                           );
   U422 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_20_port, A2 => RST, ZN => N198
                           );
   U423 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_21_port, A2 => RST, ZN => N199
                           );
   U424 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_22_port, A2 => RST, ZN => N200
                           );
   U425 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_23_port, A2 => RST, ZN => N201
                           );
   U426 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_24_port, A2 => RST, ZN => N202
                           );
   U427 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_25_port, A2 => RST, ZN => N203
                           );
   U428 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_26_port, A2 => RST, ZN => N204
                           );
   U429 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_27_port, A2 => RST, ZN => N205
                           );
   U430 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_28_port, A2 => RST, ZN => N206
                           );
   U431 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_29_port, A2 => RST, ZN => N207
                           );
   U432 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_30_port, A2 => RST, ZN => N208
                           );
   U433 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_31_port, A2 => net31066, ZN =>
                           N209);
   U434 : AND2_X1 port map( A1 => IR_OUT_11_port, A2 => net31068, ZN => N45);
   U435 : AND2_X1 port map( A1 => IR_OUT_12_port, A2 => net31068, ZN => N46);
   U436 : AND2_X1 port map( A1 => IR_OUT_13_port, A2 => net31068, ZN => N47);
   U437 : AND2_X1 port map( A1 => IR_OUT_14_port, A2 => net31068, ZN => N48);
   U438 : AND2_X1 port map( A1 => IR_OUT_15_port, A2 => net31068, ZN => N49);
   U439 : AND2_X1 port map( A1 => IR_OUT_16_port, A2 => net31068, ZN => N50);
   U440 : AND2_X1 port map( A1 => IR_OUT_17_port, A2 => net31068, ZN => N51);
   U441 : AND2_X1 port map( A1 => IR_OUT_18_port, A2 => net31068, ZN => N52);
   U442 : AND2_X1 port map( A1 => IR_OUT_19_port, A2 => net31066, ZN => N53);
   U443 : AND2_X1 port map( A1 => IR_OUT_20_port, A2 => net31066, ZN => N54);
   U444 : AND2_X1 port map( A1 => IR_OUT_21_port, A2 => net31066, ZN => N55);
   U445 : AND2_X1 port map( A1 => IR_OUT_22_port, A2 => net31066, ZN => N56);
   U446 : AND2_X1 port map( A1 => IR_OUT_23_port, A2 => net31066, ZN => N57);
   U447 : AND2_X1 port map( A1 => IR_OUT_24_port, A2 => net31066, ZN => N58);
   U448 : AND2_X1 port map( A1 => IR_OUT_25_port, A2 => net31066, ZN => N59);
   U449 : AND2_X1 port map( A1 => RF_WE, A2 => net31068, ZN => N98);
   U450 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_4_port, A2 => RST, ZN => N113);
   U451 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_4_port, A2 => net31088, ZN => 
                           N108);
   U452 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_1_port, A2 => net31088, ZN => 
                           N105);
   U453 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_0_port, A2 => net31088, ZN => 
                           N104);
   U454 : CLKBUF_X1 port map( A => ID_EX_RS2_NEXT_0_port, Z => n11_port);
   U455 : CLKBUF_X1 port map( A => ID_EX_RS2_NEXT_1_port, Z => n12_port);
   U456 : CLKBUF_X1 port map( A => ID_EX_RS2_NEXT_4_port, Z => n13_port);
   U457 : INV_X1 port map( A => n14_port, ZN => n15_port);
   U458 : INV_X1 port map( A => n16_port, ZN => n17_port);

end SYN_DLX_DATAPATH_ARCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18 is

   port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, PC_LATCH_EN, NPC_LATCH_EN, RF_WE, RegA_LATCH_EN, 
         RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
         EQ_COND : out std_logic;  ALU_OPCODE : out std_logic_vector (0 to 6); 
         DRAM_RE, DRAM_WE, LMD_LATCH_EN, JUMP_EN, JUMP_COND, WB_MUX_SEL, 
         JAL_MUX_SEL : out std_logic);

end DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18;

architecture SYN_DLX_CU_HW of 
   DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal aluOpcode1_6_port, aluOpcode1_5_port, aluOpcode1_4_port, 
      aluOpcode1_3_port, aluOpcode1_2_port, aluOpcode1_1_port, 
      aluOpcode1_0_port, aluOpcode2_6_port, aluOpcode2_5_port, 
      aluOpcode2_4_port, aluOpcode2_3_port, aluOpcode2_2_port, 
      aluOpcode2_1_port, aluOpcode2_0_port, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88
      , n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102
      , n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, IR_LATCH_EN_port, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729 : std_logic;

begin
   IR_LATCH_EN <= IR_LATCH_EN_port;
   PC_LATCH_EN <= IR_LATCH_EN_port;
   NPC_LATCH_EN <= IR_LATCH_EN_port;
   
   aluOpcode2_reg_6_inst : DFFS_X1 port map( D => aluOpcode1_6_port, CK => CLK,
                           SN => RST, Q => aluOpcode2_6_port, QN => n_1716);
   aluOpcode2_reg_5_inst : DFFS_X1 port map( D => aluOpcode1_5_port, CK => CLK,
                           SN => RST, Q => aluOpcode2_5_port, QN => n_1717);
   aluOpcode2_reg_4_inst : DFFR_X1 port map( D => aluOpcode1_4_port, CK => CLK,
                           RN => RST, Q => aluOpcode2_4_port, QN => n_1718);
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => aluOpcode1_3_port, CK => CLK,
                           RN => RST, Q => aluOpcode2_3_port, QN => n_1719);
   aluOpcode2_reg_2_inst : DFFS_X1 port map( D => aluOpcode1_2_port, CK => CLK,
                           SN => RST, Q => aluOpcode2_2_port, QN => n_1720);
   aluOpcode2_reg_1_inst : DFFS_X1 port map( D => aluOpcode1_1_port, CK => CLK,
                           SN => RST, Q => aluOpcode2_1_port, QN => n_1721);
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => aluOpcode1_0_port, CK => CLK,
                           RN => RST, Q => aluOpcode2_0_port, QN => n_1722);
   aluOpcode3_reg_6_inst : DFFS_X1 port map( D => aluOpcode2_6_port, CK => CLK,
                           SN => RST, Q => ALU_OPCODE(0), QN => n_1723);
   aluOpcode3_reg_5_inst : DFFS_X1 port map( D => aluOpcode2_5_port, CK => CLK,
                           SN => RST, Q => ALU_OPCODE(1), QN => n_1724);
   aluOpcode3_reg_4_inst : DFFR_X1 port map( D => aluOpcode2_4_port, CK => CLK,
                           RN => RST, Q => ALU_OPCODE(2), QN => n_1725);
   aluOpcode3_reg_3_inst : DFFR_X1 port map( D => aluOpcode2_3_port, CK => CLK,
                           RN => RST, Q => ALU_OPCODE(3), QN => n_1726);
   aluOpcode3_reg_2_inst : DFFS_X1 port map( D => aluOpcode2_2_port, CK => CLK,
                           SN => RST, Q => ALU_OPCODE(4), QN => n_1727);
   aluOpcode3_reg_1_inst : DFFS_X1 port map( D => aluOpcode2_1_port, CK => CLK,
                           SN => RST, Q => ALU_OPCODE(5), QN => n_1728);
   aluOpcode3_reg_0_inst : DFFR_X1 port map( D => aluOpcode2_0_port, CK => CLK,
                           RN => RST, Q => ALU_OPCODE(6), QN => n_1729);
   JAL_MUX_SEL <= '0';
   WB_MUX_SEL <= '0';
   JUMP_COND <= '0';
   JUMP_EN <= '0';
   LMD_LATCH_EN <= '0';
   DRAM_WE <= '0';
   DRAM_RE <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   RF_WE <= '0';
   U153 : NAND3_X1 port map( A1 => n52, A2 => n69, A3 => n30, ZN => n39);
   U154 : NAND3_X1 port map( A1 => n88, A2 => n89, A3 => n90, ZN => n40);
   U155 : NAND3_X1 port map( A1 => n91, A2 => n36, A3 => n92, ZN => n88);
   U156 : NAND3_X1 port map( A1 => n118, A2 => n119, A3 => n120, ZN => n117);
   U157 : NAND3_X1 port map( A1 => n112, A2 => IR_IN(26), A3 => n20, ZN => n67)
                           ;
   U158 : NAND3_X1 port map( A1 => n87, A2 => n86, A3 => n10, ZN => n116);
   U159 : NAND3_X1 port map( A1 => n27, A2 => IR_IN(2), A3 => n80, ZN => n87);
   U160 : NAND3_X1 port map( A1 => n112, A2 => n21, A3 => n20, ZN => n60);
   U161 : NAND3_X1 port map( A1 => n63, A2 => n21, A3 => n113, ZN => n123);
   U162 : NAND3_X1 port map( A1 => n92, A2 => n33, A3 => n27, ZN => n54);
   U163 : NAND3_X1 port map( A1 => IR_IN(1), A2 => n35, A3 => n91, ZN => n90);
   U164 : NAND3_X1 port map( A1 => IR_IN(2), A2 => n139, A3 => n142, ZN => n98)
                           ;
   U165 : NAND3_X1 port map( A1 => n37, A2 => n33, A3 => n79, ZN => n77);
   U166 : NAND3_X1 port map( A1 => n126, A2 => n68, A3 => n103, ZN => n134);
   U167 : NAND3_X1 port map( A1 => n63, A2 => n21, A3 => n66, ZN => n126);
   IR_LATCH_EN_port <= '0';
   U18 : NOR4_X1 port map( A1 => n12, A2 => n9, A3 => n65, A4 => n3, ZN => n111
                           );
   U19 : OAI221_X1 port map( B1 => n12, B2 => n8, C1 => n38, C2 => n39, A => 
                           RST, ZN => aluOpcode1_6_port);
   U20 : NAND4_X1 port map( A1 => n53, A2 => n25, A3 => n23, A4 => n54, ZN => 
                           n38);
   U21 : INV_X1 port map( A => n123, ZN => n12);
   U22 : OAI211_X1 port map( C1 => n40, C2 => n38, A => n41, B => RST, ZN => 
                           aluOpcode1_5_port);
   U23 : NAND4_X1 port map( A1 => n42, A2 => n13, A3 => n43, A4 => n44, ZN => 
                           n41);
   U24 : NOR4_X1 port map( A1 => n12, A2 => n3, A3 => n4, A4 => n45, ZN => n44)
                           ;
   U25 : INV_X1 port map( A => n60, ZN => n4);
   U26 : INV_X1 port map( A => n71, ZN => n27);
   U27 : NAND4_X1 port map( A1 => n25, A2 => n23, A3 => n30, A4 => n69, ZN => 
                           n61);
   U28 : INV_X1 port map( A => n40, ZN => n30);
   U29 : NAND2_X1 port map( A1 => n42, A2 => n51, ZN => n62);
   U30 : INV_X1 port map( A => n51, ZN => n8);
   U31 : INV_X1 port map( A => n57, ZN => n3);
   U32 : INV_X1 port map( A => n47, ZN => n15);
   U33 : INV_X1 port map( A => n114, ZN => n9);
   U34 : INV_X1 port map( A => n127, ZN => n7);
   U35 : INV_X1 port map( A => n77, ZN => n24);
   U36 : AOI211_X1 port map( C1 => n63, C2 => n64, A => n9, B => n65, ZN => n51
                           );
   U37 : AOI211_X1 port map( C1 => n63, C2 => n66, A => n2, B => n5, ZN => n42)
                           ;
   U38 : INV_X1 port map( A => n68, ZN => n2);
   U39 : INV_X1 port map( A => n67, ZN => n5);
   U40 : AOI211_X1 port map( C1 => n104, C2 => n66, A => n105, B => n106, ZN =>
                           n49);
   U41 : AOI211_X1 port map( C1 => n101, C2 => n102, A => n7, B => n6, ZN => 
                           n100);
   U42 : INV_X1 port map( A => n103, ZN => n6);
   U43 : NOR4_X1 port map( A1 => n121, A2 => n106, A3 => n15, A4 => n105, ZN =>
                           n120);
   U44 : NAND4_X1 port map( A1 => n48, A2 => n110, A3 => n109, A4 => n123, ZN 
                           => n121);
   U45 : NOR2_X1 port map( A1 => n21, A2 => n108, ZN => n104);
   U46 : AOI211_X1 port map( C1 => n124, C2 => n113, A => n45, B => n128, ZN =>
                           n118);
   U47 : OAI221_X1 port map( B1 => n81, B2 => n82, C1 => n83, C2 => n84, A => 
                           RST, ZN => aluOpcode1_2_port);
   U48 : OR2_X1 port map( A1 => n39, A2 => n74, ZN => n84);
   U49 : NAND4_X1 port map( A1 => n59, A2 => n58, A3 => n60, A4 => n111, ZN => 
                           n81);
   U50 : NAND4_X1 port map( A1 => n13, A2 => n99, A3 => n49, A4 => n100, ZN => 
                           n82);
   U51 : OAI211_X1 port map( C1 => n14, C2 => n129, A => n59, B => n58, ZN => 
                           n45);
   U52 : AOI21_X1 port map( B1 => n136, B2 => n137, A => n123, ZN => n135);
   U53 : AOI211_X1 port map( C1 => n34, C2 => n27, A => n138, B => n22, ZN => 
                           n137);
   U54 : NOR4_X1 port map( A1 => n24, A2 => n96, A3 => n140, A4 => n28, ZN => 
                           n136);
   U55 : INV_X1 port map( A => n73, ZN => n22);
   U56 : OAI211_X1 port map( C1 => n37, C2 => n90, A => n89, B => n54, ZN => 
                           n138);
   U57 : NAND2_X1 port map( A1 => n27, A2 => n35, ZN => n85);
   U58 : NAND2_X1 port map( A1 => n112, A2 => n122, ZN => n58);
   U59 : OAI211_X1 port map( C1 => n14, C2 => n21, A => n114, B => n58, ZN => 
                           n132);
   U60 : AND2_X1 port map( A1 => n133, A2 => n18, ZN => n112);
   U61 : OAI21_X1 port map( B1 => n85, B2 => n95, A => n75, ZN => n83);
   U62 : INV_X1 port map( A => n64, ZN => n14);
   U63 : NAND2_X1 port map( A1 => n34, A2 => n79, ZN => n73);
   U64 : NAND2_X1 port map( A1 => n112, A2 => n124, ZN => n59);
   U65 : NAND2_X1 port map( A1 => n141, A2 => n36, ZN => n71);
   U66 : NAND2_X1 port map( A1 => n122, A2 => n64, ZN => n109);
   U67 : AND2_X1 port map( A1 => n66, A2 => n102, ZN => n105);
   U68 : NAND2_X1 port map( A1 => n124, A2 => n64, ZN => n110);
   U69 : AOI21_X1 port map( B1 => n130, B2 => n131, A => n1, ZN => 
                           aluOpcode1_0_port);
   U70 : NOR4_X1 port map( A1 => n134, A2 => n135, A3 => n7, A4 => n128, ZN => 
                           n130);
   U71 : NOR4_X1 port map( A1 => n132, A2 => n105, A3 => n4, A4 => n15, ZN => 
                           n131);
   U72 : AOI21_X1 port map( B1 => n55, B2 => n56, A => n1, ZN => 
                           aluOpcode1_3_port);
   U73 : AND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           n56);
   U74 : AOI211_X1 port map( C1 => n53, C2 => n61, A => n62, B => n16, ZN => 
                           n55);
   U75 : INV_X1 port map( A => n48, ZN => n16);
   U76 : AOI21_X1 port map( B1 => n46, B2 => n43, A => n1, ZN => 
                           aluOpcode1_4_port);
   U77 : AOI21_X1 port map( B1 => n11, B2 => n50, A => n8, ZN => n46);
   U78 : INV_X1 port map( A => n38, ZN => n11);
   U79 : NAND2_X1 port map( A1 => n30, A2 => n52, ZN => n50);
   U80 : OAI211_X1 port map( C1 => n115, C2 => n116, A => n117, B => RST, ZN =>
                           aluOpcode1_1_port);
   U81 : NAND4_X1 port map( A1 => n76, A2 => n72, A3 => n73, A4 => n90, ZN => 
                           n115);
   U82 : NAND2_X1 port map( A1 => n104, A2 => n113, ZN => n114);
   U83 : NAND2_X1 port map( A1 => n79, A2 => n37, ZN => n72);
   U84 : AND3_X1 port map( A1 => n47, A2 => n48, A3 => n49, ZN => n43);
   U85 : NAND2_X1 port map( A1 => n93, A2 => n37, ZN => n69);
   U86 : INV_X1 port map( A => n74, ZN => n25);
   U87 : NAND2_X1 port map( A1 => n101, A2 => n124, ZN => n99);
   U88 : NAND2_X1 port map( A1 => n101, A2 => n122, ZN => n127);
   U89 : AND2_X1 port map( A1 => n122, A2 => n113, ZN => n128);
   U90 : AND2_X1 port map( A1 => n102, A2 => n113, ZN => n65);
   U91 : NAND2_X1 port map( A1 => n80, A2 => n26, ZN => n76);
   U92 : INV_X1 port map( A => n85, ZN => n26);
   U93 : NAND2_X1 port map( A1 => n112, A2 => n102, ZN => n57);
   U94 : INV_X1 port map( A => n95, ZN => n34);
   U95 : AND2_X1 port map( A1 => n66, A2 => n122, ZN => n106);
   U96 : NAND2_X1 port map( A1 => n125, A2 => n18, ZN => n47);
   U97 : NAND2_X1 port map( A1 => n66, A2 => n124, ZN => n68);
   U98 : NAND2_X1 port map( A1 => n101, A2 => n104, ZN => n103);
   U99 : AND4_X1 port map( A1 => n75, A2 => n76, A3 => n77, A4 => n78, ZN => 
                           n53);
   U100 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n78);
   U101 : INV_X1 port map( A => n86, ZN => n28);
   U102 : INV_X1 port map( A => n70, ZN => n23);
   U103 : OAI211_X1 port map( C1 => n33, C2 => n71, A => n72, B => n73, ZN => 
                           n70);
   U104 : INV_X1 port map( A => n107, ZN => n13);
   U105 : OAI211_X1 port map( C1 => n14, C2 => n108, A => n109, B => n110, ZN 
                           => n107);
   U106 : INV_X1 port map( A => n129, ZN => n20);
   U107 : INV_X1 port map( A => n97, ZN => n10);
   U108 : AND4_X1 port map( A1 => n126, A2 => n67, A3 => n127, A4 => n99, ZN =>
                           n119);
   U109 : NOR3_X1 port map( A1 => IR_IN(30), A2 => IR_IN(31), A3 => n18, ZN => 
                           n64);
   U110 : NOR3_X1 port map( A1 => IR_IN(30), A2 => IR_IN(31), A3 => IR_IN(29), 
                           ZN => n113);
   U111 : AOI211_X1 port map( C1 => IR_IN(1), C2 => n31, A => n96, B => n97, ZN
                           => n75);
   U112 : INV_X1 port map( A => n98, ZN => n31);
   U113 : NOR3_X1 port map( A1 => n29, A2 => IR_IN(4), A3 => n32, ZN => n141);
   U114 : INV_X1 port map( A => n139, ZN => n29);
   U115 : NOR3_X1 port map( A1 => IR_IN(6), A2 => IR_IN(10), A3 => n143, ZN => 
                           n139);
   U116 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN 
                           => n143);
   U117 : NOR3_X1 port map( A1 => IR_IN(0), A2 => IR_IN(3), A3 => n85, ZN => 
                           n96);
   U118 : NOR2_X1 port map( A1 => n108, A2 => IR_IN(26), ZN => n102);
   U119 : NOR3_X1 port map( A1 => IR_IN(3), A2 => IR_IN(5), A3 => IR_IN(4), ZN 
                           => n142);
   U120 : NOR2_X1 port map( A1 => IR_IN(28), A2 => IR_IN(27), ZN => n63);
   U121 : NOR3_X1 port map( A1 => n98, A2 => IR_IN(0), A3 => n36, ZN => n140);
   U122 : OAI21_X1 port map( B1 => IR_IN(0), B2 => n98, A => n12, ZN => n97);
   U123 : NOR2_X1 port map( A1 => n37, A2 => IR_IN(3), ZN => n80);
   U124 : NAND4_X1 port map( A1 => n141, A2 => n92, A3 => IR_IN(1), A4 => n33, 
                           ZN => n86);
   U125 : NAND4_X1 port map( A1 => n91, A2 => IR_IN(0), A3 => IR_IN(2), A4 => 
                           n36, ZN => n89);
   U126 : OAI211_X1 port map( C1 => IR_IN(0), C2 => n85, A => n86, B => n87, ZN
                           => n74);
   U127 : NOR2_X1 port map( A1 => n35, A2 => IR_IN(0), ZN => n92);
   U128 : AND3_X1 port map( A1 => n21, A2 => n19, A3 => IR_IN(27), ZN => n124);
   U129 : INV_X1 port map( A => IR_IN(0), ZN => n37);
   U130 : AND3_X1 port map( A1 => IR_IN(26), A2 => n19, A3 => IR_IN(27), ZN => 
                           n122);
   U131 : NAND2_X1 port map( A1 => IR_IN(0), A2 => IR_IN(3), ZN => n95);
   U132 : AND2_X1 port map( A1 => n133, A2 => IR_IN(29), ZN => n66);
   U133 : NAND2_X1 port map( A1 => IR_IN(0), A2 => n93, ZN => n52);
   U134 : AND3_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), A3 => IR_IN(31), 
                           ZN => n101);
   U135 : INV_X1 port map( A => IR_IN(26), ZN => n21);
   U136 : INV_X1 port map( A => IR_IN(1), ZN => n36);
   U137 : AND3_X1 port map( A1 => IR_IN(1), A2 => n35, A3 => n141, ZN => n79);
   U138 : INV_X1 port map( A => IR_IN(3), ZN => n33);
   U139 : INV_X1 port map( A => IR_IN(2), ZN => n35);
   U140 : NOR2_X1 port map( A1 => n17, A2 => IR_IN(31), ZN => n133);
   U141 : NAND2_X1 port map( A1 => n125, A2 => IR_IN(29), ZN => n48);
   U142 : INV_X1 port map( A => IR_IN(29), ZN => n18);
   U143 : NAND2_X1 port map( A1 => IR_IN(27), A2 => IR_IN(28), ZN => n129);
   U144 : OR2_X1 port map( A1 => n19, A2 => IR_IN(27), ZN => n108);
   U145 : AND3_X1 port map( A1 => n122, A2 => n17, A3 => IR_IN(31), ZN => n125)
                           ;
   U146 : AND3_X1 port map( A1 => IR_IN(3), A2 => n139, A3 => IR_IN(4), ZN => 
                           n94);
   U147 : INV_X1 port map( A => IR_IN(5), ZN => n32);
   U148 : AND2_X1 port map( A1 => IR_IN(5), A2 => n94, ZN => n91);
   U149 : AND4_X1 port map( A1 => IR_IN(2), A2 => IR_IN(1), A3 => n94, A4 => 
                           n32, ZN => n93);
   U150 : INV_X1 port map( A => IR_IN(28), ZN => n19);
   U151 : INV_X1 port map( A => IR_IN(30), ZN => n17);
   U152 : INV_X1 port map( A => RST, ZN => n1);

end SYN_DLX_CU_HW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( CLK, RST : in std_logic);

end DLX;

architecture SYN_DLX_RTL of DLX is

   component DLX_DRAM_N256_NW32
      port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector 
            (31 downto 0);  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component DLX_IRAM_RAM_DEPTH256_I_SIZE32
      port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  
            DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32
      port( CLK, RST : in std_logic;  IR_IN, DRAM_OUT : in std_logic_vector (31
            downto 0);  IR_LATCH_EN, PC_LATCH_EN, NPC_LATCH_EN, RF_WE, 
            RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, 
            ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
            std_logic_vector (0 to 6);  LMD_LATCH_EN, JUMP_EN, JUMP_COND, 
            WB_MUX_SEL, JAL_MUX_SEL : in std_logic;  IR_OUT, PC_OUT, ALU_OUT, 
            DRAM_IN : out std_logic_vector (31 downto 0));
   end component;
   
   component 
      DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18
      port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, PC_LATCH_EN, NPC_LATCH_EN, RF_WE, RegA_LATCH_EN, 
            RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
            EQ_COND : out std_logic;  ALU_OPCODE : out std_logic_vector (0 to 
            6);  DRAM_RE, DRAM_WE, LMD_LATCH_EN, JUMP_EN, JUMP_COND, WB_MUX_SEL
            , JAL_MUX_SEL : out std_logic);
   end component;
   
   signal IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, 
      IR_26_port, IR_25_port, IR_24_port, IR_23_port, IR_22_port, IR_21_port, 
      IR_20_port, IR_19_port, IR_18_port, IR_17_port, IR_16_port, IR_15_port, 
      IR_14_port, IR_13_port, IR_12_port, IR_11_port, IR_10_port, IR_9_port, 
      IR_8_port, IR_7_port, IR_6_port, IR_5_port, IR_4_port, IR_3_port, 
      IR_2_port, IR_1_port, IR_0_port, IR_LATCH_EN_i, PC_LATCH_EN_i, 
      NPC_LATCH_EN_i, RF_WE_i, RegA_LATCH_EN_i, RegB_LATCH_EN_i, 
      RegIMM_LATCH_EN_i, MUXA_SEL_i, MUXB_SEL_i, ALU_OUTREG_EN_i, EQ_COND_i, 
      ALU_OPCODE_i_0_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_4_port, ALU_OPCODE_i_5_port, 
      ALU_OPCODE_i_6_port, DRAM_RE_i, DRAM_WE_i, LMD_LATCH_EN_i, JUMP_EN_i, 
      JUMP_COND_i, WB_MUX_SEL_i, JAL_MUX_SEL_i, IR_BUS_31_port, IR_BUS_30_port,
      IR_BUS_29_port, IR_BUS_28_port, IR_BUS_27_port, IR_BUS_26_port, 
      IR_BUS_25_port, IR_BUS_24_port, IR_BUS_23_port, IR_BUS_22_port, 
      IR_BUS_21_port, IR_BUS_20_port, IR_BUS_19_port, IR_BUS_18_port, 
      IR_BUS_17_port, IR_BUS_16_port, IR_BUS_15_port, IR_BUS_14_port, 
      IR_BUS_13_port, IR_BUS_12_port, IR_BUS_11_port, IR_BUS_10_port, 
      IR_BUS_9_port, IR_BUS_8_port, IR_BUS_7_port, IR_BUS_6_port, IR_BUS_5_port
      , IR_BUS_4_port, IR_BUS_3_port, IR_BUS_2_port, IR_BUS_1_port, 
      IR_BUS_0_port, DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, PC_31_port, PC_30_port, PC_29_port, PC_28_port, 
      PC_27_port, PC_26_port, PC_25_port, PC_24_port, PC_23_port, PC_22_port, 
      PC_21_port, PC_20_port, PC_19_port, PC_18_port, PC_17_port, PC_16_port, 
      PC_15_port, PC_14_port, PC_13_port, PC_12_port, PC_11_port, PC_10_port, 
      PC_9_port, PC_8_port, PC_7_port, PC_6_port, PC_5_port, PC_4_port, 
      PC_3_port, PC_2_port, PC_1_port, PC_0_port, DATA_ADDR_31_port, 
      DATA_ADDR_30_port, DATA_ADDR_29_port, DATA_ADDR_28_port, 
      DATA_ADDR_27_port, DATA_ADDR_26_port, DATA_ADDR_25_port, 
      DATA_ADDR_24_port, DATA_ADDR_23_port, DATA_ADDR_22_port, 
      DATA_ADDR_21_port, DATA_ADDR_20_port, DATA_ADDR_19_port, 
      DATA_ADDR_18_port, DATA_ADDR_17_port, DATA_ADDR_16_port, 
      DATA_ADDR_15_port, DATA_ADDR_14_port, DATA_ADDR_13_port, 
      DATA_ADDR_12_port, DATA_ADDR_11_port, DATA_ADDR_10_port, DATA_ADDR_9_port
      , DATA_ADDR_8_port, DATA_ADDR_7_port, DATA_ADDR_6_port, DATA_ADDR_5_port,
      DATA_ADDR_4_port, DATA_ADDR_3_port, DATA_ADDR_2_port, DATA_ADDR_1_port, 
      DATA_ADDR_0_port, DATA_IN_31_port, DATA_IN_30_port, DATA_IN_29_port, 
      DATA_IN_28_port, DATA_IN_27_port, DATA_IN_26_port, DATA_IN_25_port, 
      DATA_IN_24_port, DATA_IN_23_port, DATA_IN_22_port, DATA_IN_21_port, 
      DATA_IN_20_port, DATA_IN_19_port, DATA_IN_18_port, DATA_IN_17_port, 
      DATA_IN_16_port, DATA_IN_15_port, DATA_IN_14_port, DATA_IN_13_port, 
      DATA_IN_12_port, DATA_IN_11_port, DATA_IN_10_port, DATA_IN_9_port, 
      DATA_IN_8_port, DATA_IN_7_port, DATA_IN_6_port, DATA_IN_5_port, 
      DATA_IN_4_port, DATA_IN_3_port, DATA_IN_2_port, DATA_IN_1_port, 
      DATA_IN_0_port, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, 
      n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, 
      n_1746, n_1747 : std_logic;

begin
   
   CU_I : DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18 
                           port map( CLK => CLK, RST => RST, IR_IN(31) => 
                           IR_31_port, IR_IN(30) => IR_30_port, IR_IN(29) => 
                           IR_29_port, IR_IN(28) => IR_28_port, IR_IN(27) => 
                           IR_27_port, IR_IN(26) => IR_26_port, IR_IN(25) => 
                           IR_25_port, IR_IN(24) => IR_24_port, IR_IN(23) => 
                           IR_23_port, IR_IN(22) => IR_22_port, IR_IN(21) => 
                           IR_21_port, IR_IN(20) => IR_20_port, IR_IN(19) => 
                           IR_19_port, IR_IN(18) => IR_18_port, IR_IN(17) => 
                           IR_17_port, IR_IN(16) => IR_16_port, IR_IN(15) => 
                           IR_15_port, IR_IN(14) => IR_14_port, IR_IN(13) => 
                           IR_13_port, IR_IN(12) => IR_12_port, IR_IN(11) => 
                           IR_11_port, IR_IN(10) => IR_10_port, IR_IN(9) => 
                           IR_9_port, IR_IN(8) => IR_8_port, IR_IN(7) => 
                           IR_7_port, IR_IN(6) => IR_6_port, IR_IN(5) => 
                           IR_5_port, IR_IN(4) => IR_4_port, IR_IN(3) => 
                           IR_3_port, IR_IN(2) => IR_2_port, IR_IN(1) => 
                           IR_1_port, IR_IN(0) => IR_0_port, IR_LATCH_EN => 
                           n_1730, PC_LATCH_EN => n_1731, NPC_LATCH_EN => 
                           n_1732, RF_WE => n_1733, RegA_LATCH_EN => n_1734, 
                           RegB_LATCH_EN => n_1735, RegIMM_LATCH_EN => n_1736, 
                           MUXA_SEL => n_1737, MUXB_SEL => n_1738, 
                           ALU_OUTREG_EN => n_1739, EQ_COND => n_1740, 
                           ALU_OPCODE(0) => ALU_OPCODE_i_0_port, ALU_OPCODE(1) 
                           => ALU_OPCODE_i_1_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_4_port, ALU_OPCODE(5) => 
                           ALU_OPCODE_i_5_port, ALU_OPCODE(6) => 
                           ALU_OPCODE_i_6_port, DRAM_RE => n_1741, DRAM_WE => 
                           n_1742, LMD_LATCH_EN => n_1743, JUMP_EN => n_1744, 
                           JUMP_COND => n_1745, WB_MUX_SEL => n_1746, 
                           JAL_MUX_SEL => n_1747);
   DATAPATH_I : 
                           DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32 
                           port map( CLK => CLK, RST => RST, IR_IN(31) => 
                           IR_BUS_31_port, IR_IN(30) => IR_BUS_30_port, 
                           IR_IN(29) => IR_BUS_29_port, IR_IN(28) => 
                           IR_BUS_28_port, IR_IN(27) => IR_BUS_27_port, 
                           IR_IN(26) => IR_BUS_26_port, IR_IN(25) => 
                           IR_BUS_25_port, IR_IN(24) => IR_BUS_24_port, 
                           IR_IN(23) => IR_BUS_23_port, IR_IN(22) => 
                           IR_BUS_22_port, IR_IN(21) => IR_BUS_21_port, 
                           IR_IN(20) => IR_BUS_20_port, IR_IN(19) => 
                           IR_BUS_19_port, IR_IN(18) => IR_BUS_18_port, 
                           IR_IN(17) => IR_BUS_17_port, IR_IN(16) => 
                           IR_BUS_16_port, IR_IN(15) => IR_BUS_15_port, 
                           IR_IN(14) => IR_BUS_14_port, IR_IN(13) => 
                           IR_BUS_13_port, IR_IN(12) => IR_BUS_12_port, 
                           IR_IN(11) => IR_BUS_11_port, IR_IN(10) => 
                           IR_BUS_10_port, IR_IN(9) => IR_BUS_9_port, IR_IN(8) 
                           => IR_BUS_8_port, IR_IN(7) => IR_BUS_7_port, 
                           IR_IN(6) => IR_BUS_6_port, IR_IN(5) => IR_BUS_5_port
                           , IR_IN(4) => IR_BUS_4_port, IR_IN(3) => 
                           IR_BUS_3_port, IR_IN(2) => IR_BUS_2_port, IR_IN(1) 
                           => IR_BUS_1_port, IR_IN(0) => IR_BUS_0_port, 
                           DRAM_OUT(31) => DATA_OUT_31_port, DRAM_OUT(30) => 
                           DATA_OUT_30_port, DRAM_OUT(29) => DATA_OUT_29_port, 
                           DRAM_OUT(28) => DATA_OUT_28_port, DRAM_OUT(27) => 
                           DATA_OUT_27_port, DRAM_OUT(26) => DATA_OUT_26_port, 
                           DRAM_OUT(25) => DATA_OUT_25_port, DRAM_OUT(24) => 
                           DATA_OUT_24_port, DRAM_OUT(23) => DATA_OUT_23_port, 
                           DRAM_OUT(22) => DATA_OUT_22_port, DRAM_OUT(21) => 
                           DATA_OUT_21_port, DRAM_OUT(20) => DATA_OUT_20_port, 
                           DRAM_OUT(19) => DATA_OUT_19_port, DRAM_OUT(18) => 
                           DATA_OUT_18_port, DRAM_OUT(17) => DATA_OUT_17_port, 
                           DRAM_OUT(16) => DATA_OUT_16_port, DRAM_OUT(15) => 
                           DATA_OUT_15_port, DRAM_OUT(14) => DATA_OUT_14_port, 
                           DRAM_OUT(13) => DATA_OUT_13_port, DRAM_OUT(12) => 
                           DATA_OUT_12_port, DRAM_OUT(11) => DATA_OUT_11_port, 
                           DRAM_OUT(10) => DATA_OUT_10_port, DRAM_OUT(9) => 
                           DATA_OUT_9_port, DRAM_OUT(8) => DATA_OUT_8_port, 
                           DRAM_OUT(7) => DATA_OUT_7_port, DRAM_OUT(6) => 
                           DATA_OUT_6_port, DRAM_OUT(5) => DATA_OUT_5_port, 
                           DRAM_OUT(4) => DATA_OUT_4_port, DRAM_OUT(3) => 
                           DATA_OUT_3_port, DRAM_OUT(2) => DATA_OUT_2_port, 
                           DRAM_OUT(1) => DATA_OUT_1_port, DRAM_OUT(0) => 
                           DATA_OUT_0_port, IR_LATCH_EN => IR_LATCH_EN_i, 
                           PC_LATCH_EN => PC_LATCH_EN_i, NPC_LATCH_EN => 
                           NPC_LATCH_EN_i, RF_WE => RF_WE_i, RegA_LATCH_EN => 
                           RegA_LATCH_EN_i, RegB_LATCH_EN => RegB_LATCH_EN_i, 
                           RegIMM_LATCH_EN => RegIMM_LATCH_EN_i, MUXA_SEL => 
                           MUXA_SEL_i, MUXB_SEL => MUXB_SEL_i, ALU_OUTREG_EN =>
                           ALU_OUTREG_EN_i, EQ_COND => EQ_COND_i, ALU_OPCODE(0)
                           => ALU_OPCODE_i_0_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_4_port, ALU_OPCODE(5) => 
                           ALU_OPCODE_i_5_port, ALU_OPCODE(6) => 
                           ALU_OPCODE_i_6_port, LMD_LATCH_EN => LMD_LATCH_EN_i,
                           JUMP_EN => JUMP_EN_i, JUMP_COND => JUMP_COND_i, 
                           WB_MUX_SEL => WB_MUX_SEL_i, JAL_MUX_SEL => 
                           JAL_MUX_SEL_i, IR_OUT(31) => IR_31_port, IR_OUT(30) 
                           => IR_30_port, IR_OUT(29) => IR_29_port, IR_OUT(28) 
                           => IR_28_port, IR_OUT(27) => IR_27_port, IR_OUT(26) 
                           => IR_26_port, IR_OUT(25) => IR_25_port, IR_OUT(24) 
                           => IR_24_port, IR_OUT(23) => IR_23_port, IR_OUT(22) 
                           => IR_22_port, IR_OUT(21) => IR_21_port, IR_OUT(20) 
                           => IR_20_port, IR_OUT(19) => IR_19_port, IR_OUT(18) 
                           => IR_18_port, IR_OUT(17) => IR_17_port, IR_OUT(16) 
                           => IR_16_port, IR_OUT(15) => IR_15_port, IR_OUT(14) 
                           => IR_14_port, IR_OUT(13) => IR_13_port, IR_OUT(12) 
                           => IR_12_port, IR_OUT(11) => IR_11_port, IR_OUT(10) 
                           => IR_10_port, IR_OUT(9) => IR_9_port, IR_OUT(8) => 
                           IR_8_port, IR_OUT(7) => IR_7_port, IR_OUT(6) => 
                           IR_6_port, IR_OUT(5) => IR_5_port, IR_OUT(4) => 
                           IR_4_port, IR_OUT(3) => IR_3_port, IR_OUT(2) => 
                           IR_2_port, IR_OUT(1) => IR_1_port, IR_OUT(0) => 
                           IR_0_port, PC_OUT(31) => PC_31_port, PC_OUT(30) => 
                           PC_30_port, PC_OUT(29) => PC_29_port, PC_OUT(28) => 
                           PC_28_port, PC_OUT(27) => PC_27_port, PC_OUT(26) => 
                           PC_26_port, PC_OUT(25) => PC_25_port, PC_OUT(24) => 
                           PC_24_port, PC_OUT(23) => PC_23_port, PC_OUT(22) => 
                           PC_22_port, PC_OUT(21) => PC_21_port, PC_OUT(20) => 
                           PC_20_port, PC_OUT(19) => PC_19_port, PC_OUT(18) => 
                           PC_18_port, PC_OUT(17) => PC_17_port, PC_OUT(16) => 
                           PC_16_port, PC_OUT(15) => PC_15_port, PC_OUT(14) => 
                           PC_14_port, PC_OUT(13) => PC_13_port, PC_OUT(12) => 
                           PC_12_port, PC_OUT(11) => PC_11_port, PC_OUT(10) => 
                           PC_10_port, PC_OUT(9) => PC_9_port, PC_OUT(8) => 
                           PC_8_port, PC_OUT(7) => PC_7_port, PC_OUT(6) => 
                           PC_6_port, PC_OUT(5) => PC_5_port, PC_OUT(4) => 
                           PC_4_port, PC_OUT(3) => PC_3_port, PC_OUT(2) => 
                           PC_2_port, PC_OUT(1) => PC_1_port, PC_OUT(0) => 
                           PC_0_port, ALU_OUT(31) => DATA_ADDR_31_port, 
                           ALU_OUT(30) => DATA_ADDR_30_port, ALU_OUT(29) => 
                           DATA_ADDR_29_port, ALU_OUT(28) => DATA_ADDR_28_port,
                           ALU_OUT(27) => DATA_ADDR_27_port, ALU_OUT(26) => 
                           DATA_ADDR_26_port, ALU_OUT(25) => DATA_ADDR_25_port,
                           ALU_OUT(24) => DATA_ADDR_24_port, ALU_OUT(23) => 
                           DATA_ADDR_23_port, ALU_OUT(22) => DATA_ADDR_22_port,
                           ALU_OUT(21) => DATA_ADDR_21_port, ALU_OUT(20) => 
                           DATA_ADDR_20_port, ALU_OUT(19) => DATA_ADDR_19_port,
                           ALU_OUT(18) => DATA_ADDR_18_port, ALU_OUT(17) => 
                           DATA_ADDR_17_port, ALU_OUT(16) => DATA_ADDR_16_port,
                           ALU_OUT(15) => DATA_ADDR_15_port, ALU_OUT(14) => 
                           DATA_ADDR_14_port, ALU_OUT(13) => DATA_ADDR_13_port,
                           ALU_OUT(12) => DATA_ADDR_12_port, ALU_OUT(11) => 
                           DATA_ADDR_11_port, ALU_OUT(10) => DATA_ADDR_10_port,
                           ALU_OUT(9) => DATA_ADDR_9_port, ALU_OUT(8) => 
                           DATA_ADDR_8_port, ALU_OUT(7) => DATA_ADDR_7_port, 
                           ALU_OUT(6) => DATA_ADDR_6_port, ALU_OUT(5) => 
                           DATA_ADDR_5_port, ALU_OUT(4) => DATA_ADDR_4_port, 
                           ALU_OUT(3) => DATA_ADDR_3_port, ALU_OUT(2) => 
                           DATA_ADDR_2_port, ALU_OUT(1) => DATA_ADDR_1_port, 
                           ALU_OUT(0) => DATA_ADDR_0_port, DRAM_IN(31) => 
                           DATA_IN_31_port, DRAM_IN(30) => DATA_IN_30_port, 
                           DRAM_IN(29) => DATA_IN_29_port, DRAM_IN(28) => 
                           DATA_IN_28_port, DRAM_IN(27) => DATA_IN_27_port, 
                           DRAM_IN(26) => DATA_IN_26_port, DRAM_IN(25) => 
                           DATA_IN_25_port, DRAM_IN(24) => DATA_IN_24_port, 
                           DRAM_IN(23) => DATA_IN_23_port, DRAM_IN(22) => 
                           DATA_IN_22_port, DRAM_IN(21) => DATA_IN_21_port, 
                           DRAM_IN(20) => DATA_IN_20_port, DRAM_IN(19) => 
                           DATA_IN_19_port, DRAM_IN(18) => DATA_IN_18_port, 
                           DRAM_IN(17) => DATA_IN_17_port, DRAM_IN(16) => 
                           DATA_IN_16_port, DRAM_IN(15) => DATA_IN_15_port, 
                           DRAM_IN(14) => DATA_IN_14_port, DRAM_IN(13) => 
                           DATA_IN_13_port, DRAM_IN(12) => DATA_IN_12_port, 
                           DRAM_IN(11) => DATA_IN_11_port, DRAM_IN(10) => 
                           DATA_IN_10_port, DRAM_IN(9) => DATA_IN_9_port, 
                           DRAM_IN(8) => DATA_IN_8_port, DRAM_IN(7) => 
                           DATA_IN_7_port, DRAM_IN(6) => DATA_IN_6_port, 
                           DRAM_IN(5) => DATA_IN_5_port, DRAM_IN(4) => 
                           DATA_IN_4_port, DRAM_IN(3) => DATA_IN_3_port, 
                           DRAM_IN(2) => DATA_IN_2_port, DRAM_IN(1) => 
                           DATA_IN_1_port, DRAM_IN(0) => DATA_IN_0_port);
   IRAM_I : DLX_IRAM_RAM_DEPTH256_I_SIZE32 port map( RST => RST, ADDR(31) => 
                           PC_31_port, ADDR(30) => PC_30_port, ADDR(29) => 
                           PC_29_port, ADDR(28) => PC_28_port, ADDR(27) => 
                           PC_27_port, ADDR(26) => PC_26_port, ADDR(25) => 
                           PC_25_port, ADDR(24) => PC_24_port, ADDR(23) => 
                           PC_23_port, ADDR(22) => PC_22_port, ADDR(21) => 
                           PC_21_port, ADDR(20) => PC_20_port, ADDR(19) => 
                           PC_19_port, ADDR(18) => PC_18_port, ADDR(17) => 
                           PC_17_port, ADDR(16) => PC_16_port, ADDR(15) => 
                           PC_15_port, ADDR(14) => PC_14_port, ADDR(13) => 
                           PC_13_port, ADDR(12) => PC_12_port, ADDR(11) => 
                           PC_11_port, ADDR(10) => PC_10_port, ADDR(9) => 
                           PC_9_port, ADDR(8) => PC_8_port, ADDR(7) => 
                           PC_7_port, ADDR(6) => PC_6_port, ADDR(5) => 
                           PC_5_port, ADDR(4) => PC_4_port, ADDR(3) => 
                           PC_3_port, ADDR(2) => PC_2_port, ADDR(1) => 
                           PC_1_port, ADDR(0) => PC_0_port, DOUT(31) => 
                           IR_BUS_31_port, DOUT(30) => IR_BUS_30_port, DOUT(29)
                           => IR_BUS_29_port, DOUT(28) => IR_BUS_28_port, 
                           DOUT(27) => IR_BUS_27_port, DOUT(26) => 
                           IR_BUS_26_port, DOUT(25) => IR_BUS_25_port, DOUT(24)
                           => IR_BUS_24_port, DOUT(23) => IR_BUS_23_port, 
                           DOUT(22) => IR_BUS_22_port, DOUT(21) => 
                           IR_BUS_21_port, DOUT(20) => IR_BUS_20_port, DOUT(19)
                           => IR_BUS_19_port, DOUT(18) => IR_BUS_18_port, 
                           DOUT(17) => IR_BUS_17_port, DOUT(16) => 
                           IR_BUS_16_port, DOUT(15) => IR_BUS_15_port, DOUT(14)
                           => IR_BUS_14_port, DOUT(13) => IR_BUS_13_port, 
                           DOUT(12) => IR_BUS_12_port, DOUT(11) => 
                           IR_BUS_11_port, DOUT(10) => IR_BUS_10_port, DOUT(9) 
                           => IR_BUS_9_port, DOUT(8) => IR_BUS_8_port, DOUT(7) 
                           => IR_BUS_7_port, DOUT(6) => IR_BUS_6_port, DOUT(5) 
                           => IR_BUS_5_port, DOUT(4) => IR_BUS_4_port, DOUT(3) 
                           => IR_BUS_3_port, DOUT(2) => IR_BUS_2_port, DOUT(1) 
                           => IR_BUS_1_port, DOUT(0) => IR_BUS_0_port);
   DRAM_I : DLX_DRAM_N256_NW32 port map( CLK => CLK, RST => RST, RE => 
                           DRAM_RE_i, WE => DRAM_WE_i, ADDR(31) => 
                           DATA_ADDR_31_port, ADDR(30) => DATA_ADDR_30_port, 
                           ADDR(29) => DATA_ADDR_29_port, ADDR(28) => 
                           DATA_ADDR_28_port, ADDR(27) => DATA_ADDR_27_port, 
                           ADDR(26) => DATA_ADDR_26_port, ADDR(25) => 
                           DATA_ADDR_25_port, ADDR(24) => DATA_ADDR_24_port, 
                           ADDR(23) => DATA_ADDR_23_port, ADDR(22) => 
                           DATA_ADDR_22_port, ADDR(21) => DATA_ADDR_21_port, 
                           ADDR(20) => DATA_ADDR_20_port, ADDR(19) => 
                           DATA_ADDR_19_port, ADDR(18) => DATA_ADDR_18_port, 
                           ADDR(17) => DATA_ADDR_17_port, ADDR(16) => 
                           DATA_ADDR_16_port, ADDR(15) => DATA_ADDR_15_port, 
                           ADDR(14) => DATA_ADDR_14_port, ADDR(13) => 
                           DATA_ADDR_13_port, ADDR(12) => DATA_ADDR_12_port, 
                           ADDR(11) => DATA_ADDR_11_port, ADDR(10) => 
                           DATA_ADDR_10_port, ADDR(9) => DATA_ADDR_9_port, 
                           ADDR(8) => DATA_ADDR_8_port, ADDR(7) => 
                           DATA_ADDR_7_port, ADDR(6) => DATA_ADDR_6_port, 
                           ADDR(5) => DATA_ADDR_5_port, ADDR(4) => 
                           DATA_ADDR_4_port, ADDR(3) => DATA_ADDR_3_port, 
                           ADDR(2) => DATA_ADDR_2_port, ADDR(1) => 
                           DATA_ADDR_1_port, ADDR(0) => DATA_ADDR_0_port, 
                           DIN(31) => DATA_IN_31_port, DIN(30) => 
                           DATA_IN_30_port, DIN(29) => DATA_IN_29_port, DIN(28)
                           => DATA_IN_28_port, DIN(27) => DATA_IN_27_port, 
                           DIN(26) => DATA_IN_26_port, DIN(25) => 
                           DATA_IN_25_port, DIN(24) => DATA_IN_24_port, DIN(23)
                           => DATA_IN_23_port, DIN(22) => DATA_IN_22_port, 
                           DIN(21) => DATA_IN_21_port, DIN(20) => 
                           DATA_IN_20_port, DIN(19) => DATA_IN_19_port, DIN(18)
                           => DATA_IN_18_port, DIN(17) => DATA_IN_17_port, 
                           DIN(16) => DATA_IN_16_port, DIN(15) => 
                           DATA_IN_15_port, DIN(14) => DATA_IN_14_port, DIN(13)
                           => DATA_IN_13_port, DIN(12) => DATA_IN_12_port, 
                           DIN(11) => DATA_IN_11_port, DIN(10) => 
                           DATA_IN_10_port, DIN(9) => DATA_IN_9_port, DIN(8) =>
                           DATA_IN_8_port, DIN(7) => DATA_IN_7_port, DIN(6) => 
                           DATA_IN_6_port, DIN(5) => DATA_IN_5_port, DIN(4) => 
                           DATA_IN_4_port, DIN(3) => DATA_IN_3_port, DIN(2) => 
                           DATA_IN_2_port, DIN(1) => DATA_IN_1_port, DIN(0) => 
                           DATA_IN_0_port, DOUT(31) => DATA_OUT_31_port, 
                           DOUT(30) => DATA_OUT_30_port, DOUT(29) => 
                           DATA_OUT_29_port, DOUT(28) => DATA_OUT_28_port, 
                           DOUT(27) => DATA_OUT_27_port, DOUT(26) => 
                           DATA_OUT_26_port, DOUT(25) => DATA_OUT_25_port, 
                           DOUT(24) => DATA_OUT_24_port, DOUT(23) => 
                           DATA_OUT_23_port, DOUT(22) => DATA_OUT_22_port, 
                           DOUT(21) => DATA_OUT_21_port, DOUT(20) => 
                           DATA_OUT_20_port, DOUT(19) => DATA_OUT_19_port, 
                           DOUT(18) => DATA_OUT_18_port, DOUT(17) => 
                           DATA_OUT_17_port, DOUT(16) => DATA_OUT_16_port, 
                           DOUT(15) => DATA_OUT_15_port, DOUT(14) => 
                           DATA_OUT_14_port, DOUT(13) => DATA_OUT_13_port, 
                           DOUT(12) => DATA_OUT_12_port, DOUT(11) => 
                           DATA_OUT_11_port, DOUT(10) => DATA_OUT_10_port, 
                           DOUT(9) => DATA_OUT_9_port, DOUT(8) => 
                           DATA_OUT_8_port, DOUT(7) => DATA_OUT_7_port, DOUT(6)
                           => DATA_OUT_6_port, DOUT(5) => DATA_OUT_5_port, 
                           DOUT(4) => DATA_OUT_4_port, DOUT(3) => 
                           DATA_OUT_3_port, DOUT(2) => DATA_OUT_2_port, DOUT(1)
                           => DATA_OUT_1_port, DOUT(0) => DATA_OUT_0_port);
   JAL_MUX_SEL_i <= '0';
   WB_MUX_SEL_i <= '0';
   JUMP_COND_i <= '0';
   JUMP_EN_i <= '0';
   LMD_LATCH_EN_i <= '0';
   DRAM_WE_i <= '0';
   DRAM_RE_i <= '0';
   EQ_COND_i <= '0';
   ALU_OUTREG_EN_i <= '0';
   MUXB_SEL_i <= '0';
   MUXA_SEL_i <= '0';
   RegIMM_LATCH_EN_i <= '0';
   RegB_LATCH_EN_i <= '0';
   RegA_LATCH_EN_i <= '0';
   RF_WE_i <= '0';
   NPC_LATCH_EN_i <= '0';
   PC_LATCH_EN_i <= '0';
   IR_LATCH_EN_i <= '0';

end SYN_DLX_RTL;

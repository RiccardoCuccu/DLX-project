
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (OP_SLL, OP_SRL, OP_SRA, OP_ADD, OP_ADDU, OP_SUB, OP_SUBU, 
   OP_AND, OP_OR, OP_XOR, OP_SEQ, OP_SNE, OP_SLT, OP_SGT, OP_SLE, OP_SGE, 
   OP_MOVI2S, OP_MOVS2I, OP_MOVF, OP_MOVD, OP_MOVFP2I, OP_MOVI2FP, OP_MOVI2T, 
   OP_MOVT2I, OP_SLTU, OP_SGTU, OP_SLEU, OP_SGEU, OP_ADDF, OP_SUBF, OP_MULTF, 
   OP_DIVF, OP_ADDD, OP_SUBD, OP_MULTD, OP_DIVD, OP_CVTF2D, OP_CVTF2I, 
   OP_CVTD2F, OP_CVTD2I, OP_CVTI2F, OP_CVTI2D, OP_MULT, OP_DIV, OP_EQF, OP_NEF,
   OP_LTF, OP_GTF, OP_LEF, OP_GEF, OP_MULTU, OP_DIVU, OP_EQD, OP_NED, OP_LTD, 
   OP_GTD, OP_LED, OP_GED, OP_BEQZ, OP_BNEZ, OP_BFPT, OP_BFPF, OP_ADDI, 
   OP_ADDUI, OP_SUBI, OP_SUBUI, OP_ANDI, OP_ORI, OP_XORI, OP_LHI, OP_RFE, 
   OP_TRAP, OP_JR, OP_JALR, OP_SLLI, OP_SRLI, OP_SRAI, OP_SEQI, OP_SNEI, 
   OP_SLTI, OP_SGTI, OP_SLEI, OP_SGEI, OP_LB, OP_LH, OP_LW, OP_LBU, OP_LHU, 
   OP_LF, OP_LD, OP_SB, OP_SH, OP_SW, OP_SF, OP_SD, OP_ITLB, OP_SLTUI, 
   OP_SGTUI, OP_SLEUI, OP_SGEUI, OP_J, OP_JAL, OP_NOP);
attribute ENUM_ENCODING of aluOp : type is 
   "0000000 0000001 0000010 0000011 0000100 0000101 0000110 0000111 0001000 0001001 0001010 0001011 0001100 0001101 0001110 0001111 0010000 0010001 0010010 0010011 0010100 0010101 0010110 0010111 0011000 0011001 0011010 0011011 0011100 0011101 0011110 0011111 0100000 0100001 0100010 0100011 0100100 0100101 0100110 0100111 0101000 0101001 0101010 0101011 0101100 0101101 0101110 0101111 0110000 0110001 0110010 0110011 0110100 0110101 0110110 0110111 0111000 0111001 0111010 0111011 0111100 0111101 0111110 0111111 1000000 1000001 1000010 1000011 1000100 1000101 1000110 1000111 1001000 1001001 1001010 1001011 1001100 1001101 1001110 1001111 1010000 1010001 1010010 1010011 1010100 1010101 1010110 1010111 1011000 1011001 1011010 1011011 1011100 1011101 1011110 1011111 1100000 1100001 1100010 1100011 1100100 1100101 1100110";
   
   -- Declarations for conversion functions.
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when OP_SLL => return "0000000";
         when OP_SRL => return "0000001";
         when OP_SRA => return "0000010";
         when OP_ADD => return "0000011";
         when OP_ADDU => return "0000100";
         when OP_SUB => return "0000101";
         when OP_SUBU => return "0000110";
         when OP_AND => return "0000111";
         when OP_OR => return "0001000";
         when OP_XOR => return "0001001";
         when OP_SEQ => return "0001010";
         when OP_SNE => return "0001011";
         when OP_SLT => return "0001100";
         when OP_SGT => return "0001101";
         when OP_SLE => return "0001110";
         when OP_SGE => return "0001111";
         when OP_MOVI2S => return "0010000";
         when OP_MOVS2I => return "0010001";
         when OP_MOVF => return "0010010";
         when OP_MOVD => return "0010011";
         when OP_MOVFP2I => return "0010100";
         when OP_MOVI2FP => return "0010101";
         when OP_MOVI2T => return "0010110";
         when OP_MOVT2I => return "0010111";
         when OP_SLTU => return "0011000";
         when OP_SGTU => return "0011001";
         when OP_SLEU => return "0011010";
         when OP_SGEU => return "0011011";
         when OP_ADDF => return "0011100";
         when OP_SUBF => return "0011101";
         when OP_MULTF => return "0011110";
         when OP_DIVF => return "0011111";
         when OP_ADDD => return "0100000";
         when OP_SUBD => return "0100001";
         when OP_MULTD => return "0100010";
         when OP_DIVD => return "0100011";
         when OP_CVTF2D => return "0100100";
         when OP_CVTF2I => return "0100101";
         when OP_CVTD2F => return "0100110";
         when OP_CVTD2I => return "0100111";
         when OP_CVTI2F => return "0101000";
         when OP_CVTI2D => return "0101001";
         when OP_MULT => return "0101010";
         when OP_DIV => return "0101011";
         when OP_EQF => return "0101100";
         when OP_NEF => return "0101101";
         when OP_LTF => return "0101110";
         when OP_GTF => return "0101111";
         when OP_LEF => return "0110000";
         when OP_GEF => return "0110001";
         when OP_MULTU => return "0110010";
         when OP_DIVU => return "0110011";
         when OP_EQD => return "0110100";
         when OP_NED => return "0110101";
         when OP_LTD => return "0110110";
         when OP_GTD => return "0110111";
         when OP_LED => return "0111000";
         when OP_GED => return "0111001";
         when OP_BEQZ => return "0111010";
         when OP_BNEZ => return "0111011";
         when OP_BFPT => return "0111100";
         when OP_BFPF => return "0111101";
         when OP_ADDI => return "0111110";
         when OP_ADDUI => return "0111111";
         when OP_SUBI => return "1000000";
         when OP_SUBUI => return "1000001";
         when OP_ANDI => return "1000010";
         when OP_ORI => return "1000011";
         when OP_XORI => return "1000100";
         when OP_LHI => return "1000101";
         when OP_RFE => return "1000110";
         when OP_TRAP => return "1000111";
         when OP_JR => return "1001000";
         when OP_JALR => return "1001001";
         when OP_SLLI => return "1001010";
         when OP_SRLI => return "1001011";
         when OP_SRAI => return "1001100";
         when OP_SEQI => return "1001101";
         when OP_SNEI => return "1001110";
         when OP_SLTI => return "1001111";
         when OP_SGTI => return "1010000";
         when OP_SLEI => return "1010001";
         when OP_SGEI => return "1010010";
         when OP_LB => return "1010011";
         when OP_LH => return "1010100";
         when OP_LW => return "1010101";
         when OP_LBU => return "1010110";
         when OP_LHU => return "1010111";
         when OP_LF => return "1011000";
         when OP_LD => return "1011001";
         when OP_SB => return "1011010";
         when OP_SH => return "1011011";
         when OP_SW => return "1011100";
         when OP_SF => return "1011101";
         when OP_SD => return "1011110";
         when OP_ITLB => return "1011111";
         when OP_SLTUI => return "1100000";
         when OP_SGTUI => return "1100001";
         when OP_SLEUI => return "1100010";
         when OP_SGEUI => return "1100011";
         when OP_J => return "1100100";
         when OP_JAL => return "1100101";
         when OP_NOP => return "1100110";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

   port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  DOUT :
         out std_logic_vector (31 downto 0));

end DLX_IRAM_RAM_DEPTH256_I_SIZE32;

architecture SYN_BEHAVIORAL of DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_DRAM_N256_NW32 is

   port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector (31 
         downto 0);  DOUT : out std_logic_vector (31 downto 0));

end DLX_DRAM_N256_NW32;

architecture SYN_BEHAVIORAL of DLX_DRAM_N256_NW32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RF_N32_NA5 is

   port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
         ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_N32_NA5;

architecture SYN_BEHAVIORAL of RF_N32_NA5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REG_0_31_port, REG_0_30_port, REG_0_29_port, REG_0_28_port, 
      REG_0_27_port, REG_0_26_port, REG_0_25_port, REG_0_24_port, REG_0_23_port
      , REG_0_22_port, REG_0_21_port, REG_0_20_port, REG_0_19_port, 
      REG_0_18_port, REG_0_17_port, REG_0_16_port, REG_0_15_port, REG_0_14_port
      , REG_0_13_port, REG_0_12_port, REG_0_11_port, REG_0_10_port, 
      REG_0_9_port, REG_0_8_port, REG_0_7_port, REG_0_6_port, REG_0_5_port, 
      REG_0_4_port, REG_0_3_port, REG_0_2_port, REG_0_1_port, REG_0_0_port, 
      REG_31_31_port, REG_31_30_port, REG_31_29_port, REG_31_28_port, 
      REG_31_27_port, REG_31_26_port, REG_31_25_port, REG_31_24_port, 
      REG_31_23_port, REG_31_22_port, REG_31_21_port, REG_31_20_port, 
      REG_31_19_port, REG_31_18_port, REG_31_17_port, REG_31_16_port, 
      REG_31_15_port, REG_31_14_port, REG_31_13_port, REG_31_12_port, 
      REG_31_11_port, REG_31_10_port, REG_31_9_port, REG_31_8_port, 
      REG_31_7_port, REG_31_6_port, REG_31_5_port, REG_31_4_port, REG_31_3_port
      , REG_31_2_port, REG_31_1_port, REG_31_0_port, N156, N157, N158, N159, 
      N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, 
      N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, 
      N184, N185, N186, N187, N219, N220, N221, N222, N223, N224, N225, N226, 
      N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, 
      N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, 
      n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51 : 
      std_logic;

begin
   
   REG_reg_0_31_inst : DLH_X1 port map( G => n10, D => N250, Q => REG_0_31_port
                           );
   REG_reg_0_30_inst : DLH_X1 port map( G => n10, D => N249, Q => REG_0_30_port
                           );
   REG_reg_0_29_inst : DLH_X1 port map( G => n10, D => N248, Q => REG_0_29_port
                           );
   REG_reg_0_28_inst : DLH_X1 port map( G => n10, D => N247, Q => REG_0_28_port
                           );
   REG_reg_0_27_inst : DLH_X1 port map( G => n11, D => N246, Q => REG_0_27_port
                           );
   REG_reg_0_26_inst : DLH_X1 port map( G => n11, D => N245, Q => REG_0_26_port
                           );
   REG_reg_0_25_inst : DLH_X1 port map( G => n11, D => N244, Q => REG_0_25_port
                           );
   REG_reg_0_24_inst : DLH_X1 port map( G => n11, D => N243, Q => REG_0_24_port
                           );
   REG_reg_0_23_inst : DLH_X1 port map( G => n11, D => N242, Q => REG_0_23_port
                           );
   REG_reg_0_22_inst : DLH_X1 port map( G => n11, D => N241, Q => REG_0_22_port
                           );
   REG_reg_0_21_inst : DLH_X1 port map( G => n12, D => N240, Q => REG_0_21_port
                           );
   REG_reg_0_20_inst : DLH_X1 port map( G => n12, D => N239, Q => REG_0_20_port
                           );
   REG_reg_0_19_inst : DLH_X1 port map( G => n12, D => N238, Q => REG_0_19_port
                           );
   REG_reg_0_18_inst : DLH_X1 port map( G => n12, D => N237, Q => REG_0_18_port
                           );
   REG_reg_0_17_inst : DLH_X1 port map( G => n10, D => N236, Q => REG_0_17_port
                           );
   REG_reg_0_16_inst : DLH_X1 port map( G => n10, D => N235, Q => REG_0_16_port
                           );
   REG_reg_0_15_inst : DLH_X1 port map( G => n10, D => N234, Q => REG_0_15_port
                           );
   REG_reg_0_14_inst : DLH_X1 port map( G => n10, D => N233, Q => REG_0_14_port
                           );
   REG_reg_0_13_inst : DLH_X1 port map( G => n10, D => N232, Q => REG_0_13_port
                           );
   REG_reg_0_12_inst : DLH_X1 port map( G => n10, D => N231, Q => REG_0_12_port
                           );
   REG_reg_0_11_inst : DLH_X1 port map( G => n12, D => N230, Q => REG_0_11_port
                           );
   REG_reg_0_10_inst : DLH_X1 port map( G => n12, D => N229, Q => REG_0_10_port
                           );
   REG_reg_0_9_inst : DLH_X1 port map( G => n12, D => N228, Q => REG_0_9_port);
   REG_reg_0_8_inst : DLH_X1 port map( G => n12, D => N227, Q => REG_0_8_port);
   REG_reg_0_7_inst : DLH_X1 port map( G => n12, D => N226, Q => REG_0_7_port);
   REG_reg_0_6_inst : DLH_X1 port map( G => n12, D => N225, Q => REG_0_6_port);
   REG_reg_0_5_inst : DLH_X1 port map( G => n12, D => N224, Q => REG_0_5_port);
   REG_reg_0_4_inst : DLH_X1 port map( G => n12, D => N223, Q => REG_0_4_port);
   REG_reg_0_3_inst : DLH_X1 port map( G => n12, D => N222, Q => REG_0_3_port);
   REG_reg_0_2_inst : DLH_X1 port map( G => n12, D => N221, Q => REG_0_2_port);
   REG_reg_0_1_inst : DLH_X1 port map( G => n11, D => N220, Q => REG_0_1_port);
   REG_reg_0_0_inst : DLH_X1 port map( G => n11, D => N219, Q => REG_0_0_port);
   REG_reg_31_31_inst : DLH_X1 port map( G => n12, D => N187, Q => 
                           REG_31_31_port);
   REG_reg_31_30_inst : DLH_X1 port map( G => n12, D => N186, Q => 
                           REG_31_30_port);
   REG_reg_31_29_inst : DLH_X1 port map( G => n11, D => N185, Q => 
                           REG_31_29_port);
   REG_reg_31_28_inst : DLH_X1 port map( G => n11, D => N184, Q => 
                           REG_31_28_port);
   REG_reg_31_27_inst : DLH_X1 port map( G => n12, D => N183, Q => 
                           REG_31_27_port);
   REG_reg_31_26_inst : DLH_X1 port map( G => n12, D => N182, Q => 
                           REG_31_26_port);
   REG_reg_31_25_inst : DLH_X1 port map( G => n12, D => N181, Q => 
                           REG_31_25_port);
   REG_reg_31_24_inst : DLH_X1 port map( G => n12, D => N180, Q => 
                           REG_31_24_port);
   REG_reg_31_23_inst : DLH_X1 port map( G => n11, D => N179, Q => 
                           REG_31_23_port);
   REG_reg_31_22_inst : DLH_X1 port map( G => n11, D => N178, Q => 
                           REG_31_22_port);
   REG_reg_31_21_inst : DLH_X1 port map( G => n11, D => N177, Q => 
                           REG_31_21_port);
   REG_reg_31_20_inst : DLH_X1 port map( G => n11, D => N176, Q => 
                           REG_31_20_port);
   REG_reg_31_19_inst : DLH_X1 port map( G => n11, D => N175, Q => 
                           REG_31_19_port);
   REG_reg_31_18_inst : DLH_X1 port map( G => n11, D => N174, Q => 
                           REG_31_18_port);
   REG_reg_31_17_inst : DLH_X1 port map( G => n11, D => N173, Q => 
                           REG_31_17_port);
   REG_reg_31_16_inst : DLH_X1 port map( G => n11, D => N172, Q => 
                           REG_31_16_port);
   REG_reg_31_15_inst : DLH_X1 port map( G => n11, D => N171, Q => 
                           REG_31_15_port);
   REG_reg_31_14_inst : DLH_X1 port map( G => n11, D => N170, Q => 
                           REG_31_14_port);
   REG_reg_31_13_inst : DLH_X1 port map( G => n12, D => N169, Q => 
                           REG_31_13_port);
   REG_reg_31_12_inst : DLH_X1 port map( G => n11, D => N168, Q => 
                           REG_31_12_port);
   REG_reg_31_11_inst : DLH_X1 port map( G => n11, D => N167, Q => 
                           REG_31_11_port);
   REG_reg_31_10_inst : DLH_X1 port map( G => n12, D => N166, Q => 
                           REG_31_10_port);
   REG_reg_31_9_inst : DLH_X1 port map( G => n12, D => N165, Q => REG_31_9_port
                           );
   REG_reg_31_8_inst : DLH_X1 port map( G => n12, D => N164, Q => REG_31_8_port
                           );
   REG_reg_31_7_inst : DLH_X1 port map( G => n12, D => N163, Q => REG_31_7_port
                           );
   REG_reg_31_6_inst : DLH_X1 port map( G => n12, D => N162, Q => REG_31_6_port
                           );
   REG_reg_31_5_inst : DLH_X1 port map( G => n12, D => N161, Q => REG_31_5_port
                           );
   REG_reg_31_4_inst : DLH_X1 port map( G => n12, D => N160, Q => REG_31_4_port
                           );
   REG_reg_31_3_inst : DLH_X1 port map( G => n12, D => N159, Q => REG_31_3_port
                           );
   REG_reg_31_2_inst : DLH_X1 port map( G => n12, D => N158, Q => REG_31_2_port
                           );
   REG_reg_31_1_inst : DLH_X1 port map( G => n11, D => N157, Q => REG_31_1_port
                           );
   REG_reg_31_0_inst : DLH_X1 port map( G => n11, D => N156, Q => REG_31_0_port
                           );
   U3 : CLKBUF_X2 port map( A => n51, Z => n7);
   U4 : CLKBUF_X2 port map( A => n49, Z => n8);
   U5 : INV_X1 port map( A => RST, ZN => n11);
   U6 : INV_X1 port map( A => RST, ZN => n12);
   U7 : INV_X1 port map( A => RST, ZN => n10);
   U8 : OR4_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), A3 => ADD_WR(0), A4 
                           => ADD_WR(2), ZN => n13);
   U9 : NOR2_X1 port map( A1 => ADD_WR(1), A2 => n13, ZN => n36);
   U10 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(0), ZN => n14);
   U11 : INV_X1 port map( A => n14, ZN => N156);
   U12 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(31), ZN => n46);
   U13 : INV_X1 port map( A => n46, ZN => N187);
   U14 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(30), ZN => n45);
   U15 : INV_X1 port map( A => n45, ZN => N186);
   U16 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(29), ZN => n44);
   U17 : INV_X1 port map( A => n44, ZN => N185);
   U18 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(28), ZN => n43);
   U19 : INV_X1 port map( A => n43, ZN => N184);
   U20 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(27), ZN => n42);
   U21 : INV_X1 port map( A => n42, ZN => N183);
   U22 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(26), ZN => n41);
   U23 : INV_X1 port map( A => n41, ZN => N182);
   U24 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(25), ZN => n40);
   U25 : INV_X1 port map( A => n40, ZN => N181);
   U26 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(24), ZN => n39);
   U27 : INV_X1 port map( A => n39, ZN => N180);
   U28 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(23), ZN => n38);
   U29 : INV_X1 port map( A => n38, ZN => N179);
   U30 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(22), ZN => n37);
   U31 : INV_X1 port map( A => n37, ZN => N178);
   U32 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(21), ZN => n35);
   U33 : INV_X1 port map( A => n35, ZN => N177);
   U34 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(20), ZN => n34);
   U35 : INV_X1 port map( A => n34, ZN => N176);
   U36 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(19), ZN => n33);
   U37 : INV_X1 port map( A => n33, ZN => N175);
   U38 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(18), ZN => n32);
   U39 : INV_X1 port map( A => n32, ZN => N174);
   U40 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(17), ZN => n31);
   U41 : INV_X1 port map( A => n31, ZN => N173);
   U42 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(16), ZN => n30);
   U43 : INV_X1 port map( A => n30, ZN => N172);
   U44 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(15), ZN => n29);
   U45 : INV_X1 port map( A => n29, ZN => N171);
   U46 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(14), ZN => n28);
   U47 : INV_X1 port map( A => n28, ZN => N170);
   U48 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(13), ZN => n27);
   U49 : INV_X1 port map( A => n27, ZN => N169);
   U50 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(12), ZN => n26);
   U51 : INV_X1 port map( A => n26, ZN => N168);
   U52 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(11), ZN => n25);
   U53 : INV_X1 port map( A => n25, ZN => N167);
   U54 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(10), ZN => n24);
   U55 : INV_X1 port map( A => n24, ZN => N166);
   U56 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(9), ZN => n23);
   U57 : INV_X1 port map( A => n23, ZN => N165);
   U58 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(8), ZN => n22);
   U59 : INV_X1 port map( A => n22, ZN => N164);
   U60 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(7), ZN => n21);
   U61 : INV_X1 port map( A => n21, ZN => N163);
   U62 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(6), ZN => n20);
   U63 : INV_X1 port map( A => n20, ZN => N162);
   U64 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(5), ZN => n19);
   U65 : INV_X1 port map( A => n19, ZN => N161);
   U66 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(4), ZN => n18);
   U67 : INV_X1 port map( A => n18, ZN => N160);
   U68 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(3), ZN => n17);
   U69 : INV_X1 port map( A => n17, ZN => N159);
   U70 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(2), ZN => n16);
   U71 : INV_X1 port map( A => n16, ZN => N158);
   U72 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(1), ZN => n15);
   U73 : INV_X1 port map( A => n15, ZN => N157);
   U74 : CLKBUF_X1 port map( A => n36, Z => n47);
   U75 : NOR2_X1 port map( A1 => n47, A2 => n14, ZN => N219);
   U76 : NOR2_X1 port map( A1 => n47, A2 => n15, ZN => N220);
   U77 : NOR2_X1 port map( A1 => n47, A2 => n16, ZN => N221);
   U78 : NOR2_X1 port map( A1 => n47, A2 => n17, ZN => N222);
   U79 : NOR2_X1 port map( A1 => n47, A2 => n18, ZN => N223);
   U80 : NOR2_X1 port map( A1 => n47, A2 => n19, ZN => N224);
   U81 : NOR2_X1 port map( A1 => n47, A2 => n20, ZN => N225);
   U82 : NOR2_X1 port map( A1 => n47, A2 => n21, ZN => N226);
   U83 : NOR2_X1 port map( A1 => n47, A2 => n22, ZN => N227);
   U84 : NOR2_X1 port map( A1 => n47, A2 => n23, ZN => N228);
   U85 : NOR2_X1 port map( A1 => n36, A2 => n24, ZN => N229);
   U86 : NOR2_X1 port map( A1 => n47, A2 => n25, ZN => N230);
   U87 : NOR2_X1 port map( A1 => n47, A2 => n26, ZN => N231);
   U88 : NOR2_X1 port map( A1 => n36, A2 => n27, ZN => N232);
   U89 : NOR2_X1 port map( A1 => n36, A2 => n28, ZN => N233);
   U90 : NOR2_X1 port map( A1 => n36, A2 => n29, ZN => N234);
   U91 : NOR2_X1 port map( A1 => n36, A2 => n30, ZN => N235);
   U92 : NOR2_X1 port map( A1 => n36, A2 => n31, ZN => N236);
   U93 : NOR2_X1 port map( A1 => n36, A2 => n32, ZN => N237);
   U94 : NOR2_X1 port map( A1 => n36, A2 => n33, ZN => N238);
   U95 : NOR2_X1 port map( A1 => n36, A2 => n34, ZN => N239);
   U96 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => N240);
   U97 : NOR2_X1 port map( A1 => n47, A2 => n37, ZN => N241);
   U98 : NOR2_X1 port map( A1 => n47, A2 => n38, ZN => N242);
   U99 : NOR2_X1 port map( A1 => n47, A2 => n39, ZN => N243);
   U100 : NOR2_X1 port map( A1 => n47, A2 => n40, ZN => N244);
   U101 : NOR2_X1 port map( A1 => n47, A2 => n41, ZN => N245);
   U102 : NOR2_X1 port map( A1 => n47, A2 => n42, ZN => N246);
   U103 : NOR2_X1 port map( A1 => n47, A2 => n43, ZN => N247);
   U104 : NOR2_X1 port map( A1 => n47, A2 => n44, ZN => N248);
   U105 : NOR2_X1 port map( A1 => n47, A2 => n45, ZN => N249);
   U106 : NOR2_X1 port map( A1 => n47, A2 => n46, ZN => N250);
   U107 : OR4_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => ADD_RD2(2)
                           , A4 => ADD_RD2(4), ZN => n48);
   U108 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => n48, ZN => n49);
   U109 : MUX2_X1 port map( A => REG_31_31_port, B => REG_0_31_port, S => n8, Z
                           => OUT2(31));
   U110 : MUX2_X1 port map( A => REG_31_30_port, B => REG_0_30_port, S => n8, Z
                           => OUT2(30));
   U111 : MUX2_X1 port map( A => REG_31_29_port, B => REG_0_29_port, S => n8, Z
                           => OUT2(29));
   U112 : MUX2_X1 port map( A => REG_31_28_port, B => REG_0_28_port, S => n8, Z
                           => OUT2(28));
   U113 : MUX2_X1 port map( A => REG_31_27_port, B => REG_0_27_port, S => n8, Z
                           => OUT2(27));
   U114 : MUX2_X1 port map( A => REG_31_26_port, B => REG_0_26_port, S => n8, Z
                           => OUT2(26));
   U115 : MUX2_X1 port map( A => REG_31_25_port, B => REG_0_25_port, S => n8, Z
                           => OUT2(25));
   U116 : MUX2_X1 port map( A => REG_31_24_port, B => REG_0_24_port, S => n8, Z
                           => OUT2(24));
   U117 : MUX2_X1 port map( A => REG_31_23_port, B => REG_0_23_port, S => n8, Z
                           => OUT2(23));
   U118 : MUX2_X1 port map( A => REG_31_22_port, B => REG_0_22_port, S => n8, Z
                           => OUT2(22));
   U119 : MUX2_X1 port map( A => REG_31_21_port, B => REG_0_21_port, S => n8, Z
                           => OUT2(21));
   U120 : MUX2_X1 port map( A => REG_31_20_port, B => REG_0_20_port, S => n8, Z
                           => OUT2(20));
   U121 : MUX2_X1 port map( A => REG_31_19_port, B => REG_0_19_port, S => n8, Z
                           => OUT2(19));
   U122 : MUX2_X1 port map( A => REG_31_18_port, B => REG_0_18_port, S => n49, 
                           Z => OUT2(18));
   U123 : MUX2_X1 port map( A => REG_31_17_port, B => REG_0_17_port, S => n49, 
                           Z => OUT2(17));
   U124 : MUX2_X1 port map( A => REG_31_16_port, B => REG_0_16_port, S => n49, 
                           Z => OUT2(16));
   U125 : MUX2_X1 port map( A => REG_31_15_port, B => REG_0_15_port, S => n49, 
                           Z => OUT2(15));
   U126 : MUX2_X1 port map( A => REG_31_14_port, B => REG_0_14_port, S => n49, 
                           Z => OUT2(14));
   U127 : MUX2_X1 port map( A => REG_31_13_port, B => REG_0_13_port, S => n49, 
                           Z => OUT2(13));
   U128 : MUX2_X1 port map( A => REG_31_12_port, B => REG_0_12_port, S => n49, 
                           Z => OUT2(12));
   U129 : MUX2_X1 port map( A => REG_31_11_port, B => REG_0_11_port, S => n49, 
                           Z => OUT2(11));
   U130 : MUX2_X1 port map( A => REG_31_10_port, B => REG_0_10_port, S => n49, 
                           Z => OUT2(10));
   U131 : MUX2_X1 port map( A => REG_31_9_port, B => REG_0_9_port, S => n8, Z 
                           => OUT2(9));
   U132 : MUX2_X1 port map( A => REG_31_8_port, B => REG_0_8_port, S => n8, Z 
                           => OUT2(8));
   U133 : MUX2_X1 port map( A => REG_31_7_port, B => REG_0_7_port, S => n8, Z 
                           => OUT2(7));
   U134 : MUX2_X1 port map( A => REG_31_6_port, B => REG_0_6_port, S => n8, Z 
                           => OUT2(6));
   U135 : MUX2_X1 port map( A => REG_31_5_port, B => REG_0_5_port, S => n8, Z 
                           => OUT2(5));
   U136 : MUX2_X1 port map( A => REG_31_4_port, B => REG_0_4_port, S => n8, Z 
                           => OUT2(4));
   U137 : MUX2_X1 port map( A => REG_31_3_port, B => REG_0_3_port, S => n8, Z 
                           => OUT2(3));
   U138 : MUX2_X1 port map( A => REG_31_2_port, B => REG_0_2_port, S => n8, Z 
                           => OUT2(2));
   U139 : MUX2_X1 port map( A => REG_31_1_port, B => REG_0_1_port, S => n8, Z 
                           => OUT2(1));
   U140 : MUX2_X1 port map( A => REG_31_0_port, B => REG_0_0_port, S => n8, Z 
                           => OUT2(0));
   U141 : OR4_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => ADD_RD1(2)
                           , A4 => ADD_RD1(4), ZN => n50);
   U142 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => n50, ZN => n51);
   U143 : MUX2_X1 port map( A => REG_31_31_port, B => REG_0_31_port, S => n7, Z
                           => OUT1(31));
   U144 : MUX2_X1 port map( A => REG_31_30_port, B => REG_0_30_port, S => n7, Z
                           => OUT1(30));
   U145 : MUX2_X1 port map( A => REG_31_29_port, B => REG_0_29_port, S => n7, Z
                           => OUT1(29));
   U146 : MUX2_X1 port map( A => REG_31_28_port, B => REG_0_28_port, S => n7, Z
                           => OUT1(28));
   U147 : MUX2_X1 port map( A => REG_31_27_port, B => REG_0_27_port, S => n7, Z
                           => OUT1(27));
   U148 : MUX2_X1 port map( A => REG_31_26_port, B => REG_0_26_port, S => n7, Z
                           => OUT1(26));
   U149 : MUX2_X1 port map( A => REG_31_25_port, B => REG_0_25_port, S => n7, Z
                           => OUT1(25));
   U150 : MUX2_X1 port map( A => REG_31_24_port, B => REG_0_24_port, S => n7, Z
                           => OUT1(24));
   U151 : MUX2_X1 port map( A => REG_31_23_port, B => REG_0_23_port, S => n7, Z
                           => OUT1(23));
   U152 : MUX2_X1 port map( A => REG_31_22_port, B => REG_0_22_port, S => n7, Z
                           => OUT1(22));
   U153 : MUX2_X1 port map( A => REG_31_21_port, B => REG_0_21_port, S => n7, Z
                           => OUT1(21));
   U154 : MUX2_X1 port map( A => REG_31_20_port, B => REG_0_20_port, S => n7, Z
                           => OUT1(20));
   U155 : MUX2_X1 port map( A => REG_31_19_port, B => REG_0_19_port, S => n7, Z
                           => OUT1(19));
   U156 : MUX2_X1 port map( A => REG_31_18_port, B => REG_0_18_port, S => n51, 
                           Z => OUT1(18));
   U157 : MUX2_X1 port map( A => REG_31_17_port, B => REG_0_17_port, S => n51, 
                           Z => OUT1(17));
   U158 : MUX2_X1 port map( A => REG_31_16_port, B => REG_0_16_port, S => n51, 
                           Z => OUT1(16));
   U159 : MUX2_X1 port map( A => REG_31_15_port, B => REG_0_15_port, S => n51, 
                           Z => OUT1(15));
   U160 : MUX2_X1 port map( A => REG_31_14_port, B => REG_0_14_port, S => n51, 
                           Z => OUT1(14));
   U161 : MUX2_X1 port map( A => REG_31_13_port, B => REG_0_13_port, S => n51, 
                           Z => OUT1(13));
   U162 : MUX2_X1 port map( A => REG_31_12_port, B => REG_0_12_port, S => n51, 
                           Z => OUT1(12));
   U163 : MUX2_X1 port map( A => REG_31_11_port, B => REG_0_11_port, S => n51, 
                           Z => OUT1(11));
   U164 : MUX2_X1 port map( A => REG_31_10_port, B => REG_0_10_port, S => n51, 
                           Z => OUT1(10));
   U165 : MUX2_X1 port map( A => REG_31_9_port, B => REG_0_9_port, S => n7, Z 
                           => OUT1(9));
   U166 : MUX2_X1 port map( A => REG_31_8_port, B => REG_0_8_port, S => n7, Z 
                           => OUT1(8));
   U167 : MUX2_X1 port map( A => REG_31_7_port, B => REG_0_7_port, S => n7, Z 
                           => OUT1(7));
   U168 : MUX2_X1 port map( A => REG_31_6_port, B => REG_0_6_port, S => n7, Z 
                           => OUT1(6));
   U169 : MUX2_X1 port map( A => REG_31_5_port, B => REG_0_5_port, S => n7, Z 
                           => OUT1(5));
   U170 : MUX2_X1 port map( A => REG_31_4_port, B => REG_0_4_port, S => n7, Z 
                           => OUT1(4));
   U171 : MUX2_X1 port map( A => REG_31_3_port, B => REG_0_3_port, S => n7, Z 
                           => OUT1(3));
   U172 : MUX2_X1 port map( A => REG_31_2_port, B => REG_0_2_port, S => n7, Z 
                           => OUT1(2));
   U173 : MUX2_X1 port map( A => REG_31_1_port, B => REG_0_1_port, S => n7, Z 
                           => OUT1(1));
   U174 : MUX2_X1 port map( A => REG_31_0_port, B => REG_0_0_port, S => n7, Z 
                           => OUT1(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_NB8 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
         std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);  Z
         : out std_logic);

end ALU_N32_NB8;

architecture SYN_BEHAVIORAL of ALU_N32_NB8 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X2
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal N96, OP_A_31_port, OP_A_30_port, OP_A_29_port, OP_A_28_port, 
      OP_A_27_port, OP_A_26_port, OP_A_25_port, OP_A_24_port, OP_A_23_port, 
      OP_A_22_port, OP_A_21_port, OP_A_20_port, OP_A_19_port, OP_A_18_port, 
      OP_A_17_port, OP_A_16_port, OP_A_15_port, OP_A_14_port, OP_A_13_port, 
      OP_A_12_port, OP_A_11_port, OP_A_10_port, OP_A_9_port, OP_A_8_port, 
      OP_A_7_port, OP_A_6_port, OP_A_5_port, OP_A_4_port, OP_A_3_port, 
      OP_A_2_port, OP_A_1_port, OP_A_0_port, OP_B_31_port, OP_B_30_port, 
      OP_B_29_port, OP_B_28_port, OP_B_27_port, OP_B_26_port, OP_B_25_port, 
      OP_B_24_port, OP_B_23_port, OP_B_22_port, OP_B_21_port, OP_B_20_port, 
      OP_B_19_port, OP_B_18_port, OP_B_17_port, OP_B_16_port, OP_B_15_port, 
      OP_B_14_port, OP_B_13_port, OP_B_12_port, OP_B_11_port, OP_B_10_port, 
      OP_B_9_port, OP_B_8_port, OP_B_7_port, OP_B_6_port, OP_B_5_port, 
      OP_B_4_port, OP_B_3_port, OP_B_2_port, OP_B_1_port, OP_B_0_port, OP_Ci, 
      OP_LOGIC_1_port, OP_LOGIC_0_port, OP_SHIFT, OP_COMPARE_3_port, 
      OP_COMPARE_2_port, OP_COMPARE_1_port, OP_COMPARE_0_port, N246, N247, N248
      , N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
      N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, 
      N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, 
      N285, N286, N287, N288, N289, C431_DATA4_3, C431_DATA4_4, C431_DATA4_5, 
      C431_DATA4_6, C431_DATA4_7, C431_DATA4_8, C431_DATA4_9, C431_DATA4_10, 
      C431_DATA4_11, C431_DATA4_12, C431_DATA4_13, C431_DATA4_14, C431_DATA4_15
      , C431_DATA4_16, C431_DATA4_17, C430_DATA4_5, C430_DATA4_6, C430_DATA4_7,
      C430_DATA4_8, C430_DATA4_9, C430_DATA4_10, C430_DATA4_11, C430_DATA4_12, 
      C430_DATA4_13, C430_DATA4_14, C430_DATA4_15, C430_DATA4_16, C430_DATA4_17
      , C430_DATA4_18, C430_DATA4_19, C429_DATA4_7, C429_DATA4_8, C429_DATA4_9,
      C429_DATA4_10, C429_DATA4_11, C429_DATA4_12, C429_DATA4_13, C429_DATA4_14
      , C429_DATA4_15, C429_DATA4_16, C429_DATA4_17, C429_DATA4_18, 
      C429_DATA4_19, C429_DATA4_20, C429_DATA4_21, C428_DATA4_1, C428_DATA4_2, 
      C428_DATA4_3, C428_DATA4_4, C428_DATA4_5, C428_DATA4_6, C428_DATA4_7, 
      C428_DATA4_8, C428_DATA4_9, C428_DATA4_10, C428_DATA4_11, C428_DATA4_12, 
      C428_DATA4_13, C428_DATA4_14, C428_DATA4_15, C2_DATA1_2, C2_DATA1_4, 
      C2_DATA1_6, DP_OP_440J3_122_9847_n80, DP_OP_440J3_122_9847_n79, 
      DP_OP_440J3_122_9847_n78, DP_OP_440J3_122_9847_n77, 
      DP_OP_440J3_122_9847_n76, DP_OP_440J3_122_9847_n75, 
      DP_OP_440J3_122_9847_n74, DP_OP_440J3_122_9847_n73, 
      DP_OP_440J3_122_9847_n72, DP_OP_440J3_122_9847_n71, 
      DP_OP_440J3_122_9847_n70, DP_OP_440J3_122_9847_n69, 
      DP_OP_440J3_122_9847_n68, DP_OP_440J3_122_9847_n67, 
      DP_OP_440J3_122_9847_n66, DP_OP_440J3_122_9847_n35, 
      DP_OP_440J3_122_9847_n34, DP_OP_440J3_122_9847_n33, 
      DP_OP_440J3_122_9847_n32, DP_OP_440J3_122_9847_n31, 
      DP_OP_440J3_122_9847_n30, DP_OP_440J3_122_9847_n29, 
      DP_OP_440J3_122_9847_n28, DP_OP_440J3_122_9847_n27, 
      DP_OP_440J3_122_9847_n26, DP_OP_440J3_122_9847_n25, 
      DP_OP_440J3_122_9847_n24, DP_OP_440J3_122_9847_n23, 
      DP_OP_440J3_122_9847_n22, DP_OP_440J3_122_9847_n21, 
      DP_OP_440J3_122_9847_n20, DP_OP_446J3_125_4819_n87, 
      DP_OP_446J3_125_4819_n86, DP_OP_446J3_125_4819_n85, 
      DP_OP_446J3_125_4819_n84, DP_OP_446J3_125_4819_n83, 
      DP_OP_446J3_125_4819_n82, DP_OP_446J3_125_4819_n81, 
      DP_OP_446J3_125_4819_n80, DP_OP_446J3_125_4819_n79, 
      DP_OP_446J3_125_4819_n78, DP_OP_446J3_125_4819_n77, 
      DP_OP_446J3_125_4819_n76, DP_OP_446J3_125_4819_n75, 
      DP_OP_446J3_125_4819_n74, DP_OP_446J3_125_4819_n73, 
      DP_OP_446J3_125_4819_n72, DP_OP_446J3_125_4819_n27, 
      DP_OP_446J3_125_4819_n26, DP_OP_446J3_125_4819_n25, 
      DP_OP_446J3_125_4819_n24, DP_OP_446J3_125_4819_n23, 
      DP_OP_446J3_125_4819_n22, DP_OP_446J3_125_4819_n21, 
      DP_OP_446J3_125_4819_n20, DP_OP_446J3_125_4819_n19, 
      DP_OP_446J3_125_4819_n18, DP_OP_446J3_125_4819_n17, 
      DP_OP_446J3_125_4819_n16, DP_OP_446J3_125_4819_n15, 
      DP_OP_446J3_125_4819_n14, DP_OP_446J3_125_4819_n13, 
      DP_OP_446J3_125_4819_n12, DP_OP_451J3_128_3502_n85, 
      DP_OP_451J3_128_3502_n84, DP_OP_451J3_128_3502_n83, 
      DP_OP_451J3_128_3502_n82, DP_OP_451J3_128_3502_n81, 
      DP_OP_451J3_128_3502_n80, DP_OP_451J3_128_3502_n79, 
      DP_OP_451J3_128_3502_n78, DP_OP_451J3_128_3502_n77, 
      DP_OP_451J3_128_3502_n76, DP_OP_451J3_128_3502_n75, 
      DP_OP_451J3_128_3502_n74, DP_OP_451J3_128_3502_n73, 
      DP_OP_451J3_128_3502_n72, DP_OP_451J3_128_3502_n71, 
      DP_OP_451J3_128_3502_n70, DP_OP_451J3_128_3502_n30, 
      DP_OP_451J3_128_3502_n29, DP_OP_451J3_128_3502_n28, 
      DP_OP_451J3_128_3502_n27, DP_OP_451J3_128_3502_n26, 
      DP_OP_451J3_128_3502_n25, DP_OP_451J3_128_3502_n24, 
      DP_OP_451J3_128_3502_n23, DP_OP_451J3_128_3502_n22, 
      DP_OP_451J3_128_3502_n21, DP_OP_451J3_128_3502_n20, 
      DP_OP_451J3_128_3502_n19, DP_OP_451J3_128_3502_n18, 
      DP_OP_451J3_128_3502_n17, DP_OP_451J3_128_3502_n16, 
      DP_OP_451J3_128_3502_n15, DP_OP_456J3_131_2158_n82, 
      DP_OP_456J3_131_2158_n81, DP_OP_456J3_131_2158_n80, 
      DP_OP_456J3_131_2158_n79, DP_OP_456J3_131_2158_n78, 
      DP_OP_456J3_131_2158_n77, DP_OP_456J3_131_2158_n76, 
      DP_OP_456J3_131_2158_n75, DP_OP_456J3_131_2158_n74, 
      DP_OP_456J3_131_2158_n73, DP_OP_456J3_131_2158_n72, 
      DP_OP_456J3_131_2158_n71, DP_OP_456J3_131_2158_n70, 
      DP_OP_456J3_131_2158_n69, DP_OP_456J3_131_2158_n68, 
      DP_OP_456J3_131_2158_n67, DP_OP_456J3_131_2158_n32, 
      DP_OP_456J3_131_2158_n31, DP_OP_456J3_131_2158_n30, 
      DP_OP_456J3_131_2158_n29, DP_OP_456J3_131_2158_n28, 
      DP_OP_456J3_131_2158_n27, DP_OP_456J3_131_2158_n26, 
      DP_OP_456J3_131_2158_n25, DP_OP_456J3_131_2158_n24, 
      DP_OP_456J3_131_2158_n23, DP_OP_456J3_131_2158_n22, 
      DP_OP_456J3_131_2158_n21, DP_OP_456J3_131_2158_n20, 
      DP_OP_456J3_131_2158_n19, DP_OP_456J3_131_2158_n18, 
      DP_OP_456J3_131_2158_n17, intadd_0_A_16_port, intadd_0_A_12_port, 
      intadd_0_A_11_port, intadd_0_A_10_port, intadd_0_A_9_port, 
      intadd_0_A_8_port, intadd_0_A_7_port, intadd_0_A_6_port, 
      intadd_0_A_5_port, intadd_0_A_4_port, intadd_0_A_3_port, 
      intadd_0_A_2_port, intadd_0_A_1_port, intadd_0_A_0_port, 
      intadd_0_B_14_port, intadd_0_B_13_port, intadd_0_B_12_port, 
      intadd_0_B_11_port, intadd_0_B_10_port, intadd_0_B_9_port, 
      intadd_0_B_8_port, intadd_0_B_7_port, intadd_0_B_6_port, 
      intadd_0_B_5_port, intadd_0_B_4_port, intadd_0_B_3_port, 
      intadd_0_B_2_port, intadd_0_B_1_port, intadd_0_B_0_port, intadd_0_CI, 
      intadd_0_SUM_26_port, intadd_0_SUM_25_port, intadd_0_SUM_24_port, 
      intadd_0_SUM_23_port, intadd_0_SUM_22_port, intadd_0_SUM_21_port, 
      intadd_0_SUM_20_port, intadd_0_SUM_19_port, intadd_0_SUM_18_port, 
      intadd_0_SUM_17_port, intadd_0_SUM_16_port, intadd_0_SUM_15_port, 
      intadd_0_SUM_14_port, intadd_0_SUM_13_port, intadd_0_SUM_12_port, 
      intadd_0_SUM_11_port, intadd_0_SUM_10_port, intadd_0_SUM_9_port, 
      intadd_0_SUM_8_port, intadd_0_SUM_7_port, intadd_0_SUM_6_port, 
      intadd_0_SUM_5_port, intadd_0_SUM_4_port, intadd_0_SUM_3_port, 
      intadd_0_SUM_2_port, intadd_0_SUM_1_port, intadd_0_SUM_0_port, 
      intadd_0_n27, intadd_0_n26, intadd_0_n25, intadd_0_n24, intadd_0_n23, 
      intadd_0_n22, intadd_0_n21, intadd_0_n20, intadd_0_n19, intadd_0_n18, 
      intadd_0_n17, intadd_0_n16, intadd_0_n15, intadd_0_n14, intadd_0_n13, 
      intadd_0_n12, intadd_0_n11, intadd_0_n10, intadd_0_n9, intadd_0_n8, 
      intadd_0_n7, intadd_0_n6, intadd_0_n5, intadd_0_n4, intadd_0_n3, 
      intadd_0_n2, intadd_0_n1, intadd_1_A_0_port, intadd_1_B_18_port, 
      intadd_1_B_14_port, intadd_1_B_13_port, intadd_1_B_12_port, 
      intadd_1_B_11_port, intadd_1_B_10_port, intadd_1_B_9_port, 
      intadd_1_B_8_port, intadd_1_B_7_port, intadd_1_B_6_port, 
      intadd_1_B_5_port, intadd_1_B_4_port, intadd_1_B_3_port, 
      intadd_1_B_2_port, intadd_1_B_1_port, intadd_1_B_0_port, 
      intadd_1_SUM_24_port, intadd_1_SUM_23_port, intadd_1_SUM_22_port, 
      intadd_1_SUM_21_port, intadd_1_SUM_20_port, intadd_1_SUM_19_port, 
      intadd_1_SUM_18_port, intadd_1_SUM_17_port, intadd_1_SUM_16_port, 
      intadd_1_SUM_15_port, intadd_1_SUM_14_port, intadd_1_SUM_13_port, 
      intadd_1_SUM_12_port, intadd_1_SUM_11_port, intadd_1_SUM_10_port, 
      intadd_1_SUM_9_port, intadd_1_SUM_8_port, intadd_1_SUM_7_port, 
      intadd_1_SUM_6_port, intadd_1_SUM_5_port, intadd_1_SUM_4_port, 
      intadd_1_SUM_3_port, intadd_1_SUM_2_port, intadd_1_SUM_1_port, 
      intadd_1_SUM_0_port, intadd_1_n25, intadd_1_n24, intadd_1_n23, 
      intadd_1_n22, intadd_1_n21, intadd_1_n20, intadd_1_n19, intadd_1_n18, 
      intadd_1_n17, intadd_1_n16, intadd_1_n15, intadd_1_n14, intadd_1_n13, 
      intadd_1_n12, intadd_1_n11, intadd_1_n10, intadd_1_n9, intadd_1_n8, 
      intadd_1_n7, intadd_1_n6, intadd_1_n5, intadd_1_n4, intadd_1_n3, 
      intadd_1_n2, intadd_1_n1, intadd_2_A_9_port, intadd_2_A_8_port, 
      intadd_2_A_7_port, intadd_2_A_6_port, intadd_2_A_5_port, 
      intadd_2_A_4_port, intadd_2_A_3_port, intadd_2_A_2_port, 
      intadd_2_A_1_port, intadd_2_A_0_port, intadd_2_B_0_port, 
      intadd_2_SUM_9_port, intadd_2_SUM_8_port, intadd_2_SUM_7_port, 
      intadd_2_SUM_6_port, intadd_2_SUM_5_port, intadd_2_SUM_4_port, 
      intadd_2_SUM_3_port, intadd_2_SUM_2_port, intadd_2_SUM_1_port, 
      intadd_2_SUM_0_port, intadd_2_n10, intadd_2_n9, intadd_2_n8, intadd_2_n7,
      intadd_2_n6, intadd_2_n5, intadd_2_n4, intadd_2_n3, intadd_2_n2, 
      intadd_2_n1, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
      n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96_port, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246_port, n247_port, n248_port, 
      n249_port, n250_port, n251_port, n252_port, n253_port, n254_port, 
      n255_port, n256_port, n257_port, n258_port, n259_port, n260_port, 
      n261_port, n262_port, n263_port, n264_port, n265_port, n266_port, 
      n267_port, n268_port, n269_port, n270_port, n271_port, n272_port, 
      n273_port, n274_port, n275_port, n276_port, n277_port, n278_port, 
      n279_port, n280_port, n281_port, n282_port, n283_port, n284_port, 
      n285_port, n286_port, n287_port, n288_port, n289_port, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
      n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, 
      n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
      n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
      n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
      n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, 
      n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
      n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
      n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n_1170 : std_logic;

begin
   
   OP_COMPARE_reg_3_inst : DLH_X1 port map( G => N285, D => N289, Q => 
                           OP_COMPARE_3_port);
   OP_COMPARE_reg_2_inst : DLH_X1 port map( G => N285, D => N288, Q => 
                           OP_COMPARE_2_port);
   OP_COMPARE_reg_1_inst : DLH_X1 port map( G => N285, D => N287, Q => 
                           OP_COMPARE_1_port);
   OP_COMPARE_reg_0_inst : DLH_X1 port map( G => N285, D => N286, Q => 
                           OP_COMPARE_0_port);
   OP_A_reg_31_inst : DLH_X1 port map( G => n1411, D => OP1(31), Q => 
                           OP_A_31_port);
   OP_A_reg_30_inst : DLH_X1 port map( G => n1411, D => OP1(30), Q => 
                           OP_A_30_port);
   OP_A_reg_29_inst : DLH_X1 port map( G => n1411, D => OP1(29), Q => 
                           OP_A_29_port);
   OP_A_reg_28_inst : DLH_X1 port map( G => n1411, D => OP1(28), Q => 
                           OP_A_28_port);
   OP_A_reg_27_inst : DLH_X1 port map( G => N246, D => OP1(27), Q => 
                           OP_A_27_port);
   OP_A_reg_26_inst : DLH_X1 port map( G => N246, D => OP1(26), Q => 
                           OP_A_26_port);
   OP_A_reg_25_inst : DLH_X1 port map( G => N246, D => OP1(25), Q => 
                           OP_A_25_port);
   OP_A_reg_24_inst : DLH_X1 port map( G => n1411, D => OP1(24), Q => 
                           OP_A_24_port);
   OP_A_reg_23_inst : DLH_X1 port map( G => N246, D => OP1(23), Q => 
                           OP_A_23_port);
   OP_A_reg_22_inst : DLH_X1 port map( G => n1411, D => OP1(22), Q => 
                           OP_A_22_port);
   OP_A_reg_21_inst : DLH_X1 port map( G => n1411, D => OP1(21), Q => 
                           OP_A_21_port);
   OP_A_reg_20_inst : DLH_X1 port map( G => N246, D => OP1(20), Q => 
                           OP_A_20_port);
   OP_A_reg_19_inst : DLH_X1 port map( G => N246, D => OP1(19), Q => 
                           OP_A_19_port);
   OP_A_reg_18_inst : DLH_X1 port map( G => n1411, D => OP1(18), Q => 
                           OP_A_18_port);
   OP_A_reg_17_inst : DLH_X1 port map( G => n1411, D => OP1(17), Q => 
                           OP_A_17_port);
   OP_A_reg_16_inst : DLH_X1 port map( G => n1411, D => OP1(16), Q => 
                           OP_A_16_port);
   OP_B_reg_31_inst : DLH_X1 port map( G => N246, D => N278, Q => OP_B_31_port)
                           ;
   OP_B_reg_30_inst : DLH_X1 port map( G => n1411, D => N277, Q => OP_B_30_port
                           );
   OP_B_reg_29_inst : DLH_X1 port map( G => N246, D => N276, Q => OP_B_29_port)
                           ;
   OP_B_reg_28_inst : DLH_X1 port map( G => N246, D => N275, Q => OP_B_28_port)
                           ;
   OP_B_reg_27_inst : DLH_X1 port map( G => N246, D => N274, Q => OP_B_27_port)
                           ;
   OP_B_reg_26_inst : DLH_X1 port map( G => N246, D => N273, Q => OP_B_26_port)
                           ;
   OP_B_reg_25_inst : DLH_X1 port map( G => N246, D => N272, Q => OP_B_25_port)
                           ;
   OP_B_reg_24_inst : DLH_X1 port map( G => N246, D => N271, Q => OP_B_24_port)
                           ;
   OP_B_reg_23_inst : DLH_X1 port map( G => N246, D => N270, Q => OP_B_23_port)
                           ;
   OP_B_reg_22_inst : DLH_X1 port map( G => N246, D => N269, Q => OP_B_22_port)
                           ;
   OP_B_reg_21_inst : DLH_X1 port map( G => N246, D => N268, Q => OP_B_21_port)
                           ;
   OP_B_reg_20_inst : DLH_X1 port map( G => N246, D => N267, Q => OP_B_20_port)
                           ;
   OP_B_reg_19_inst : DLH_X1 port map( G => n1411, D => N266, Q => OP_B_19_port
                           );
   OP_B_reg_18_inst : DLH_X1 port map( G => n1411, D => N265, Q => OP_B_18_port
                           );
   OP_B_reg_17_inst : DLH_X1 port map( G => n1411, D => N264, Q => OP_B_17_port
                           );
   OP_B_reg_16_inst : DLH_X1 port map( G => n1411, D => N263, Q => OP_B_16_port
                           );
   OP_B_reg_15_inst : DLH_X1 port map( G => n1411, D => N262, Q => OP_B_15_port
                           );
   OP_B_reg_14_inst : DLH_X1 port map( G => n1411, D => N261, Q => OP_B_14_port
                           );
   OP_B_reg_13_inst : DLH_X1 port map( G => n1411, D => N260, Q => OP_B_13_port
                           );
   OP_B_reg_12_inst : DLH_X1 port map( G => n1411, D => N259, Q => OP_B_12_port
                           );
   OP_B_reg_11_inst : DLH_X1 port map( G => n1411, D => N258, Q => OP_B_11_port
                           );
   OP_B_reg_10_inst : DLH_X1 port map( G => n1411, D => N257, Q => OP_B_10_port
                           );
   OP_B_reg_9_inst : DLH_X1 port map( G => N246, D => N256, Q => OP_B_9_port);
   OP_B_reg_8_inst : DLH_X1 port map( G => N246, D => N255, Q => OP_B_8_port);
   OP_B_reg_7_inst : DLH_X1 port map( G => n1411, D => N254, Q => OP_B_7_port);
   OP_B_reg_6_inst : DLH_X1 port map( G => N246, D => N253, Q => OP_B_6_port);
   OP_B_reg_0_inst : DLH_X1 port map( G => n1411, D => N247, Q => OP_B_0_port);
   OP_Ci_reg : DLH_X1 port map( G => N279, D => N280, Q => OP_Ci);
   OP_LOGIC_reg_1_inst : DLH_X1 port map( G => N281, D => N283, Q => 
                           OP_LOGIC_1_port);
   OP_LOGIC_reg_0_inst : DLH_X1 port map( G => N281, D => N282, Q => 
                           OP_LOGIC_0_port);
   OP_SHIFT_reg : DLH_X1 port map( G => N284, D => N96, Q => OP_SHIFT);
   DP_OP_440J3_122_9847_U43 : HA_X1 port map( A => DP_OP_440J3_122_9847_n35, B 
                           => DP_OP_440J3_122_9847_n66, CO => 
                           DP_OP_440J3_122_9847_n34, S => C428_DATA4_1);
   DP_OP_440J3_122_9847_U42 : HA_X1 port map( A => DP_OP_440J3_122_9847_n34, B 
                           => DP_OP_440J3_122_9847_n67, CO => 
                           DP_OP_440J3_122_9847_n33, S => C428_DATA4_2);
   DP_OP_440J3_122_9847_U41 : HA_X1 port map( A => DP_OP_440J3_122_9847_n33, B 
                           => DP_OP_440J3_122_9847_n68, CO => 
                           DP_OP_440J3_122_9847_n32, S => C428_DATA4_3);
   DP_OP_440J3_122_9847_U40 : HA_X1 port map( A => DP_OP_440J3_122_9847_n32, B 
                           => DP_OP_440J3_122_9847_n69, CO => 
                           DP_OP_440J3_122_9847_n31, S => C428_DATA4_4);
   DP_OP_440J3_122_9847_U39 : HA_X1 port map( A => DP_OP_440J3_122_9847_n31, B 
                           => DP_OP_440J3_122_9847_n70, CO => 
                           DP_OP_440J3_122_9847_n30, S => C428_DATA4_5);
   DP_OP_440J3_122_9847_U38 : HA_X1 port map( A => DP_OP_440J3_122_9847_n30, B 
                           => DP_OP_440J3_122_9847_n71, CO => 
                           DP_OP_440J3_122_9847_n29, S => C428_DATA4_6);
   DP_OP_440J3_122_9847_U37 : HA_X1 port map( A => DP_OP_440J3_122_9847_n29, B 
                           => DP_OP_440J3_122_9847_n72, CO => 
                           DP_OP_440J3_122_9847_n28, S => C428_DATA4_7);
   DP_OP_440J3_122_9847_U36 : HA_X1 port map( A => DP_OP_440J3_122_9847_n28, B 
                           => DP_OP_440J3_122_9847_n73, CO => 
                           DP_OP_440J3_122_9847_n27, S => C428_DATA4_8);
   DP_OP_440J3_122_9847_U35 : HA_X1 port map( A => DP_OP_440J3_122_9847_n27, B 
                           => DP_OP_440J3_122_9847_n74, CO => 
                           DP_OP_440J3_122_9847_n26, S => C428_DATA4_9);
   DP_OP_440J3_122_9847_U34 : HA_X1 port map( A => DP_OP_440J3_122_9847_n26, B 
                           => DP_OP_440J3_122_9847_n75, CO => 
                           DP_OP_440J3_122_9847_n25, S => C428_DATA4_10);
   DP_OP_440J3_122_9847_U33 : HA_X1 port map( A => DP_OP_440J3_122_9847_n25, B 
                           => DP_OP_440J3_122_9847_n76, CO => 
                           DP_OP_440J3_122_9847_n24, S => C428_DATA4_11);
   DP_OP_440J3_122_9847_U32 : HA_X1 port map( A => DP_OP_440J3_122_9847_n24, B 
                           => DP_OP_440J3_122_9847_n77, CO => 
                           DP_OP_440J3_122_9847_n23, S => C428_DATA4_12);
   DP_OP_440J3_122_9847_U31 : HA_X1 port map( A => DP_OP_440J3_122_9847_n23, B 
                           => DP_OP_440J3_122_9847_n78, CO => 
                           DP_OP_440J3_122_9847_n22, S => C428_DATA4_13);
   DP_OP_440J3_122_9847_U30 : HA_X1 port map( A => DP_OP_440J3_122_9847_n22, B 
                           => DP_OP_440J3_122_9847_n79, CO => 
                           DP_OP_440J3_122_9847_n21, S => C428_DATA4_14);
   DP_OP_440J3_122_9847_U29 : HA_X1 port map( A => DP_OP_440J3_122_9847_n21, B 
                           => DP_OP_440J3_122_9847_n80, CO => 
                           DP_OP_440J3_122_9847_n20, S => C428_DATA4_15);
   DP_OP_446J3_125_4819_U33 : HA_X1 port map( A => n1413, B => 
                           DP_OP_446J3_125_4819_n72, CO => 
                           DP_OP_446J3_125_4819_n27, S => C2_DATA1_6);
   DP_OP_446J3_125_4819_U32 : HA_X1 port map( A => DP_OP_446J3_125_4819_n27, B 
                           => DP_OP_446J3_125_4819_n73, CO => 
                           DP_OP_446J3_125_4819_n26, S => C429_DATA4_7);
   DP_OP_446J3_125_4819_U31 : HA_X1 port map( A => DP_OP_446J3_125_4819_n26, B 
                           => DP_OP_446J3_125_4819_n74, CO => 
                           DP_OP_446J3_125_4819_n25, S => C429_DATA4_8);
   DP_OP_446J3_125_4819_U30 : HA_X1 port map( A => DP_OP_446J3_125_4819_n25, B 
                           => DP_OP_446J3_125_4819_n75, CO => 
                           DP_OP_446J3_125_4819_n24, S => C429_DATA4_9);
   DP_OP_446J3_125_4819_U29 : HA_X1 port map( A => DP_OP_446J3_125_4819_n24, B 
                           => DP_OP_446J3_125_4819_n76, CO => 
                           DP_OP_446J3_125_4819_n23, S => C429_DATA4_10);
   DP_OP_446J3_125_4819_U28 : HA_X1 port map( A => DP_OP_446J3_125_4819_n23, B 
                           => DP_OP_446J3_125_4819_n77, CO => 
                           DP_OP_446J3_125_4819_n22, S => C429_DATA4_11);
   DP_OP_446J3_125_4819_U27 : HA_X1 port map( A => DP_OP_446J3_125_4819_n22, B 
                           => DP_OP_446J3_125_4819_n78, CO => 
                           DP_OP_446J3_125_4819_n21, S => C429_DATA4_12);
   DP_OP_446J3_125_4819_U26 : HA_X1 port map( A => DP_OP_446J3_125_4819_n21, B 
                           => DP_OP_446J3_125_4819_n79, CO => 
                           DP_OP_446J3_125_4819_n20, S => C429_DATA4_13);
   DP_OP_446J3_125_4819_U25 : HA_X1 port map( A => DP_OP_446J3_125_4819_n20, B 
                           => DP_OP_446J3_125_4819_n80, CO => 
                           DP_OP_446J3_125_4819_n19, S => C429_DATA4_14);
   DP_OP_446J3_125_4819_U24 : HA_X1 port map( A => DP_OP_446J3_125_4819_n19, B 
                           => DP_OP_446J3_125_4819_n81, CO => 
                           DP_OP_446J3_125_4819_n18, S => C429_DATA4_15);
   DP_OP_446J3_125_4819_U23 : HA_X1 port map( A => DP_OP_446J3_125_4819_n18, B 
                           => DP_OP_446J3_125_4819_n82, CO => 
                           DP_OP_446J3_125_4819_n17, S => C429_DATA4_16);
   DP_OP_446J3_125_4819_U22 : HA_X1 port map( A => DP_OP_446J3_125_4819_n17, B 
                           => DP_OP_446J3_125_4819_n83, CO => 
                           DP_OP_446J3_125_4819_n16, S => C429_DATA4_17);
   DP_OP_446J3_125_4819_U21 : HA_X1 port map( A => DP_OP_446J3_125_4819_n16, B 
                           => DP_OP_446J3_125_4819_n84, CO => 
                           DP_OP_446J3_125_4819_n15, S => C429_DATA4_18);
   DP_OP_446J3_125_4819_U20 : HA_X1 port map( A => DP_OP_446J3_125_4819_n15, B 
                           => DP_OP_446J3_125_4819_n85, CO => 
                           DP_OP_446J3_125_4819_n14, S => C429_DATA4_19);
   DP_OP_446J3_125_4819_U19 : HA_X1 port map( A => DP_OP_446J3_125_4819_n14, B 
                           => DP_OP_446J3_125_4819_n86, CO => 
                           DP_OP_446J3_125_4819_n13, S => C429_DATA4_20);
   DP_OP_446J3_125_4819_U18 : HA_X1 port map( A => DP_OP_446J3_125_4819_n13, B 
                           => DP_OP_446J3_125_4819_n87, CO => 
                           DP_OP_446J3_125_4819_n12, S => C429_DATA4_21);
   DP_OP_451J3_128_3502_U37 : HA_X1 port map( A => n1412, B => 
                           DP_OP_451J3_128_3502_n70, CO => 
                           DP_OP_451J3_128_3502_n30, S => C2_DATA1_4);
   DP_OP_451J3_128_3502_U36 : HA_X1 port map( A => DP_OP_451J3_128_3502_n30, B 
                           => DP_OP_451J3_128_3502_n71, CO => 
                           DP_OP_451J3_128_3502_n29, S => C430_DATA4_5);
   DP_OP_451J3_128_3502_U35 : HA_X1 port map( A => DP_OP_451J3_128_3502_n29, B 
                           => DP_OP_451J3_128_3502_n72, CO => 
                           DP_OP_451J3_128_3502_n28, S => C430_DATA4_6);
   DP_OP_451J3_128_3502_U34 : HA_X1 port map( A => DP_OP_451J3_128_3502_n28, B 
                           => DP_OP_451J3_128_3502_n73, CO => 
                           DP_OP_451J3_128_3502_n27, S => C430_DATA4_7);
   DP_OP_451J3_128_3502_U33 : HA_X1 port map( A => DP_OP_451J3_128_3502_n27, B 
                           => DP_OP_451J3_128_3502_n74, CO => 
                           DP_OP_451J3_128_3502_n26, S => C430_DATA4_8);
   DP_OP_451J3_128_3502_U32 : HA_X1 port map( A => DP_OP_451J3_128_3502_n26, B 
                           => DP_OP_451J3_128_3502_n75, CO => 
                           DP_OP_451J3_128_3502_n25, S => C430_DATA4_9);
   DP_OP_451J3_128_3502_U31 : HA_X1 port map( A => DP_OP_451J3_128_3502_n25, B 
                           => DP_OP_451J3_128_3502_n76, CO => 
                           DP_OP_451J3_128_3502_n24, S => C430_DATA4_10);
   DP_OP_451J3_128_3502_U30 : HA_X1 port map( A => DP_OP_451J3_128_3502_n24, B 
                           => DP_OP_451J3_128_3502_n77, CO => 
                           DP_OP_451J3_128_3502_n23, S => C430_DATA4_11);
   DP_OP_451J3_128_3502_U29 : HA_X1 port map( A => DP_OP_451J3_128_3502_n23, B 
                           => DP_OP_451J3_128_3502_n78, CO => 
                           DP_OP_451J3_128_3502_n22, S => C430_DATA4_12);
   DP_OP_451J3_128_3502_U28 : HA_X1 port map( A => DP_OP_451J3_128_3502_n22, B 
                           => DP_OP_451J3_128_3502_n79, CO => 
                           DP_OP_451J3_128_3502_n21, S => C430_DATA4_13);
   DP_OP_451J3_128_3502_U27 : HA_X1 port map( A => DP_OP_451J3_128_3502_n21, B 
                           => DP_OP_451J3_128_3502_n80, CO => 
                           DP_OP_451J3_128_3502_n20, S => C430_DATA4_14);
   DP_OP_451J3_128_3502_U26 : HA_X1 port map( A => DP_OP_451J3_128_3502_n20, B 
                           => DP_OP_451J3_128_3502_n81, CO => 
                           DP_OP_451J3_128_3502_n19, S => C430_DATA4_15);
   DP_OP_451J3_128_3502_U25 : HA_X1 port map( A => DP_OP_451J3_128_3502_n19, B 
                           => DP_OP_451J3_128_3502_n82, CO => 
                           DP_OP_451J3_128_3502_n18, S => C430_DATA4_16);
   DP_OP_451J3_128_3502_U24 : HA_X1 port map( A => DP_OP_451J3_128_3502_n18, B 
                           => DP_OP_451J3_128_3502_n83, CO => 
                           DP_OP_451J3_128_3502_n17, S => C430_DATA4_17);
   DP_OP_451J3_128_3502_U23 : HA_X1 port map( A => DP_OP_451J3_128_3502_n17, B 
                           => DP_OP_451J3_128_3502_n84, CO => 
                           DP_OP_451J3_128_3502_n16, S => C430_DATA4_18);
   DP_OP_451J3_128_3502_U22 : HA_X1 port map( A => DP_OP_451J3_128_3502_n16, B 
                           => DP_OP_451J3_128_3502_n85, CO => 
                           DP_OP_451J3_128_3502_n15, S => C430_DATA4_19);
   DP_OP_456J3_131_2158_U40 : HA_X1 port map( A => n1414, B => 
                           DP_OP_456J3_131_2158_n67, CO => 
                           DP_OP_456J3_131_2158_n32, S => C2_DATA1_2);
   DP_OP_456J3_131_2158_U39 : HA_X1 port map( A => DP_OP_456J3_131_2158_n32, B 
                           => DP_OP_456J3_131_2158_n68, CO => 
                           DP_OP_456J3_131_2158_n31, S => C431_DATA4_3);
   DP_OP_456J3_131_2158_U38 : HA_X1 port map( A => DP_OP_456J3_131_2158_n31, B 
                           => DP_OP_456J3_131_2158_n69, CO => 
                           DP_OP_456J3_131_2158_n30, S => C431_DATA4_4);
   DP_OP_456J3_131_2158_U37 : HA_X1 port map( A => DP_OP_456J3_131_2158_n30, B 
                           => DP_OP_456J3_131_2158_n70, CO => 
                           DP_OP_456J3_131_2158_n29, S => C431_DATA4_5);
   DP_OP_456J3_131_2158_U36 : HA_X1 port map( A => DP_OP_456J3_131_2158_n29, B 
                           => DP_OP_456J3_131_2158_n71, CO => 
                           DP_OP_456J3_131_2158_n28, S => C431_DATA4_6);
   DP_OP_456J3_131_2158_U35 : HA_X1 port map( A => DP_OP_456J3_131_2158_n28, B 
                           => DP_OP_456J3_131_2158_n72, CO => 
                           DP_OP_456J3_131_2158_n27, S => C431_DATA4_7);
   DP_OP_456J3_131_2158_U34 : HA_X1 port map( A => DP_OP_456J3_131_2158_n27, B 
                           => DP_OP_456J3_131_2158_n73, CO => 
                           DP_OP_456J3_131_2158_n26, S => C431_DATA4_8);
   DP_OP_456J3_131_2158_U33 : HA_X1 port map( A => DP_OP_456J3_131_2158_n26, B 
                           => DP_OP_456J3_131_2158_n74, CO => 
                           DP_OP_456J3_131_2158_n25, S => C431_DATA4_9);
   DP_OP_456J3_131_2158_U32 : HA_X1 port map( A => DP_OP_456J3_131_2158_n25, B 
                           => DP_OP_456J3_131_2158_n75, CO => 
                           DP_OP_456J3_131_2158_n24, S => C431_DATA4_10);
   DP_OP_456J3_131_2158_U31 : HA_X1 port map( A => DP_OP_456J3_131_2158_n24, B 
                           => DP_OP_456J3_131_2158_n76, CO => 
                           DP_OP_456J3_131_2158_n23, S => C431_DATA4_11);
   DP_OP_456J3_131_2158_U30 : HA_X1 port map( A => DP_OP_456J3_131_2158_n23, B 
                           => DP_OP_456J3_131_2158_n77, CO => 
                           DP_OP_456J3_131_2158_n22, S => C431_DATA4_12);
   DP_OP_456J3_131_2158_U29 : HA_X1 port map( A => DP_OP_456J3_131_2158_n22, B 
                           => DP_OP_456J3_131_2158_n78, CO => 
                           DP_OP_456J3_131_2158_n21, S => C431_DATA4_13);
   DP_OP_456J3_131_2158_U28 : HA_X1 port map( A => DP_OP_456J3_131_2158_n21, B 
                           => DP_OP_456J3_131_2158_n79, CO => 
                           DP_OP_456J3_131_2158_n20, S => C431_DATA4_14);
   DP_OP_456J3_131_2158_U27 : HA_X1 port map( A => DP_OP_456J3_131_2158_n20, B 
                           => DP_OP_456J3_131_2158_n80, CO => 
                           DP_OP_456J3_131_2158_n19, S => C431_DATA4_15);
   DP_OP_456J3_131_2158_U26 : HA_X1 port map( A => DP_OP_456J3_131_2158_n19, B 
                           => DP_OP_456J3_131_2158_n81, CO => 
                           DP_OP_456J3_131_2158_n18, S => C431_DATA4_16);
   DP_OP_456J3_131_2158_U25 : HA_X1 port map( A => DP_OP_456J3_131_2158_n18, B 
                           => DP_OP_456J3_131_2158_n82, CO => 
                           DP_OP_456J3_131_2158_n17, S => C431_DATA4_17);
   intadd_0_U28 : FA_X1 port map( A => intadd_0_A_0_port, B => 
                           intadd_0_B_0_port, CI => intadd_0_CI, CO => 
                           intadd_0_n27, S => intadd_0_SUM_0_port);
   intadd_0_U27 : FA_X1 port map( A => intadd_0_A_1_port, B => 
                           intadd_0_B_1_port, CI => intadd_0_n27, CO => 
                           intadd_0_n26, S => intadd_0_SUM_1_port);
   intadd_0_U26 : FA_X1 port map( A => intadd_0_A_2_port, B => 
                           intadd_0_B_2_port, CI => intadd_0_n26, CO => 
                           intadd_0_n25, S => intadd_0_SUM_2_port);
   intadd_0_U25 : FA_X1 port map( A => intadd_0_A_3_port, B => 
                           intadd_0_B_3_port, CI => intadd_0_n25, CO => 
                           intadd_0_n24, S => intadd_0_SUM_3_port);
   intadd_0_U24 : FA_X1 port map( A => intadd_0_A_4_port, B => 
                           intadd_0_B_4_port, CI => intadd_0_n24, CO => 
                           intadd_0_n23, S => intadd_0_SUM_4_port);
   intadd_0_U23 : FA_X1 port map( A => intadd_0_A_5_port, B => 
                           intadd_0_B_5_port, CI => intadd_0_n23, CO => 
                           intadd_0_n22, S => intadd_0_SUM_5_port);
   intadd_0_U22 : FA_X1 port map( A => intadd_0_A_6_port, B => 
                           intadd_0_B_6_port, CI => intadd_0_n22, CO => 
                           intadd_0_n21, S => intadd_0_SUM_6_port);
   intadd_0_U21 : FA_X1 port map( A => intadd_0_A_7_port, B => 
                           intadd_0_B_7_port, CI => intadd_0_n21, CO => 
                           intadd_0_n20, S => intadd_0_SUM_7_port);
   intadd_0_U20 : FA_X1 port map( A => intadd_0_A_8_port, B => 
                           intadd_0_B_8_port, CI => intadd_0_n20, CO => 
                           intadd_0_n19, S => intadd_0_SUM_8_port);
   intadd_0_U19 : FA_X1 port map( A => intadd_0_A_9_port, B => 
                           intadd_0_B_9_port, CI => intadd_0_n19, CO => 
                           intadd_0_n18, S => intadd_0_SUM_9_port);
   intadd_0_U18 : FA_X1 port map( A => intadd_0_A_10_port, B => 
                           intadd_0_B_10_port, CI => intadd_0_n18, CO => 
                           intadd_0_n17, S => intadd_0_SUM_10_port);
   intadd_0_U17 : FA_X1 port map( A => intadd_0_A_11_port, B => 
                           intadd_0_B_11_port, CI => intadd_0_n17, CO => 
                           intadd_0_n16, S => intadd_0_SUM_11_port);
   intadd_0_U16 : FA_X1 port map( A => intadd_0_A_12_port, B => 
                           intadd_0_B_12_port, CI => intadd_0_n16, CO => 
                           intadd_0_n15, S => intadd_0_SUM_12_port);
   intadd_0_U15 : FA_X1 port map( A => intadd_0_A_16_port, B => 
                           intadd_0_B_13_port, CI => intadd_0_n15, CO => 
                           intadd_0_n14, S => intadd_0_SUM_13_port);
   intadd_0_U14 : FA_X1 port map( A => intadd_0_A_16_port, B => 
                           intadd_0_B_14_port, CI => intadd_0_n14, CO => 
                           intadd_0_n13, S => intadd_0_SUM_14_port);
   intadd_0_U13 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n13, CO => intadd_0_n12, S => 
                           intadd_0_SUM_15_port);
   intadd_0_U12 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n12, CO => intadd_0_n11, S => 
                           intadd_0_SUM_16_port);
   intadd_0_U11 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n11, CO => intadd_0_n10, S => 
                           intadd_0_SUM_17_port);
   intadd_0_U10 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n10, CO => intadd_0_n9, S => 
                           intadd_0_SUM_18_port);
   intadd_0_U9 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n9, CO => intadd_0_n8, S => 
                           intadd_0_SUM_19_port);
   intadd_0_U8 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n8, CO => intadd_0_n7, S => 
                           intadd_0_SUM_20_port);
   intadd_0_U7 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n7, CO => intadd_0_n6, S => 
                           intadd_0_SUM_21_port);
   intadd_0_U6 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n6, CO => intadd_0_n5, S => 
                           intadd_0_SUM_22_port);
   intadd_0_U5 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n5, CO => intadd_0_n4, S => 
                           intadd_0_SUM_23_port);
   intadd_0_U4 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n4, CO => intadd_0_n3, S => 
                           intadd_0_SUM_24_port);
   intadd_0_U3 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n3, CO => intadd_0_n2, S => 
                           intadd_0_SUM_25_port);
   intadd_0_U2 : FA_X1 port map( A => intadd_0_A_16_port, B => n64, CI => 
                           intadd_0_n2, CO => intadd_0_n1, S => 
                           intadd_0_SUM_26_port);
   intadd_1_U26 : FA_X1 port map( A => intadd_1_A_0_port, B => 
                           intadd_1_B_0_port, CI => intadd_0_SUM_2_port, CO => 
                           intadd_1_n25, S => intadd_1_SUM_0_port);
   intadd_1_U25 : FA_X1 port map( A => intadd_0_SUM_3_port, B => 
                           intadd_1_B_1_port, CI => intadd_1_n25, CO => 
                           intadd_1_n24, S => intadd_1_SUM_1_port);
   intadd_1_U24 : FA_X1 port map( A => intadd_0_SUM_4_port, B => 
                           intadd_1_B_2_port, CI => intadd_1_n24, CO => 
                           intadd_1_n23, S => intadd_1_SUM_2_port);
   intadd_1_U23 : FA_X1 port map( A => intadd_0_SUM_5_port, B => 
                           intadd_1_B_3_port, CI => intadd_1_n23, CO => 
                           intadd_1_n22, S => intadd_1_SUM_3_port);
   intadd_1_U22 : FA_X1 port map( A => intadd_0_SUM_6_port, B => 
                           intadd_1_B_4_port, CI => intadd_1_n22, CO => 
                           intadd_1_n21, S => intadd_1_SUM_4_port);
   intadd_1_U21 : FA_X1 port map( A => intadd_0_SUM_7_port, B => 
                           intadd_1_B_5_port, CI => intadd_1_n21, CO => 
                           intadd_1_n20, S => intadd_1_SUM_5_port);
   intadd_1_U20 : FA_X1 port map( A => intadd_0_SUM_8_port, B => 
                           intadd_1_B_6_port, CI => intadd_1_n20, CO => 
                           intadd_1_n19, S => intadd_1_SUM_6_port);
   intadd_1_U19 : FA_X1 port map( A => intadd_0_SUM_9_port, B => 
                           intadd_1_B_7_port, CI => intadd_1_n19, CO => 
                           intadd_1_n18, S => intadd_1_SUM_7_port);
   intadd_1_U18 : FA_X1 port map( A => intadd_0_SUM_10_port, B => 
                           intadd_1_B_8_port, CI => intadd_1_n18, CO => 
                           intadd_1_n17, S => intadd_1_SUM_8_port);
   intadd_1_U17 : FA_X1 port map( A => intadd_0_SUM_11_port, B => 
                           intadd_1_B_9_port, CI => intadd_1_n17, CO => 
                           intadd_1_n16, S => intadd_1_SUM_9_port);
   intadd_1_U16 : FA_X1 port map( A => intadd_0_SUM_12_port, B => 
                           intadd_1_B_10_port, CI => intadd_1_n16, CO => 
                           intadd_1_n15, S => intadd_1_SUM_10_port);
   intadd_1_U15 : FA_X1 port map( A => intadd_0_SUM_13_port, B => 
                           intadd_1_B_11_port, CI => intadd_1_n15, CO => 
                           intadd_1_n14, S => intadd_1_SUM_11_port);
   intadd_1_U14 : FA_X1 port map( A => intadd_0_SUM_14_port, B => 
                           intadd_1_B_12_port, CI => intadd_1_n14, CO => 
                           intadd_1_n13, S => intadd_1_SUM_12_port);
   intadd_1_U13 : FA_X1 port map( A => intadd_0_SUM_15_port, B => 
                           intadd_1_B_13_port, CI => intadd_1_n13, CO => 
                           intadd_1_n12, S => intadd_1_SUM_13_port);
   intadd_1_U12 : FA_X1 port map( A => intadd_0_SUM_16_port, B => 
                           intadd_1_B_14_port, CI => intadd_1_n12, CO => 
                           intadd_1_n11, S => intadd_1_SUM_14_port);
   intadd_1_U11 : FA_X1 port map( A => intadd_0_SUM_17_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n11, CO => 
                           intadd_1_n10, S => intadd_1_SUM_15_port);
   intadd_1_U10 : FA_X1 port map( A => intadd_0_SUM_18_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n10, CO => 
                           intadd_1_n9, S => intadd_1_SUM_16_port);
   intadd_1_U9 : FA_X1 port map( A => intadd_0_SUM_19_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n9, CO => 
                           intadd_1_n8, S => intadd_1_SUM_17_port);
   intadd_1_U8 : FA_X1 port map( A => intadd_0_SUM_20_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n8, CO => 
                           intadd_1_n7, S => intadd_1_SUM_18_port);
   intadd_1_U7 : FA_X1 port map( A => intadd_0_SUM_21_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n7, CO => 
                           intadd_1_n6, S => intadd_1_SUM_19_port);
   intadd_1_U6 : FA_X1 port map( A => intadd_0_SUM_22_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n6, CO => 
                           intadd_1_n5, S => intadd_1_SUM_20_port);
   intadd_1_U5 : FA_X1 port map( A => intadd_0_SUM_23_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n5, CO => 
                           intadd_1_n4, S => intadd_1_SUM_21_port);
   intadd_1_U4 : FA_X1 port map( A => intadd_0_SUM_24_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n4, CO => 
                           intadd_1_n3, S => intadd_1_SUM_22_port);
   intadd_1_U3 : FA_X1 port map( A => intadd_0_SUM_25_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n3, CO => 
                           intadd_1_n2, S => intadd_1_SUM_23_port);
   intadd_1_U2 : FA_X1 port map( A => intadd_0_SUM_26_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n2, CO => 
                           intadd_1_n1, S => intadd_1_SUM_24_port);
   intadd_2_U11 : FA_X1 port map( A => intadd_2_A_0_port, B => 
                           intadd_2_B_0_port, CI => intadd_1_SUM_2_port, CO => 
                           intadd_2_n10, S => intadd_2_SUM_0_port);
   intadd_2_U10 : FA_X1 port map( A => intadd_2_A_1_port, B => 
                           intadd_1_SUM_3_port, CI => intadd_2_n10, CO => 
                           intadd_2_n9, S => intadd_2_SUM_1_port);
   intadd_2_U9 : FA_X1 port map( A => intadd_2_A_2_port, B => 
                           intadd_1_SUM_4_port, CI => intadd_2_n9, CO => 
                           intadd_2_n8, S => intadd_2_SUM_2_port);
   intadd_2_U8 : FA_X1 port map( A => intadd_2_A_3_port, B => 
                           intadd_1_SUM_5_port, CI => intadd_2_n8, CO => 
                           intadd_2_n7, S => intadd_2_SUM_3_port);
   intadd_2_U7 : FA_X1 port map( A => intadd_2_A_4_port, B => 
                           intadd_1_SUM_6_port, CI => intadd_2_n7, CO => 
                           intadd_2_n6, S => intadd_2_SUM_4_port);
   intadd_2_U6 : FA_X1 port map( A => intadd_2_A_5_port, B => 
                           intadd_1_SUM_7_port, CI => intadd_2_n6, CO => 
                           intadd_2_n5, S => intadd_2_SUM_5_port);
   intadd_2_U5 : FA_X1 port map( A => intadd_2_A_6_port, B => 
                           intadd_1_SUM_8_port, CI => intadd_2_n5, CO => 
                           intadd_2_n4, S => intadd_2_SUM_6_port);
   intadd_2_U4 : FA_X1 port map( A => intadd_2_A_7_port, B => 
                           intadd_1_SUM_9_port, CI => intadd_2_n4, CO => 
                           intadd_2_n3, S => intadd_2_SUM_7_port);
   intadd_2_U3 : FA_X1 port map( A => intadd_2_A_8_port, B => 
                           intadd_1_SUM_10_port, CI => intadd_2_n3, CO => 
                           intadd_2_n2, S => intadd_2_SUM_8_port);
   intadd_2_U2 : FA_X1 port map( A => intadd_2_A_9_port, B => 
                           intadd_1_SUM_11_port, CI => intadd_2_n2, CO => 
                           intadd_2_n1, S => intadd_2_SUM_9_port);
   OP_A_reg_7_inst : DLH_X1 port map( G => N246, D => OP1(7), Q => OP_A_7_port)
                           ;
   OP_A_reg_12_inst : DLH_X1 port map( G => N246, D => OP1(12), Q => 
                           OP_A_12_port);
   OP_A_reg_13_inst : DLH_X1 port map( G => n1411, D => OP1(13), Q => 
                           OP_A_13_port);
   OP_A_reg_10_inst : DLH_X1 port map( G => n1411, D => OP1(10), Q => 
                           OP_A_10_port);
   OP_A_reg_0_inst : DLH_X1 port map( G => n1411, D => OP1(0), Q => OP_A_0_port
                           );
   OP_A_reg_4_inst : DLH_X1 port map( G => N246, D => OP1(4), Q => OP_A_4_port)
                           ;
   OP_A_reg_8_inst : DLH_X1 port map( G => n1411, D => OP1(8), Q => OP_A_8_port
                           );
   OP_A_reg_6_inst : DLH_X1 port map( G => N246, D => OP1(6), Q => OP_A_6_port)
                           ;
   OP_A_reg_11_inst : DLH_X1 port map( G => n1411, D => OP1(11), Q => 
                           OP_A_11_port);
   OP_A_reg_14_inst : DLH_X1 port map( G => n1411, D => OP1(14), Q => 
                           OP_A_14_port);
   OP_A_reg_1_inst : DLH_X1 port map( G => N246, D => OP1(1), Q => OP_A_1_port)
                           ;
   OP_A_reg_3_inst : DLH_X1 port map( G => N246, D => OP1(3), Q => OP_A_3_port)
                           ;
   OP_A_reg_9_inst : DLH_X1 port map( G => n1411, D => OP1(9), Q => OP_A_9_port
                           );
   OP_A_reg_5_inst : DLH_X1 port map( G => n1411, D => OP1(5), Q => OP_A_5_port
                           );
   OP_B_reg_2_inst : DLH_X1 port map( G => N246, D => N249, Q => OP_B_2_port);
   OP_B_reg_5_inst : DLH_X1 port map( G => n1411, D => N252, Q => OP_B_5_port);
   OP_B_reg_3_inst : DLH_X1 port map( G => N246, D => N250, Q => OP_B_3_port);
   OP_A_reg_15_inst : DLH_X1 port map( G => n1411, D => OP1(15), Q => 
                           OP_A_15_port);
   OP_B_reg_4_inst : DLH_X1 port map( G => N246, D => N251, Q => OP_B_4_port);
   OP_A_reg_2_inst : DLH_X1 port map( G => N246, D => OP1(2), Q => OP_A_2_port)
                           ;
   OP_B_reg_1_inst : DLH_X2 port map( G => N246, D => N248, Q => OP_B_1_port);
   U3 : CLKBUF_X1 port map( A => n150, Z => n62);
   U4 : CLKBUF_X2 port map( A => n196, Z => n58);
   U5 : INV_X1 port map( A => n1367, ZN => n1366);
   U6 : INV_X2 port map( A => n577, ZN => n55);
   U7 : INV_X2 port map( A => n510, ZN => n56);
   U8 : INV_X2 port map( A => n607, ZN => n57);
   U9 : INV_X2 port map( A => N280, ZN => n198);
   U10 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_15, B1 => 
                           OP_A_11_port, B2 => n161, C1 => n162, C2 => 
                           OP_A_10_port, ZN => intadd_1_B_9_port);
   U11 : AOI211_X1 port map( C1 => n66, C2 => n863, A => n541, B => n540, ZN =>
                           n964);
   U12 : NOR2_X2 port map( A1 => DP_OP_446J3_125_4819_n12, A2 => n1091, ZN => 
                           n59);
   U13 : OR2_X1 port map( A1 => n147, A2 => n114, ZN => n60);
   U14 : OR3_X1 port map( A1 => n1081, A2 => OP_B_7_port, A3 => n163, ZN => n61
                           );
   U15 : NOR2_X2 port map( A1 => OP_B_2_port, A2 => n1159, ZN => n855);
   U16 : NOR2_X2 port map( A1 => OP_B_7_port, A2 => n164, ZN => n1027);
   U17 : NOR2_X2 port map( A1 => n225, A2 => n742, ZN => n149);
   U18 : NOR2_X2 port map( A1 => OP_B_5_port, A2 => n156, ZN => n162);
   U19 : AOI21_X2 port map( B1 => OP_B_3_port, B2 => OP_B_4_port, A => n298, ZN
                           => n1412);
   U20 : NOR2_X2 port map( A1 => OP_B_3_port, A2 => OP_B_2_port, ZN => n894);
   U21 : INV_X1 port map( A => n61, ZN => n63);
   U22 : INV_X1 port map( A => n60, ZN => n64);
   U23 : NOR2_X2 port map( A1 => n900, A2 => n1260, ZN => n1227);
   U24 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n581, ZN => n65);
   U25 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n581, ZN => n66);
   U26 : NOR2_X2 port map( A1 => n1380, A2 => n116, ZN => intadd_1_B_18_port);
   U27 : AOI21_X2 port map( B1 => OP_B_2_port, B2 => OP_B_1_port, A => n1159, 
                           ZN => n1414);
   U28 : NOR3_X4 port map( A1 => n152, A2 => OP_B_5_port, A3 => n155, ZN => 
                           n161);
   U29 : NOR2_X4 port map( A1 => n128, A2 => n111, ZN => intadd_0_A_16_port);
   U30 : NOR3_X4 port map( A1 => n1081, A2 => OP_B_7_port, A3 => n1080, ZN => 
                           n1379);
   U31 : OR2_X1 port map( A1 => n1412, A2 => n1380, ZN => n67);
   U32 : INV_X1 port map( A => OPC(4), ZN => n71);
   U33 : NOR3_X1 port map( A1 => N284, A2 => N285, A3 => n109, ZN => n196);
   U34 : INV_X1 port map( A => OPC(6), ZN => n173);
   U35 : NOR3_X1 port map( A1 => OPC(5), A2 => n71, A3 => n173, ZN => n82);
   U36 : NAND2_X1 port map( A1 => OPC(4), A2 => OPC(5), ZN => n83);
   U37 : NOR2_X1 port map( A1 => OPC(6), A2 => n83, ZN => n79);
   U38 : NOR2_X1 port map( A1 => n82, A2 => n79, ZN => n178);
   U39 : NOR2_X1 port map( A1 => OPC(2), A2 => OPC(1), ZN => n74);
   U40 : INV_X1 port map( A => OPC(3), ZN => n68);
   U41 : INV_X1 port map( A => OPC(0), ZN => n69);
   U42 : NAND3_X1 port map( A1 => n74, A2 => n68, A3 => n69, ZN => n98);
   U43 : INV_X1 port map( A => OPC(5), ZN => n70);
   U44 : NAND2_X1 port map( A1 => n71, A2 => n70, ZN => n217);
   U45 : NOR2_X1 port map( A1 => OPC(3), A2 => n69, ZN => n85);
   U46 : NAND2_X1 port map( A1 => n74, A2 => n85, ZN => n1410);
   U47 : OAI22_X1 port map( A1 => n178, A2 => n98, B1 => n217, B2 => n1410, ZN 
                           => N280);
   U48 : NOR2_X1 port map( A1 => OPC(4), A2 => n70, ZN => n90);
   U49 : NAND2_X1 port map( A1 => n90, A2 => n173, ZN => n174);
   U50 : NOR3_X1 port map( A1 => OPC(6), A2 => OPC(5), A3 => n71, ZN => n102);
   U51 : INV_X1 port map( A => n102, ZN => n1409);
   U52 : NAND3_X1 port map( A1 => OPC(3), A2 => OPC(0), A3 => n74, ZN => n216);
   U53 : OAI22_X1 port map( A1 => n174, A2 => n98, B1 => n1409, B2 => n216, ZN 
                           => N96);
   U54 : NAND3_X1 port map( A1 => OPC(6), A2 => OPC(5), A3 => n71, ZN => n1405)
                           ;
   U55 : INV_X1 port map( A => n98, ZN => n104);
   U56 : INV_X1 port map( A => n217, ZN => n103);
   U57 : NAND2_X1 port map( A1 => OPC(6), A2 => n103, ZN => n1408);
   U58 : INV_X1 port map( A => n1408, ZN => n72);
   U59 : AOI21_X1 port map( B1 => n104, B2 => n72, A => N96, ZN => n73);
   U60 : OAI21_X1 port map( B1 => n1405, B2 => n216, A => n73, ZN => N284);
   U61 : NAND2_X1 port map( A1 => OPC(3), A2 => n74, ZN => n75);
   U62 : NOR2_X1 port map( A1 => OPC(0), A2 => n75, ZN => n88);
   U63 : INV_X1 port map( A => n88, ZN => n1407);
   U64 : INV_X1 port map( A => n216, ZN => n80);
   U65 : NAND2_X1 port map( A1 => OPC(2), A2 => OPC(3), ZN => n76);
   U66 : NOR2_X1 port map( A1 => OPC(0), A2 => n76, ZN => n96_port);
   U67 : INV_X1 port map( A => OPC(1), ZN => n106);
   U68 : INV_X1 port map( A => OPC(2), ZN => n77);
   U69 : NAND3_X1 port map( A1 => OPC(1), A2 => n85, A3 => n77, ZN => n95);
   U70 : INV_X1 port map( A => n95, ZN => n78);
   U71 : AOI21_X1 port map( B1 => n96_port, B2 => n106, A => n78, ZN => n181);
   U72 : NOR2_X1 port map( A1 => OPC(4), A2 => n181, ZN => n171);
   U73 : AOI21_X1 port map( B1 => n80, B2 => n79, A => n171, ZN => n81);
   U74 : OAI21_X1 port map( B1 => n1405, B2 => n1407, A => n81, ZN => N286);
   U75 : INV_X1 port map( A => n82, ZN => n218);
   U76 : AOI21_X1 port map( B1 => n174, B2 => n218, A => n1407, ZN => n86);
   U77 : NAND2_X1 port map( A1 => OPC(4), A2 => n173, ZN => n84);
   U78 : OR2_X1 port map( A1 => n173, A2 => n83, ZN => n92);
   U79 : OAI22_X1 port map( A1 => n84, A2 => n1407, B1 => n216, B2 => n92, ZN 
                           => n170);
   U80 : NAND3_X1 port map( A1 => OPC(2), A2 => n85, A3 => n106, ZN => n94);
   U81 : OAI22_X1 port map( A1 => n174, A2 => n94, B1 => n1407, B2 => n92, ZN 
                           => n179);
   U82 : NOR4_X1 port map( A1 => n86, A2 => n170, A3 => N286, A4 => n179, ZN =>
                           n87);
   U83 : OR2_X1 port map( A1 => n217, A2 => n94, ZN => n176);
   U84 : OAI211_X1 port map( C1 => n216, C2 => n218, A => n87, B => n176, ZN =>
                           N285);
   U85 : NAND2_X1 port map( A1 => n103, A2 => n88, ZN => n1406);
   U86 : INV_X1 port map( A => n1410, ZN => n89);
   U87 : OAI21_X1 port map( B1 => n90, B2 => n102, A => n89, ZN => n91);
   U88 : OAI211_X1 port map( C1 => n98, C2 => n92, A => n1406, B => n91, ZN => 
                           N281);
   U89 : NAND3_X1 port map( A1 => OPC(2), A2 => OPC(3), A3 => OPC(0), ZN => n93
                           );
   U90 : OAI211_X1 port map( C1 => OPC(1), C2 => n93, A => n95, B => n98, ZN =>
                           n101);
   U91 : AOI21_X1 port map( B1 => n95, B2 => n94, A => n218, ZN => n100);
   U92 : NAND3_X1 port map( A1 => OPC(5), A2 => OPC(1), A3 => n96_port, ZN => 
                           n97);
   U93 : OAI21_X1 port map( B1 => n98, B2 => n1405, A => n97, ZN => n99);
   U94 : AOI211_X1 port map( C1 => n102, C2 => n101, A => n100, B => n99, ZN =>
                           n117);
   U95 : INV_X1 port map( A => N281, ZN => n220);
   U96 : NAND3_X1 port map( A1 => n104, A2 => n103, A3 => n173, ZN => n105);
   U97 : OAI21_X1 port map( B1 => n216, B2 => n174, A => n105, ZN => n1365);
   U98 : INV_X1 port map( A => n1365, ZN => n900);
   U99 : INV_X1 port map( A => n174, ZN => n108);
   U100 : AOI211_X1 port map( C1 => OPC(3), C2 => OPC(2), A => OPC(0), B => 
                           n106, ZN => n107);
   U101 : OAI211_X1 port map( C1 => OPC(2), C2 => OPC(3), A => n108, B => n107,
                           ZN => n1395);
   U102 : NAND4_X1 port map( A1 => n117, A2 => n220, A3 => n900, A4 => n1395, 
                           ZN => n109);
   U103 : NAND2_X1 port map( A1 => n198, A2 => n58, ZN => N246);
   U104 : CLKBUF_X1 port map( A => N246, Z => n1411);
   U105 : INV_X1 port map( A => OP_A_15_port, ZN => n1080);
   U106 : INV_X1 port map( A => OP_B_1_port, ZN => n225);
   U107 : INV_X1 port map( A => OP_B_0_port, ZN => n224);
   U108 : OR2_X1 port map( A1 => OP_B_1_port, A2 => n224, ZN => n510);
   U109 : NOR2_X1 port map( A1 => n1080, A2 => n510, ZN => n128);
   U110 : NOR2_X1 port map( A1 => OP_B_0_port, A2 => n225, ZN => n603);
   U111 : INV_X1 port map( A => n603, ZN => n575);
   U112 : OR2_X1 port map( A1 => n225, A2 => n224, ZN => n577);
   U113 : NAND2_X1 port map( A1 => n55, A2 => n1080, ZN => n118);
   U114 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n575, A => n118, ZN => 
                           n110);
   U115 : INV_X1 port map( A => n110, ZN => n125);
   U116 : NOR2_X1 port map( A1 => DP_OP_440J3_122_9847_n20, A2 => n125, ZN => 
                           n111);
   U117 : INV_X1 port map( A => OP_B_2_port, ZN => n581);
   U118 : AOI211_X1 port map( C1 => n581, C2 => n225, A => OP_B_3_port, B => 
                           n1080, ZN => n147);
   U119 : INV_X1 port map( A => OP_B_3_port, ZN => n1159);
   U120 : NAND2_X1 port map( A1 => n855, A2 => n225, ZN => n120);
   U121 : NAND2_X1 port map( A1 => OP_B_3_port, A2 => OP_B_2_port, ZN => n857);
   U122 : NAND2_X1 port map( A1 => OP_B_1_port, A2 => n855, ZN => n112);
   U123 : OAI21_X1 port map( B1 => OP_B_1_port, B2 => n857, A => n112, ZN => 
                           n139);
   U124 : NAND2_X1 port map( A1 => n1080, A2 => n139, ZN => n119);
   U125 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n120, A => n119, ZN => 
                           n113);
   U126 : INV_X1 port map( A => n113, ZN => n144);
   U127 : NOR2_X1 port map( A1 => DP_OP_456J3_131_2158_n17, A2 => n144, ZN => 
                           n114);
   U128 : INV_X1 port map( A => OP_B_7_port, ZN => n296);
   U129 : AOI21_X1 port map( B1 => OP_B_6_port, B2 => OP_B_5_port, A => n296, 
                           ZN => n1413);
   U130 : INV_X1 port map( A => OP_B_5_port, ZN => n298);
   U131 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => OP_B_3_port, ZN => n152);
   U132 : NOR3_X1 port map( A1 => n152, A2 => OP_B_5_port, A3 => n1080, ZN => 
                           n1380);
   U133 : NAND2_X1 port map( A1 => n152, A2 => OP_B_5_port, ZN => n123);
   U134 : INV_X1 port map( A => OP_B_4_port, ZN => n1362);
   U135 : NOR2_X1 port map( A1 => n1159, A2 => n1362, ZN => n155);
   U136 : NOR3_X1 port map( A1 => n152, A2 => n155, A3 => n298, ZN => n153);
   U137 : NAND2_X1 port map( A1 => n153, A2 => n1080, ZN => n122);
   U138 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n123, A => n122, ZN => 
                           n115);
   U139 : INV_X1 port map( A => n115, ZN => n159);
   U140 : OR2_X1 port map( A1 => DP_OP_451J3_128_3502_n15, A2 => n159, ZN => 
                           n1382);
   U141 : INV_X1 port map( A => n1382, ZN => n116);
   U142 : NAND2_X1 port map( A1 => n198, A2 => n117, ZN => N279);
   U143 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n575, A => n118, ZN => 
                           DP_OP_440J3_122_9847_n80);
   U144 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n577, B1 => OP_A_13_port
                           , B2 => n575, ZN => DP_OP_440J3_122_9847_n79);
   U145 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n577, B1 => OP_A_12_port
                           , B2 => n575, ZN => DP_OP_440J3_122_9847_n78);
   U146 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n575, B1 => OP_A_12_port
                           , B2 => n577, ZN => DP_OP_440J3_122_9847_n77);
   U147 : OAI22_X1 port map( A1 => OP_A_10_port, A2 => n575, B1 => OP_A_11_port
                           , B2 => n577, ZN => DP_OP_440J3_122_9847_n76);
   U148 : OAI22_X1 port map( A1 => OP_A_9_port, A2 => n575, B1 => OP_A_10_port,
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n75);
   U149 : OAI22_X1 port map( A1 => OP_A_8_port, A2 => n575, B1 => OP_A_9_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n74);
   U150 : OAI22_X1 port map( A1 => OP_A_7_port, A2 => n575, B1 => OP_A_8_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n73);
   U151 : OAI22_X1 port map( A1 => OP_A_6_port, A2 => n575, B1 => OP_A_7_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n72);
   U152 : OAI22_X1 port map( A1 => OP_A_5_port, A2 => n575, B1 => OP_A_6_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n71);
   U153 : OAI22_X1 port map( A1 => OP_A_4_port, A2 => n575, B1 => OP_A_5_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n70);
   U154 : OAI22_X1 port map( A1 => OP_A_3_port, A2 => n575, B1 => OP_A_4_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n69);
   U155 : OAI22_X1 port map( A1 => OP_A_2_port, A2 => n575, B1 => OP_A_3_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n68);
   U156 : OAI22_X1 port map( A1 => OP_A_2_port, A2 => n577, B1 => OP_A_1_port, 
                           B2 => n575, ZN => DP_OP_440J3_122_9847_n67);
   U157 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n577, B1 => OP_A_0_port, 
                           B2 => n575, ZN => DP_OP_440J3_122_9847_n66);
   U158 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n577, A => n575, ZN => 
                           DP_OP_440J3_122_9847_n35);
   U159 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n120, A => n119, ZN => 
                           DP_OP_456J3_131_2158_n82);
   U160 : INV_X1 port map( A => n139, ZN => n121);
   U161 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n121, B1 => OP_A_13_port
                           , B2 => n120, ZN => DP_OP_456J3_131_2158_n81);
   U162 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n121, B1 => OP_A_12_port
                           , B2 => n120, ZN => DP_OP_456J3_131_2158_n80);
   U163 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n120, B1 => OP_A_12_port
                           , B2 => n121, ZN => DP_OP_456J3_131_2158_n79);
   U164 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n121, B1 => OP_A_10_port
                           , B2 => n120, ZN => DP_OP_456J3_131_2158_n78);
   U165 : OAI22_X1 port map( A1 => n121, A2 => OP_A_10_port, B1 => OP_A_9_port,
                           B2 => n120, ZN => DP_OP_456J3_131_2158_n77);
   U166 : OAI22_X1 port map( A1 => n121, A2 => OP_A_9_port, B1 => OP_A_8_port, 
                           B2 => n120, ZN => DP_OP_456J3_131_2158_n76);
   U167 : OAI22_X1 port map( A1 => n121, A2 => OP_A_8_port, B1 => OP_A_7_port, 
                           B2 => n120, ZN => DP_OP_456J3_131_2158_n75);
   U168 : OAI22_X1 port map( A1 => n121, A2 => OP_A_7_port, B1 => OP_A_6_port, 
                           B2 => n120, ZN => DP_OP_456J3_131_2158_n74);
   U169 : OAI22_X1 port map( A1 => n121, A2 => OP_A_6_port, B1 => OP_A_5_port, 
                           B2 => n120, ZN => DP_OP_456J3_131_2158_n73);
   U170 : OAI22_X1 port map( A1 => n121, A2 => OP_A_5_port, B1 => OP_A_4_port, 
                           B2 => n120, ZN => DP_OP_456J3_131_2158_n72);
   U171 : OAI22_X1 port map( A1 => n121, A2 => OP_A_4_port, B1 => OP_A_3_port, 
                           B2 => n120, ZN => DP_OP_456J3_131_2158_n71);
   U172 : OAI22_X1 port map( A1 => n121, A2 => OP_A_3_port, B1 => OP_A_2_port, 
                           B2 => n120, ZN => DP_OP_456J3_131_2158_n70);
   U173 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n120, B1 => n121, B2 => 
                           OP_A_2_port, ZN => DP_OP_456J3_131_2158_n69);
   U174 : OAI22_X1 port map( A1 => n121, A2 => OP_A_1_port, B1 => OP_A_0_port, 
                           B2 => n120, ZN => DP_OP_456J3_131_2158_n68);
   U175 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n121, A => n120, ZN => 
                           DP_OP_456J3_131_2158_n67);
   U176 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n123, A => n122, ZN => 
                           DP_OP_451J3_128_3502_n85);
   U177 : INV_X1 port map( A => n153, ZN => n124);
   U178 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n124, B1 => OP_A_13_port
                           , B2 => n123, ZN => DP_OP_451J3_128_3502_n84);
   U179 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n124, B1 => OP_A_12_port
                           , B2 => n123, ZN => DP_OP_451J3_128_3502_n83);
   U180 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n123, B1 => OP_A_12_port
                           , B2 => n124, ZN => DP_OP_451J3_128_3502_n82);
   U181 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n124, B1 => OP_A_10_port
                           , B2 => n123, ZN => DP_OP_451J3_128_3502_n81);
   U182 : OAI22_X1 port map( A1 => OP_A_10_port, A2 => n124, B1 => OP_A_9_port,
                           B2 => n123, ZN => DP_OP_451J3_128_3502_n80);
   U183 : OAI22_X1 port map( A1 => OP_A_9_port, A2 => n124, B1 => OP_A_8_port, 
                           B2 => n123, ZN => DP_OP_451J3_128_3502_n79);
   U184 : OAI22_X1 port map( A1 => OP_A_8_port, A2 => n124, B1 => OP_A_7_port, 
                           B2 => n123, ZN => DP_OP_451J3_128_3502_n78);
   U185 : OAI22_X1 port map( A1 => OP_A_7_port, A2 => n124, B1 => OP_A_6_port, 
                           B2 => n123, ZN => DP_OP_451J3_128_3502_n77);
   U186 : OAI22_X1 port map( A1 => OP_A_6_port, A2 => n124, B1 => OP_A_5_port, 
                           B2 => n123, ZN => DP_OP_451J3_128_3502_n76);
   U187 : OAI22_X1 port map( A1 => OP_A_5_port, A2 => n124, B1 => OP_A_4_port, 
                           B2 => n123, ZN => DP_OP_451J3_128_3502_n75);
   U188 : OAI22_X1 port map( A1 => OP_A_4_port, A2 => n124, B1 => OP_A_3_port, 
                           B2 => n123, ZN => DP_OP_451J3_128_3502_n74);
   U189 : OAI22_X1 port map( A1 => OP_A_3_port, A2 => n124, B1 => OP_A_2_port, 
                           B2 => n123, ZN => DP_OP_451J3_128_3502_n73);
   U190 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n123, B1 => OP_A_2_port, 
                           B2 => n124, ZN => DP_OP_451J3_128_3502_n72);
   U191 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n124, B1 => OP_A_0_port, 
                           B2 => n123, ZN => DP_OP_451J3_128_3502_n71);
   U192 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n124, A => n123, ZN => 
                           DP_OP_451J3_128_3502_n70);
   U193 : XNOR2_X1 port map( A => DP_OP_440J3_122_9847_n20, B => n125, ZN => 
                           n126);
   U194 : INV_X1 port map( A => n128, ZN => n890);
   U195 : NAND2_X1 port map( A1 => n225, A2 => n890, ZN => n127);
   U196 : OAI21_X1 port map( B1 => n128, B2 => n126, A => n127, ZN => 
                           intadd_0_A_12_port);
   U197 : OAI21_X1 port map( B1 => n128, B2 => C428_DATA4_15, A => n127, ZN => 
                           intadd_0_A_11_port);
   U198 : NAND2_X1 port map( A1 => n56, A2 => OP_A_14_port, ZN => n852);
   U199 : INV_X1 port map( A => n852, ZN => n129);
   U200 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_14, A => n129,
                           ZN => intadd_0_A_10_port);
   U201 : NAND2_X1 port map( A1 => n56, A2 => OP_A_13_port, ZN => n819);
   U202 : INV_X1 port map( A => n819, ZN => n130);
   U203 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_13, A => n130,
                           ZN => intadd_0_A_9_port);
   U204 : NAND2_X1 port map( A1 => n56, A2 => OP_A_12_port, ZN => n804);
   U205 : INV_X1 port map( A => n804, ZN => n131);
   U206 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_12, A => n131,
                           ZN => intadd_0_A_8_port);
   U207 : NAND2_X1 port map( A1 => n56, A2 => OP_A_11_port, ZN => n769);
   U208 : INV_X1 port map( A => n769, ZN => n132);
   U209 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_11, A => n132,
                           ZN => intadd_0_A_7_port);
   U210 : NAND2_X1 port map( A1 => n56, A2 => OP_A_10_port, ZN => n740);
   U211 : INV_X1 port map( A => n740, ZN => n133);
   U212 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_10, A => n133,
                           ZN => intadd_0_A_6_port);
   U213 : NAND2_X1 port map( A1 => n56, A2 => OP_A_9_port, ZN => n726);
   U214 : INV_X1 port map( A => n726, ZN => n134);
   U215 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_9, A => n134, 
                           ZN => intadd_0_A_5_port);
   U216 : NAND2_X1 port map( A1 => n56, A2 => OP_A_8_port, ZN => n696);
   U217 : INV_X1 port map( A => n696, ZN => n135);
   U218 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_8, A => n135, 
                           ZN => intadd_0_A_4_port);
   U219 : NAND2_X1 port map( A1 => n56, A2 => OP_A_7_port, ZN => n675);
   U220 : INV_X1 port map( A => n675, ZN => n136);
   U221 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_7, A => n136, 
                           ZN => intadd_0_A_3_port);
   U222 : NAND2_X1 port map( A1 => n56, A2 => OP_A_6_port, ZN => n658);
   U223 : INV_X1 port map( A => n658, ZN => n137);
   U224 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_6, A => n137, 
                           ZN => intadd_0_A_2_port);
   U225 : NAND2_X1 port map( A1 => n56, A2 => OP_A_5_port, ZN => n628);
   U226 : INV_X1 port map( A => n628, ZN => n138);
   U227 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_5, A => n138, 
                           ZN => intadd_0_A_1_port);
   U228 : INV_X1 port map( A => n894, ZN => n765);
   U229 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n581, ZN => n853);
   U230 : INV_X1 port map( A => n853, ZN => n742);
   U231 : AOI22_X1 port map( A1 => OP_B_1_port, A2 => n765, B1 => n742, B2 => 
                           n225, ZN => n150);
   U232 : AND2_X1 port map( A1 => n139, A2 => C2_DATA1_2, ZN => n140);
   U233 : AOI21_X1 port map( B1 => n62, B2 => OP_A_0_port, A => n140, ZN => 
                           n526);
   U234 : INV_X1 port map( A => OP_A_2_port, ZN => n576);
   U235 : NOR2_X1 port map( A1 => n510, A2 => n576, ZN => n552);
   U236 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_2, A => n552, 
                           ZN => n527);
   U237 : NOR2_X1 port map( A1 => n526, A2 => n527, ZN => n538);
   U238 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_3, B1 => 
                           OP_A_0_port, B2 => n149, C1 => n62, C2 => 
                           OP_A_1_port, ZN => n142);
   U239 : INV_X1 port map( A => n142, ZN => n535);
   U240 : INV_X1 port map( A => n538, ZN => n141);
   U241 : INV_X1 port map( A => OP_A_3_port, ZN => n550);
   U242 : NOR2_X1 port map( A1 => n510, A2 => n550, ZN => n580);
   U243 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_3, A => n580, 
                           ZN => n536);
   U244 : OAI21_X1 port map( B1 => n142, B2 => n141, A => n536, ZN => n143);
   U245 : OAI21_X1 port map( B1 => n538, B2 => n535, A => n143, ZN => 
                           intadd_0_A_0_port);
   U246 : XNOR2_X1 port map( A => DP_OP_456J3_131_2158_n17, B => n144, ZN => 
                           n146);
   U247 : OR2_X1 port map( A1 => n147, A2 => n1414, ZN => n145);
   U248 : OAI21_X1 port map( B1 => n147, B2 => n146, A => n145, ZN => 
                           intadd_0_B_14_port);
   U249 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_17, B1 => 
                           OP_A_15_port, B2 => n62, C1 => OP_A_14_port, C2 => 
                           n149, ZN => intadd_0_B_13_port);
   U250 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_16, B1 => 
                           OP_A_13_port, B2 => n149, C1 => OP_A_14_port, C2 => 
                           n62, ZN => intadd_0_B_12_port);
   U251 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_15, B1 => 
                           OP_A_12_port, B2 => n149, C1 => OP_A_13_port, C2 => 
                           n62, ZN => intadd_0_B_11_port);
   U252 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_14, B1 => 
                           OP_A_12_port, B2 => n62, C1 => OP_A_11_port, C2 => 
                           n149, ZN => intadd_0_B_10_port);
   U253 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_13, B1 => 
                           OP_A_11_port, B2 => n62, C1 => n149, C2 => 
                           OP_A_10_port, ZN => intadd_0_B_9_port);
   U254 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_12, B1 => n62, B2 
                           => OP_A_10_port, C1 => n149, C2 => OP_A_9_port, ZN 
                           => intadd_0_B_8_port);
   U255 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_11, B1 => n62, B2 
                           => OP_A_9_port, C1 => n149, C2 => OP_A_8_port, ZN =>
                           intadd_0_B_7_port);
   U256 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_10, B1 => n62, B2 
                           => OP_A_8_port, C1 => n149, C2 => OP_A_7_port, ZN =>
                           intadd_0_B_6_port);
   U257 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_9, B1 => n62, B2 =>
                           OP_A_7_port, C1 => n149, C2 => OP_A_6_port, ZN => 
                           intadd_0_B_5_port);
   U258 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_8, B1 => n62, B2 =>
                           OP_A_6_port, C1 => n149, C2 => OP_A_5_port, ZN => 
                           intadd_0_B_4_port);
   U259 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_7, B1 => n62, B2 =>
                           OP_A_5_port, C1 => n149, C2 => OP_A_4_port, ZN => 
                           intadd_0_B_3_port);
   U260 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_6, B1 => n62, B2 =>
                           OP_A_4_port, C1 => n149, C2 => OP_A_3_port, ZN => 
                           intadd_0_B_2_port);
   U261 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_5, B1 => n62, B2 =>
                           OP_A_3_port, C1 => n149, C2 => OP_A_2_port, ZN => 
                           intadd_0_B_1_port);
   U262 : NAND2_X1 port map( A1 => n56, A2 => OP_A_4_port, ZN => n604);
   U263 : INV_X1 port map( A => n604, ZN => n148);
   U264 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_4, A => n148, 
                           ZN => intadd_0_B_0_port);
   U265 : AOI222_X1 port map( A1 => n1414, A2 => C431_DATA4_4, B1 => n62, B2 =>
                           OP_A_2_port, C1 => n149, C2 => OP_A_1_port, ZN => 
                           intadd_0_CI);
   U266 : NOR2_X1 port map( A1 => OP_B_5_port, A2 => OP_B_6_port, ZN => n1081);
   U267 : NAND2_X1 port map( A1 => n1081, A2 => OP_B_7_port, ZN => n1078);
   U268 : INV_X1 port map( A => OP_B_6_port, ZN => n379);
   U269 : NOR2_X1 port map( A1 => n298, A2 => n379, ZN => n163);
   U270 : NOR3_X1 port map( A1 => n1081, A2 => n163, A3 => n296, ZN => n165);
   U271 : NAND2_X1 port map( A1 => n165, A2 => n1080, ZN => n1077);
   U272 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n1078, A => n1077, ZN =>
                           DP_OP_446J3_125_4819_n87);
   U273 : INV_X1 port map( A => n165, ZN => n151);
   U274 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n151, B1 => OP_A_13_port
                           , B2 => n1078, ZN => DP_OP_446J3_125_4819_n86);
   U275 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n151, B1 => OP_A_12_port
                           , B2 => n1078, ZN => DP_OP_446J3_125_4819_n85);
   U276 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n1078, B1 => 
                           OP_A_12_port, B2 => n151, ZN => 
                           DP_OP_446J3_125_4819_n84);
   U277 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n151, B1 => OP_A_10_port
                           , B2 => n1078, ZN => DP_OP_446J3_125_4819_n83);
   U278 : OAI22_X1 port map( A1 => OP_A_10_port, A2 => n151, B1 => OP_A_9_port,
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n82);
   U279 : OAI22_X1 port map( A1 => OP_A_9_port, A2 => n151, B1 => OP_A_8_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n81);
   U280 : OAI22_X1 port map( A1 => OP_A_8_port, A2 => n151, B1 => OP_A_7_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n80);
   U281 : OAI22_X1 port map( A1 => OP_A_7_port, A2 => n151, B1 => OP_A_6_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n79);
   U282 : OAI22_X1 port map( A1 => OP_A_6_port, A2 => n151, B1 => OP_A_5_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n78);
   U283 : OAI22_X1 port map( A1 => OP_A_5_port, A2 => n151, B1 => OP_A_4_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n77);
   U284 : OAI22_X1 port map( A1 => OP_A_4_port, A2 => n151, B1 => OP_A_3_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n76);
   U285 : OAI22_X1 port map( A1 => OP_A_3_port, A2 => n151, B1 => OP_A_2_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n75);
   U286 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n1078, B1 => OP_A_2_port,
                           B2 => n151, ZN => DP_OP_446J3_125_4819_n74);
   U287 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n151, B1 => OP_A_0_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n73);
   U288 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n151, A => n1078, ZN => 
                           DP_OP_446J3_125_4819_n72);
   U289 : AND2_X1 port map( A1 => C2_DATA1_4, A2 => n153, ZN => n154);
   U290 : AOI21_X1 port map( B1 => n161, B2 => OP_A_0_port, A => n154, ZN => 
                           n565);
   U291 : NOR2_X1 port map( A1 => intadd_0_SUM_0_port, A2 => n565, ZN => n564);
   U292 : INV_X1 port map( A => intadd_0_SUM_1_port, ZN => n158);
   U293 : INV_X1 port map( A => n564, ZN => n590);
   U294 : INV_X1 port map( A => n155, ZN => n156);
   U295 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_5, B1 => 
                           OP_A_0_port, B2 => n162, C1 => OP_A_1_port, C2 => 
                           n161, ZN => n591);
   U296 : OAI21_X1 port map( B1 => intadd_0_SUM_1_port, B2 => n590, A => n591, 
                           ZN => n157);
   U297 : OAI21_X1 port map( B1 => n564, B2 => n158, A => n157, ZN => 
                           intadd_1_A_0_port);
   U298 : XNOR2_X1 port map( A => DP_OP_451J3_128_3502_n15, B => n159, ZN => 
                           n160);
   U299 : OAI21_X1 port map( B1 => n1380, B2 => n160, A => n67, ZN => 
                           intadd_1_B_14_port);
   U300 : AOI222_X1 port map( A1 => OP_A_15_port, A2 => n161, B1 => n1412, B2 
                           => C430_DATA4_19, C1 => OP_A_14_port, C2 => n162, ZN
                           => intadd_1_B_13_port);
   U301 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_18, B1 => 
                           OP_A_13_port, B2 => n162, C1 => OP_A_14_port, C2 => 
                           n161, ZN => intadd_1_B_12_port);
   U302 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_17, B1 => 
                           OP_A_12_port, B2 => n162, C1 => OP_A_13_port, C2 => 
                           n161, ZN => intadd_1_B_11_port);
   U303 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_16, B1 => 
                           OP_A_12_port, B2 => n161, C1 => OP_A_11_port, C2 => 
                           n162, ZN => intadd_1_B_10_port);
   U304 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_14, B1 => n161, B2 
                           => OP_A_10_port, C1 => n162, C2 => OP_A_9_port, ZN 
                           => intadd_1_B_8_port);
   U305 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_13, B1 => n161, B2 
                           => OP_A_9_port, C1 => n162, C2 => OP_A_8_port, ZN =>
                           intadd_1_B_7_port);
   U306 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_12, B1 => n161, B2 
                           => OP_A_8_port, C1 => n162, C2 => OP_A_7_port, ZN =>
                           intadd_1_B_6_port);
   U307 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_11, B1 => n161, B2 
                           => OP_A_7_port, C1 => n162, C2 => OP_A_6_port, ZN =>
                           intadd_1_B_5_port);
   U308 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_10, B1 => n161, B2 
                           => OP_A_6_port, C1 => n162, C2 => OP_A_5_port, ZN =>
                           intadd_1_B_4_port);
   U309 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_9, B1 => n161, B2 
                           => OP_A_5_port, C1 => n162, C2 => OP_A_4_port, ZN =>
                           intadd_1_B_3_port);
   U310 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_8, B1 => n161, B2 
                           => OP_A_4_port, C1 => n162, C2 => OP_A_3_port, ZN =>
                           intadd_1_B_2_port);
   U311 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_7, B1 => n161, B2 
                           => OP_A_3_port, C1 => n162, C2 => OP_A_2_port, ZN =>
                           intadd_1_B_1_port);
   U312 : AOI222_X1 port map( A1 => n1412, A2 => C430_DATA4_6, B1 => 
                           OP_A_1_port, B2 => n162, C1 => n161, C2 => 
                           OP_A_2_port, ZN => intadd_1_B_0_port);
   U313 : CLKBUF_X1 port map( A => n1413, Z => n169);
   U314 : INV_X1 port map( A => n163, ZN => n164);
   U315 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_17, B1 => n63, B2 =>
                           OP_A_11_port, C1 => n1027, C2 => OP_A_10_port, ZN =>
                           intadd_2_A_9_port);
   U316 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_16, B1 => n63, B2 =>
                           OP_A_10_port, C1 => n1027, C2 => OP_A_9_port, ZN => 
                           intadd_2_A_8_port);
   U317 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_15, B1 => n63, B2 =>
                           OP_A_9_port, C1 => n1027, C2 => OP_A_8_port, ZN => 
                           intadd_2_A_7_port);
   U318 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_14, B1 => n63, B2 =>
                           OP_A_8_port, C1 => n1027, C2 => OP_A_7_port, ZN => 
                           intadd_2_A_6_port);
   U319 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_13, B1 => n63, B2 =>
                           OP_A_7_port, C1 => n1027, C2 => OP_A_6_port, ZN => 
                           intadd_2_A_5_port);
   U320 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_12, B1 => n63, B2 =>
                           OP_A_6_port, C1 => n1027, C2 => OP_A_5_port, ZN => 
                           intadd_2_A_4_port);
   U321 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_11, B1 => n63, B2 =>
                           OP_A_5_port, C1 => n1027, C2 => OP_A_4_port, ZN => 
                           intadd_2_A_3_port);
   U322 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_10, B1 => n63, B2 =>
                           OP_A_4_port, C1 => n1027, C2 => OP_A_3_port, ZN => 
                           intadd_2_A_2_port);
   U323 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_9, B1 => n63, B2 => 
                           OP_A_3_port, C1 => n1027, C2 => OP_A_2_port, ZN => 
                           intadd_2_A_1_port);
   U324 : AND2_X1 port map( A1 => C2_DATA1_6, A2 => n165, ZN => n166);
   U325 : AOI21_X1 port map( B1 => OP_A_0_port, B2 => n63, A => n166, ZN => 
                           n620);
   U326 : NOR2_X1 port map( A1 => intadd_1_SUM_0_port, A2 => n620, ZN => n619);
   U327 : INV_X1 port map( A => intadd_1_SUM_1_port, ZN => n168);
   U328 : INV_X1 port map( A => n619, ZN => n641);
   U329 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_7, B1 => n63, B2 => 
                           OP_A_1_port, C1 => n1027, C2 => OP_A_0_port, ZN => 
                           n642);
   U330 : OAI21_X1 port map( B1 => intadd_1_SUM_1_port, B2 => n641, A => n642, 
                           ZN => n167);
   U331 : OAI21_X1 port map( B1 => n619, B2 => n168, A => n167, ZN => 
                           intadd_2_A_0_port);
   U332 : AOI222_X1 port map( A1 => n169, A2 => C429_DATA4_8, B1 => n63, B2 => 
                           OP_A_2_port, C1 => n1027, C2 => OP_A_1_port, ZN => 
                           intadd_2_B_0_port);
   U333 : AOI21_X1 port map( B1 => n171, B2 => n173, A => n170, ZN => n172);
   U334 : OAI21_X1 port map( B1 => n176, B2 => n173, A => n172, ZN => N287);
   U335 : AOI21_X1 port map( B1 => n174, B2 => n1408, A => n181, ZN => n175);
   U336 : INV_X1 port map( A => n175, ZN => n177);
   U337 : OAI211_X1 port map( C1 => n178, C2 => n1407, A => n177, B => n176, ZN
                           => N288);
   U338 : INV_X1 port map( A => n179, ZN => n180);
   U339 : OAI21_X1 port map( B1 => n181, B2 => n1405, A => n180, ZN => N289);
   U340 : INV_X1 port map( A => OP2(0), ZN => n219);
   U341 : AOI22_X1 port map( A1 => OP2(0), A2 => n58, B1 => n198, B2 => n219, 
                           ZN => N247);
   U342 : INV_X1 port map( A => OP2(1), ZN => n485);
   U343 : AOI22_X1 port map( A1 => OP2(1), A2 => n58, B1 => n198, B2 => n485, 
                           ZN => N248);
   U344 : INV_X1 port map( A => OP2(2), ZN => n182);
   U345 : AOI22_X1 port map( A1 => OP2(2), A2 => n58, B1 => n198, B2 => n182, 
                           ZN => N249);
   U346 : INV_X1 port map( A => OP2(3), ZN => n183);
   U347 : AOI22_X1 port map( A1 => OP2(3), A2 => n58, B1 => n198, B2 => n183, 
                           ZN => N250);
   U348 : INV_X1 port map( A => OP2(4), ZN => n184);
   U349 : AOI22_X1 port map( A1 => OP2(4), A2 => n58, B1 => n198, B2 => n184, 
                           ZN => N251);
   U350 : INV_X1 port map( A => OP2(5), ZN => n612);
   U351 : AOI22_X1 port map( A1 => OP2(5), A2 => n58, B1 => n198, B2 => n612, 
                           ZN => N252);
   U352 : INV_X1 port map( A => OP2(6), ZN => n185);
   U353 : AOI22_X1 port map( A1 => OP2(6), A2 => n58, B1 => n198, B2 => n185, 
                           ZN => N253);
   U354 : INV_X1 port map( A => OP2(7), ZN => n664);
   U355 : AOI22_X1 port map( A1 => OP2(7), A2 => n58, B1 => n198, B2 => n664, 
                           ZN => N254);
   U356 : INV_X1 port map( A => OP2(8), ZN => n186);
   U357 : AOI22_X1 port map( A1 => OP2(8), A2 => n58, B1 => n198, B2 => n186, 
                           ZN => N255);
   U358 : INV_X1 port map( A => OP2(9), ZN => n691);
   U359 : AOI22_X1 port map( A1 => OP2(9), A2 => n58, B1 => n198, B2 => n691, 
                           ZN => N256);
   U360 : INV_X1 port map( A => OP2(10), ZN => n187);
   U361 : AOI22_X1 port map( A1 => OP2(10), A2 => n58, B1 => n198, B2 => n187, 
                           ZN => N257);
   U362 : INV_X1 port map( A => OP2(11), ZN => n188);
   U363 : AOI22_X1 port map( A1 => OP2(11), A2 => n58, B1 => n198, B2 => n188, 
                           ZN => N258);
   U364 : INV_X1 port map( A => OP2(12), ZN => n776);
   U365 : AOI22_X1 port map( A1 => OP2(12), A2 => n58, B1 => n198, B2 => n776, 
                           ZN => N259);
   U366 : INV_X1 port map( A => OP2(13), ZN => n800);
   U367 : AOI22_X1 port map( A1 => OP2(13), A2 => n58, B1 => n198, B2 => n800, 
                           ZN => N260);
   U368 : INV_X1 port map( A => OP2(14), ZN => n189);
   U369 : AOI22_X1 port map( A1 => OP2(14), A2 => n58, B1 => n198, B2 => n189, 
                           ZN => N261);
   U370 : INV_X1 port map( A => OP2(15), ZN => n859);
   U371 : AOI22_X1 port map( A1 => OP2(15), A2 => n58, B1 => n198, B2 => n859, 
                           ZN => N262);
   U372 : INV_X1 port map( A => OP2(16), ZN => n190);
   U373 : AOI22_X1 port map( A1 => OP2(16), A2 => n58, B1 => n198, B2 => n190, 
                           ZN => N263);
   U374 : INV_X1 port map( A => OP2(17), ZN => n191);
   U375 : AOI22_X1 port map( A1 => OP2(17), A2 => n196, B1 => n198, B2 => n191,
                           ZN => N264);
   U376 : INV_X1 port map( A => OP2(18), ZN => n192);
   U377 : AOI22_X1 port map( A1 => OP2(18), A2 => n196, B1 => n198, B2 => n192,
                           ZN => N265);
   U378 : INV_X1 port map( A => OP2(19), ZN => n193);
   U379 : AOI22_X1 port map( A1 => OP2(19), A2 => n196, B1 => n198, B2 => n193,
                           ZN => N266);
   U380 : INV_X1 port map( A => OP2(20), ZN => n194);
   U381 : AOI22_X1 port map( A1 => OP2(20), A2 => n196, B1 => n198, B2 => n194,
                           ZN => N267);
   U382 : INV_X1 port map( A => OP2(21), ZN => n195);
   U383 : AOI22_X1 port map( A1 => OP2(21), A2 => n196, B1 => n198, B2 => n195,
                           ZN => N268);
   U384 : INV_X1 port map( A => OP2(22), ZN => n197);
   U385 : AOI22_X1 port map( A1 => OP2(22), A2 => n58, B1 => n198, B2 => n197, 
                           ZN => N269);
   U386 : INV_X1 port map( A => OP2(23), ZN => n199);
   U387 : AOI22_X1 port map( A1 => OP2(23), A2 => n58, B1 => n198, B2 => n199, 
                           ZN => N270);
   U388 : INV_X1 port map( A => OP2(24), ZN => n1137);
   U389 : AOI22_X1 port map( A1 => OP2(24), A2 => n58, B1 => n198, B2 => n1137,
                           ZN => N271);
   U390 : INV_X1 port map( A => OP2(25), ZN => n200);
   U391 : AOI22_X1 port map( A1 => OP2(25), A2 => n58, B1 => n198, B2 => n200, 
                           ZN => N272);
   U392 : INV_X1 port map( A => OP2(26), ZN => n201);
   U393 : AOI22_X1 port map( A1 => OP2(26), A2 => n58, B1 => n198, B2 => n201, 
                           ZN => N273);
   U394 : INV_X1 port map( A => OP2(27), ZN => n202);
   U395 : AOI22_X1 port map( A1 => OP2(27), A2 => n58, B1 => n198, B2 => n202, 
                           ZN => N274);
   U396 : INV_X1 port map( A => OP2(28), ZN => n203);
   U397 : AOI22_X1 port map( A1 => OP2(28), A2 => n58, B1 => n198, B2 => n203, 
                           ZN => N275);
   U398 : INV_X1 port map( A => OP2(29), ZN => n204);
   U399 : AOI22_X1 port map( A1 => OP2(29), A2 => n58, B1 => n198, B2 => n204, 
                           ZN => N276);
   U400 : INV_X1 port map( A => OP2(30), ZN => n205);
   U401 : AOI22_X1 port map( A1 => OP2(30), A2 => n58, B1 => n198, B2 => n205, 
                           ZN => N277);
   U402 : INV_X1 port map( A => OP2(31), ZN => n206);
   U403 : AOI22_X1 port map( A1 => OP2(31), A2 => n58, B1 => n198, B2 => n206, 
                           ZN => N278);
   U404 : INV_X1 port map( A => N284, ZN => n1158);
   U405 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => n55, ZN => n1203);
   U406 : NAND2_X1 port map( A1 => n56, A2 => OP_A_21_port, ZN => n1058);
   U407 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => n603, ZN => n1132);
   U408 : OR2_X1 port map( A1 => OP_B_1_port, A2 => OP_B_0_port, ZN => n607);
   U409 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => n57, ZN => n1002);
   U410 : AND4_X1 port map( A1 => n1203, A2 => n1058, A3 => n1132, A4 => n1002,
                           ZN => n784);
   U411 : NAND2_X1 port map( A1 => n56, A2 => OP_A_25_port, ZN => n1204);
   U412 : NAND2_X1 port map( A1 => OP_A_27_port, A2 => n55, ZN => n1317);
   U413 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => n57, ZN => n1129);
   U414 : CLKBUF_X1 port map( A => n603, Z => n553);
   U415 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => n553, ZN => n1271);
   U416 : NAND4_X1 port map( A1 => n1204, A2 => n1317, A3 => n1129, A4 => n1271
                           , ZN => n781);
   U417 : INV_X1 port map( A => n857, ZN => n511);
   U418 : INV_X1 port map( A => OP_A_31_port, ZN => n1369);
   U419 : AOI22_X1 port map( A1 => OP_A_30_port, A2 => n603, B1 => OP_A_28_port
                           , B2 => n57, ZN => n207);
   U420 : NAND2_X1 port map( A1 => n56, A2 => OP_A_29_port, ZN => n1318);
   U421 : OAI211_X1 port map( C1 => n577, C2 => n1369, A => n207, B => n1318, 
                           ZN => n1264);
   U422 : AOI22_X1 port map( A1 => n855, A2 => n781, B1 => n511, B2 => n1264, 
                           ZN => n209);
   U423 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => n55, ZN => n1057);
   U424 : NAND2_X1 port map( A1 => n56, A2 => OP_A_17_port, ZN => n937);
   U425 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => n553, ZN => n1005);
   U426 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n57, ZN => n887);
   U427 : NAND4_X1 port map( A1 => n1057, A2 => n937, A3 => n1005, A4 => n887, 
                           ZN => n777);
   U428 : NAND2_X1 port map( A1 => n894, A2 => n777, ZN => n208);
   U429 : OAI211_X1 port map( C1 => n784, C2 => n742, A => n209, B => n208, ZN 
                           => n898);
   U430 : NAND2_X1 port map( A1 => OP_A_15_port, A2 => n55, ZN => n936);
   U431 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => n57, ZN => n767);
   U432 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => n553, ZN => n889);
   U433 : AND4_X1 port map( A1 => n819, A2 => n936, A3 => n767, A4 => n889, ZN 
                           => n771);
   U434 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n857, ZN => n1351);
   U435 : INV_X1 port map( A => n1351, ZN => n891);
   U436 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => n55, ZN => n817);
   U437 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => n553, ZN => n768);
   U438 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => n57, ZN => n672);
   U439 : AND4_X1 port map( A1 => n817, A2 => n726, A3 => n768, A4 => n672, ZN 
                           => n681);
   U440 : INV_X1 port map( A => n855, ZN => n741);
   U441 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n741, ZN => n1349);
   U442 : INV_X1 port map( A => n1349, ZN => n566);
   U443 : OAI22_X1 port map( A1 => n771, A2 => n891, B1 => n681, B2 => n566, ZN
                           => n215);
   U444 : NAND2_X1 port map( A1 => OP_A_3_port, A2 => n55, ZN => n626);
   U445 : NAND2_X1 port map( A1 => n56, A2 => OP_A_1_port, ZN => n508);
   U446 : NAND2_X1 port map( A1 => OP_A_0_port, A2 => n57, ZN => n895);
   U447 : NAND2_X1 port map( A1 => OP_A_2_port, A2 => n553, ZN => n210);
   U448 : AND4_X1 port map( A1 => n626, A2 => n508, A3 => n895, A4 => n210, ZN 
                           => n213);
   U449 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n765, ZN => n1359);
   U450 : INV_X1 port map( A => n1359, ZN => n1260);
   U451 : NAND2_X1 port map( A1 => OP_A_7_port, A2 => n55, ZN => n725);
   U452 : NAND2_X1 port map( A1 => OP_A_4_port, A2 => n57, ZN => n211);
   U453 : NAND2_X1 port map( A1 => OP_A_6_port, A2 => n553, ZN => n674);
   U454 : NAND4_X1 port map( A1 => n725, A2 => n628, A3 => n211, A4 => n674, ZN
                           => n582);
   U455 : INV_X1 port map( A => n582, ZN => n212);
   U456 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n742, ZN => n1357);
   U457 : INV_X1 port map( A => n1357, ZN => n899);
   U458 : OAI22_X1 port map( A1 => n213, A2 => n1260, B1 => n212, B2 => n899, 
                           ZN => n214);
   U459 : AOI211_X1 port map( C1 => OP_B_4_port, C2 => n898, A => n215, B => 
                           n214, ZN => n483);
   U460 : NOR2_X1 port map( A1 => n217, A2 => n216, ZN => n1346);
   U461 : CLKBUF_X1 port map( A => n1346, Z => n1329);
   U462 : NAND2_X1 port map( A1 => OP_B_0_port, A2 => OP_A_0_port, ZN => n294);
   U463 : OR2_X1 port map( A1 => n218, A2 => n1410, ZN => n1138);
   U464 : OAI22_X1 port map( A1 => n1395, A2 => n294, B1 => n1138, B2 => n219, 
                           ZN => n222);
   U465 : NOR2_X1 port map( A1 => n220, A2 => OP_LOGIC_0_port, ZN => n476);
   U466 : INV_X1 port map( A => OP_LOGIC_1_port, ZN => n223);
   U467 : AND2_X1 port map( A1 => n476, A2 => n223, ZN => n1244);
   U468 : INV_X1 port map( A => n1244, ZN => n1368);
   U469 : INV_X1 port map( A => n1227, ZN => n1061);
   U470 : OAI22_X1 port map( A1 => n294, A2 => n1368, B1 => n895, B2 => n1061, 
                           ZN => n221);
   U471 : AOI211_X1 port map( C1 => n1329, C2 => OP1(0), A => n222, B => n221, 
                           ZN => n482);
   U472 : NAND3_X1 port map( A1 => N281, A2 => n223, A3 => OP_LOGIC_0_port, ZN 
                           => n1367);
   U473 : INV_X1 port map( A => OP_A_0_port, ZN => n549);
   U474 : NAND2_X1 port map( A1 => n224, A2 => n549, ZN => n489);
   U475 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n550, ZN => n366);
   U476 : INV_X1 port map( A => n366, ZN => n317);
   U477 : INV_X1 port map( A => OP_A_5_port, ZN => n606);
   U478 : NAND2_X1 port map( A1 => n606, A2 => OP_B_5_port, ZN => n370);
   U479 : OAI21_X1 port map( B1 => n1362, B2 => OP_A_4_port, A => n370, ZN => 
                           n321);
   U480 : INV_X1 port map( A => OP_A_1_port, ZN => n578);
   U481 : OAI21_X1 port map( B1 => n225, B2 => OP_A_1_port, A => OP_A_0_port, 
                           ZN => n316);
   U482 : OAI211_X1 port map( C1 => n578, C2 => n55, A => n607, B => n316, ZN 
                           => n367);
   U483 : NOR2_X1 port map( A1 => OP_A_3_port, A2 => n1159, ZN => n303);
   U484 : AOI21_X1 port map( B1 => n576, B2 => OP_B_2_port, A => n303, ZN => 
                           n365);
   U485 : INV_X1 port map( A => n303, ZN => n318);
   U486 : NOR2_X1 port map( A1 => n576, A2 => OP_B_2_port, ZN => n226);
   U487 : AOI22_X1 port map( A1 => n367, A2 => n365, B1 => n318, B2 => n226, ZN
                           => n228);
   U488 : INV_X1 port map( A => OP_A_4_port, ZN => n369);
   U489 : NOR2_X1 port map( A1 => n369, A2 => OP_B_4_port, ZN => n227);
   U490 : NOR2_X1 port map( A1 => n606, A2 => OP_B_5_port, ZN => n372);
   U491 : AOI21_X1 port map( B1 => n370, B2 => n227, A => n372, ZN => n320);
   U492 : OAI221_X1 port map( B1 => n317, B2 => n321, C1 => n228, C2 => n321, A
                           => n320, ZN => n234);
   U493 : NAND2_X1 port map( A1 => n379, A2 => OP_A_6_port, ZN => n229);
   U494 : NOR2_X1 port map( A1 => n296, A2 => OP_A_7_port, ZN => n380);
   U495 : NAND2_X1 port map( A1 => n296, A2 => OP_A_7_port, ZN => n381);
   U496 : OAI21_X1 port map( B1 => n229, B2 => n380, A => n381, ZN => n323);
   U497 : INV_X1 port map( A => OP_A_6_port, ZN => n373);
   U498 : AOI21_X1 port map( B1 => n373, B2 => OP_B_6_port, A => n380, ZN => 
                           n325);
   U499 : INV_X1 port map( A => OP_A_12_port, ZN => n235);
   U500 : NAND2_X1 port map( A1 => n235, A2 => OP_B_12_port, ZN => n334);
   U501 : INV_X1 port map( A => OP_A_13_port, ZN => n236);
   U502 : INV_X1 port map( A => OP_B_14_port, ZN => n230);
   U503 : NAND2_X1 port map( A1 => n1080, A2 => OP_B_15_port, ZN => n350);
   U504 : OAI21_X1 port map( B1 => n230, B2 => OP_A_14_port, A => n350, ZN => 
                           n231);
   U505 : AOI21_X1 port map( B1 => n236, B2 => OP_B_13_port, A => n231, ZN => 
                           n242);
   U506 : AND2_X1 port map( A1 => n334, A2 => n242, ZN => n232);
   U507 : INV_X1 port map( A => OP_A_10_port, ZN => n337);
   U508 : INV_X1 port map( A => OP_A_11_port, ZN => n237);
   U509 : NAND2_X1 port map( A1 => n237, A2 => OP_B_11_port, ZN => n344);
   U510 : INV_X1 port map( A => n344, ZN => n241);
   U511 : AOI21_X1 port map( B1 => OP_B_10_port, B2 => n337, A => n241, ZN => 
                           n239);
   U512 : INV_X1 port map( A => OP_A_9_port, ZN => n304);
   U513 : INV_X1 port map( A => OP_A_8_port, ZN => n238);
   U514 : AOI22_X1 port map( A1 => OP_B_9_port, A2 => n304, B1 => OP_B_8_port, 
                           B2 => n238, ZN => n340);
   U515 : NAND3_X1 port map( A1 => n232, A2 => n239, A3 => n340, ZN => n327);
   U516 : INV_X1 port map( A => n327, ZN => n233);
   U517 : OAI221_X1 port map( B1 => n234, B2 => n323, C1 => n325, C2 => n323, A
                           => n233, ZN => n250_port);
   U518 : INV_X1 port map( A => OP_A_14_port, ZN => n333);
   U519 : NOR2_X1 port map( A1 => n333, A2 => OP_B_14_port, ZN => n347);
   U520 : OAI22_X1 port map( A1 => OP_B_13_port, A2 => n236, B1 => OP_B_12_port
                           , B2 => n235, ZN => n336);
   U521 : OR2_X1 port map( A1 => n337, A2 => OP_B_10_port, ZN => n338);
   U522 : NOR2_X1 port map( A1 => n237, A2 => OP_B_11_port, ZN => n346);
   U523 : INV_X1 port map( A => n346, ZN => n339);
   U524 : INV_X1 port map( A => OP_B_9_port, ZN => n341);
   U525 : OAI22_X1 port map( A1 => OP_B_8_port, A2 => n238, B1 => OP_B_9_port, 
                           B2 => n304, ZN => n358);
   U526 : OAI211_X1 port map( C1 => OP_A_9_port, C2 => n341, A => n239, B => 
                           n358, ZN => n240);
   U527 : OAI211_X1 port map( C1 => n241, C2 => n338, A => n339, B => n240, ZN 
                           => n243);
   U528 : OAI221_X1 port map( B1 => n336, B2 => n334, C1 => n336, C2 => n243, A
                           => n242, ZN => n244);
   U529 : INV_X1 port map( A => n244, ZN => n245);
   U530 : NOR2_X1 port map( A1 => n1080, A2 => OP_B_15_port, ZN => n353);
   U531 : AOI211_X1 port map( C1 => n350, C2 => n347, A => n245, B => n353, ZN 
                           => n328);
   U532 : INV_X1 port map( A => OP_B_17_port, ZN => n257_port);
   U533 : NOR2_X1 port map( A1 => OP_A_17_port, A2 => n257_port, ZN => n395);
   U534 : INV_X1 port map( A => OP_B_16_port, ZN => n258_port);
   U535 : NOR2_X1 port map( A1 => OP_A_16_port, A2 => n258_port, ZN => n396);
   U536 : INV_X1 port map( A => OP_B_18_port, ZN => n359);
   U537 : INV_X1 port map( A => OP_A_19_port, ZN => n256_port);
   U538 : NAND2_X1 port map( A1 => OP_B_19_port, A2 => n256_port, ZN => n398);
   U539 : OAI21_X1 port map( B1 => OP_A_18_port, B2 => n359, A => n398, ZN => 
                           n259_port);
   U540 : INV_X1 port map( A => OP_A_21_port, ZN => n247_port);
   U541 : INV_X1 port map( A => OP_B_22_port, ZN => n391);
   U542 : INV_X1 port map( A => OP_A_23_port, ZN => n254_port);
   U543 : NAND2_X1 port map( A1 => OP_B_23_port, A2 => n254_port, ZN => n409);
   U544 : OAI21_X1 port map( B1 => OP_A_22_port, B2 => n391, A => n409, ZN => 
                           n246_port);
   U545 : AOI21_X1 port map( B1 => OP_B_21_port, B2 => n247_port, A => 
                           n246_port, ZN => n248_port);
   U546 : INV_X1 port map( A => n248_port, ZN => n262_port);
   U547 : INV_X1 port map( A => OP_B_20_port, ZN => n255_port);
   U548 : NOR2_X1 port map( A1 => n255_port, A2 => OP_A_20_port, ZN => n401);
   U549 : OR2_X1 port map( A1 => n262_port, A2 => n401, ZN => n249_port);
   U550 : OR4_X1 port map( A1 => n395, A2 => n396, A3 => n259_port, A4 => 
                           n249_port, ZN => n326);
   U551 : AOI21_X1 port map( B1 => n250_port, B2 => n328, A => n326, ZN => 
                           n251_port);
   U552 : INV_X1 port map( A => n251_port, ZN => n286_port);
   U553 : INV_X1 port map( A => OP_B_24_port, ZN => n418);
   U554 : INV_X1 port map( A => OP_A_25_port, ZN => n267_port);
   U555 : NAND2_X1 port map( A1 => n267_port, A2 => OP_B_25_port, ZN => n419);
   U556 : INV_X1 port map( A => OP_A_26_port, ZN => n424);
   U557 : INV_X1 port map( A => OP_A_27_port, ZN => n1247);
   U558 : NAND2_X1 port map( A1 => OP_B_27_port, A2 => n1247, ZN => n426);
   U559 : INV_X1 port map( A => n426, ZN => n272_port);
   U560 : AOI21_X1 port map( B1 => n424, B2 => OP_B_26_port, A => n272_port, ZN
                           => n268_port);
   U561 : OAI211_X1 port map( C1 => n418, C2 => OP_A_24_port, A => n419, B => 
                           n268_port, ZN => n278_port);
   U562 : INV_X1 port map( A => OP_B_28_port, ZN => n276_port);
   U563 : INV_X1 port map( A => OP_A_29_port, ZN => n1296);
   U564 : NAND2_X1 port map( A1 => n1296, A2 => OP_B_29_port, ZN => n414);
   U565 : NOR2_X1 port map( A1 => OP_B_31_port, A2 => n1369, ZN => n429);
   U566 : INV_X1 port map( A => OP_A_30_port, ZN => n253_port);
   U567 : NAND2_X1 port map( A1 => OP_B_30_port, A2 => n253_port, ZN => n453);
   U568 : INV_X1 port map( A => n453, ZN => n412);
   U569 : NOR2_X1 port map( A1 => n429, A2 => n412, ZN => n273_port);
   U570 : OAI211_X1 port map( C1 => n276_port, C2 => OP_A_28_port, A => n414, B
                           => n273_port, ZN => n252_port);
   U571 : OR2_X1 port map( A1 => n278_port, A2 => n252_port, ZN => n464);
   U572 : NOR2_X1 port map( A1 => OP_B_30_port, A2 => n253_port, ZN => n441);
   U573 : INV_X1 port map( A => n429, ZN => n451);
   U574 : NAND2_X1 port map( A1 => n1369, A2 => OP_B_31_port, ZN => n307);
   U575 : INV_X1 port map( A => n307, ZN => n454);
   U576 : AND2_X1 port map( A1 => n391, A2 => OP_A_22_port, ZN => n265_port);
   U577 : NOR2_X1 port map( A1 => OP_B_23_port, A2 => n254_port, ZN => n410);
   U578 : INV_X1 port map( A => OP_B_21_port, ZN => n403);
   U579 : AOI22_X1 port map( A1 => OP_A_21_port, A2 => n403, B1 => OP_A_20_port
                           , B2 => n255_port, ZN => n405);
   U580 : INV_X1 port map( A => OP_A_18_port, ZN => n392);
   U581 : NOR2_X1 port map( A1 => OP_B_18_port, A2 => n392, ZN => n261_port);
   U582 : NOR2_X1 port map( A1 => OP_B_19_port, A2 => n256_port, ZN => n399);
   U583 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n257_port, ZN => n394);
   U584 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n258_port, ZN => n361);
   U585 : AOI211_X1 port map( C1 => n394, C2 => n361, A => n395, B => n259_port
                           , ZN => n260_port);
   U586 : AOI211_X1 port map( C1 => n261_port, C2 => n398, A => n399, B => 
                           n260_port, ZN => n263_port);
   U587 : AOI221_X1 port map( B1 => n401, B2 => n405, C1 => n263_port, C2 => 
                           n405, A => n262_port, ZN => n264_port);
   U588 : AOI211_X1 port map( C1 => n265_port, C2 => n409, A => n410, B => 
                           n264_port, ZN => n284_port);
   U589 : INV_X1 port map( A => n414, ZN => n290);
   U590 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n276_port, ZN => 
                           n266_port);
   U591 : NOR2_X1 port map( A1 => OP_B_29_port, A2 => n1296, ZN => n416);
   U592 : INV_X1 port map( A => n416, ZN => n363);
   U593 : OAI21_X1 port map( B1 => n290, B2 => n266_port, A => n363, ZN => 
                           n282_port);
   U594 : INV_X1 port map( A => OP_A_28_port, ZN => n413);
   U595 : AOI21_X1 port map( B1 => OP_B_28_port, B2 => n413, A => n290, ZN => 
                           n281_port);
   U596 : OR2_X1 port map( A1 => n424, A2 => OP_B_26_port, ZN => n271_port);
   U597 : NOR2_X1 port map( A1 => OP_B_25_port, A2 => n267_port, ZN => n420);
   U598 : AND2_X1 port map( A1 => n418, A2 => OP_A_24_port, ZN => n269_port);
   U599 : OAI211_X1 port map( C1 => n420, C2 => n269_port, A => n419, B => 
                           n268_port, ZN => n270_port);
   U600 : OR2_X1 port map( A1 => n1247, A2 => OP_B_27_port, ZN => n423);
   U601 : OAI211_X1 port map( C1 => n272_port, C2 => n271_port, A => n270_port,
                           B => n423, ZN => n280_port);
   U602 : OAI221_X1 port map( B1 => n282_port, B2 => n281_port, C1 => n282_port
                           , C2 => n280_port, A => n273_port, ZN => n274_port);
   U603 : OAI21_X1 port map( B1 => n284_port, B2 => n464, A => n274_port, ZN =>
                           n275_port);
   U604 : AOI211_X1 port map( C1 => n441, C2 => n451, A => n454, B => n275_port
                           , ZN => n462);
   U605 : OAI21_X1 port map( B1 => n286_port, B2 => n464, A => n462, ZN => 
                           n288_port);
   U606 : NOR2_X1 port map( A1 => OP_COMPARE_1_port, A2 => OP_COMPARE_2_port, 
                           ZN => n439);
   U607 : NOR2_X1 port map( A1 => n454, A2 => n412, ZN => n279_port);
   U608 : OAI211_X1 port map( C1 => n276_port, C2 => OP_A_28_port, A => n414, B
                           => n279_port, ZN => n277_port);
   U609 : OR2_X1 port map( A1 => n278_port, A2 => n277_port, ZN => n331);
   U610 : OAI221_X1 port map( B1 => n282_port, B2 => n281_port, C1 => n282_port
                           , C2 => n280_port, A => n279_port, ZN => n283_port);
   U611 : OAI21_X1 port map( B1 => n284_port, B2 => n331, A => n283_port, ZN =>
                           n285_port);
   U612 : AOI211_X1 port map( C1 => n441, C2 => n307, A => n429, B => n285_port
                           , ZN => n330);
   U613 : OAI211_X1 port map( C1 => n331, C2 => n286_port, A => 
                           OP_COMPARE_0_port, B => n330, ZN => n287_port);
   U614 : OAI211_X1 port map( C1 => OP_COMPARE_0_port, C2 => n288_port, A => 
                           n439, B => n287_port, ZN => n475);
   U615 : INV_X1 port map( A => OP_COMPARE_3_port, ZN => n474);
   U616 : NAND2_X1 port map( A1 => n426, A2 => n423, ZN => n1240);
   U617 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => OP_B_19_port, ZN => n975
                           );
   U618 : OR2_X1 port map( A1 => OP_A_19_port, A2 => OP_B_19_port, ZN => n991);
   U619 : NAND2_X1 port map( A1 => n975, A2 => n991, ZN => n974);
   U620 : INV_X1 port map( A => n974, ZN => n983);
   U621 : NOR2_X1 port map( A1 => OP_A_23_port, A2 => OP_B_23_port, ZN => n1107
                           );
   U622 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => OP_B_23_port, ZN => 
                           n1122);
   U623 : INV_X1 port map( A => n1122, ZN => n289_port);
   U624 : NOR2_X1 port map( A1 => n1107, A2 => n289_port, ZN => n1105);
   U625 : AND2_X1 port map( A1 => OP_A_15_port, A2 => OP_B_15_port, ZN => n877)
                           ;
   U626 : NOR2_X1 port map( A1 => OP_A_15_port, A2 => OP_B_15_port, ZN => n862)
                           ;
   U627 : NOR2_X1 port map( A1 => n877, A2 => n862, ZN => n873);
   U628 : OR4_X1 port map( A1 => n1240, A2 => n983, A3 => n1105, A4 => n873, ZN
                           => n302);
   U629 : NOR2_X1 port map( A1 => n290, A2 => n416, ZN => n1301);
   U630 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => OP_B_26_port, ZN => 
                           n1236);
   U631 : OAI21_X1 port map( B1 => OP_A_26_port, B2 => OP_B_26_port, A => n1236
                           , ZN => n1199);
   U632 : NOR2_X1 port map( A1 => OP_A_30_port, A2 => OP_B_30_port, ZN => n1374
                           );
   U633 : NAND2_X1 port map( A1 => OP_A_30_port, A2 => OP_B_30_port, ZN => 
                           n1376);
   U634 : INV_X1 port map( A => n1376, ZN => n291);
   U635 : NOR2_X1 port map( A1 => n1374, A2 => n291, ZN => n1342);
   U636 : INV_X1 port map( A => n1342, ZN => n1332);
   U637 : NOR2_X1 port map( A1 => OP_A_28_port, A2 => OP_B_28_port, ZN => n1298
                           );
   U638 : INV_X1 port map( A => n1298, ZN => n292);
   U639 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => OP_B_28_port, ZN => 
                           n1300);
   U640 : NAND2_X1 port map( A1 => n292, A2 => n1300, ZN => n1266);
   U641 : NAND4_X1 port map( A1 => n1301, A2 => n1199, A3 => n1332, A4 => n1266
                           , ZN => n301);
   U642 : NAND2_X1 port map( A1 => n1362, A2 => n369, ZN => n597);
   U643 : NAND2_X1 port map( A1 => OP_B_4_port, A2 => OP_A_4_port, ZN => n570);
   U644 : NAND2_X1 port map( A1 => n597, A2 => n570, ZN => n573);
   U645 : NAND2_X1 port map( A1 => n581, A2 => n576, ZN => n546);
   U646 : NOR2_X1 port map( A1 => n581, A2 => n576, ZN => n507);
   U647 : INV_X1 port map( A => n507, ZN => n293);
   U648 : NAND2_X1 port map( A1 => n546, A2 => n293, ZN => n524);
   U649 : NOR2_X1 port map( A1 => OP_B_1_port, A2 => OP_A_1_port, ZN => n521);
   U650 : INV_X1 port map( A => n521, ZN => n503);
   U651 : NAND2_X1 port map( A1 => OP_B_1_port, A2 => OP_A_1_port, ZN => n520);
   U652 : NAND2_X1 port map( A1 => n503, A2 => n520, ZN => n506);
   U653 : NAND2_X1 port map( A1 => n294, A2 => n489, ZN => n477);
   U654 : NAND4_X1 port map( A1 => n573, A2 => n524, A3 => n506, A4 => n477, ZN
                           => n300);
   U655 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => OP_B_11_port, ZN => n749
                           );
   U656 : OR2_X1 port map( A1 => OP_A_11_port, A2 => OP_B_11_port, ZN => n773);
   U657 : NAND2_X1 port map( A1 => n749, A2 => n773, ZN => n754);
   U658 : NAND2_X1 port map( A1 => OP_B_7_port, A2 => OP_A_7_port, ZN => n645);
   U659 : INV_X1 port map( A => OP_A_7_port, ZN => n295);
   U660 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => n678);
   U661 : NAND2_X1 port map( A1 => n645, A2 => n678, ZN => n653);
   U662 : NAND2_X1 port map( A1 => OP_B_6_port, A2 => OP_A_6_port, ZN => n649);
   U663 : NOR2_X1 port map( A1 => OP_B_6_port, A2 => OP_A_6_port, ZN => n651);
   U664 : INV_X1 port map( A => n651, ZN => n297);
   U665 : NAND2_X1 port map( A1 => n649, A2 => n297, ZN => n636);
   U666 : NAND2_X1 port map( A1 => OP_B_5_port, A2 => OP_A_5_port, ZN => n593);
   U667 : NAND2_X1 port map( A1 => n298, A2 => n606, ZN => n632);
   U668 : NAND2_X1 port map( A1 => n593, A2 => n632, ZN => n600);
   U669 : NAND4_X1 port map( A1 => n754, A2 => n653, A3 => n636, A4 => n600, ZN
                           => n299);
   U670 : NOR4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN 
                           => n315);
   U671 : NOR2_X1 port map( A1 => n366, A2 => n303, ZN => n557);
   U672 : NOR2_X1 port map( A1 => OP_A_13_port, A2 => OP_B_13_port, ZN => n831)
                           ;
   U673 : INV_X1 port map( A => n831, ZN => n793);
   U674 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => OP_B_13_port, ZN => n829
                           );
   U675 : NAND2_X1 port map( A1 => n793, A2 => n829, ZN => n798);
   U676 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => OP_B_8_port, ZN => n711);
   U677 : NOR2_X1 port map( A1 => OP_A_8_port, A2 => OP_B_8_port, ZN => n715);
   U678 : INV_X1 port map( A => n715, ZN => n671);
   U679 : NAND2_X1 port map( A1 => n711, A2 => n671, ZN => n680);
   U680 : NOR2_X1 port map( A1 => OP_A_9_port, A2 => OP_B_9_port, ZN => n714);
   U681 : NOR2_X1 port map( A1 => n304, A2 => n341, ZN => n698);
   U682 : NOR2_X1 port map( A1 => n714, A2 => n698, ZN => n702);
   U683 : INV_X1 port map( A => n702, ZN => n305);
   U684 : NAND4_X1 port map( A1 => n557, A2 => n798, A3 => n680, A4 => n305, ZN
                           => n313);
   U685 : NOR2_X1 port map( A1 => OP_A_21_port, A2 => OP_B_21_port, ZN => n1050
                           );
   U686 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => OP_B_21_port, ZN => 
                           n1048);
   U687 : INV_X1 port map( A => n1048, ZN => n1021);
   U688 : NOR2_X1 port map( A1 => n1050, A2 => n1021, ZN => n1020);
   U689 : NOR2_X1 port map( A1 => OP_A_25_port, A2 => OP_B_25_port, ZN => n1195
                           );
   U690 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => OP_B_25_port, ZN => 
                           n1193);
   U691 : INV_X1 port map( A => n1193, ZN => n306);
   U692 : NOR2_X1 port map( A1 => n1195, A2 => n306, ZN => n1164);
   U693 : NOR2_X1 port map( A1 => OP_A_17_port, A2 => OP_B_17_port, ZN => n953)
                           ;
   U694 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => OP_B_17_port, ZN => n951
                           );
   U695 : INV_X1 port map( A => n951, ZN => n928);
   U696 : NOR2_X1 port map( A1 => n953, A2 => n928, ZN => n918);
   U697 : NAND2_X1 port map( A1 => n307, A2 => n451, ZN => n1370);
   U698 : OR4_X1 port map( A1 => n1020, A2 => n1164, A3 => n918, A4 => n1370, 
                           ZN => n312);
   U699 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => OP_B_18_port, ZN => n980
                           );
   U700 : INV_X1 port map( A => n980, ZN => n948);
   U701 : NOR2_X1 port map( A1 => OP_A_18_port, A2 => OP_B_18_port, ZN => n982)
                           ;
   U702 : NOR2_X1 port map( A1 => n948, A2 => n982, ZN => n958);
   U703 : INV_X1 port map( A => n958, ZN => n308);
   U704 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => OP_B_20_port, ZN => 
                           n1046);
   U705 : NOR2_X1 port map( A1 => OP_A_20_port, A2 => OP_B_20_port, ZN => n1049
                           );
   U706 : INV_X1 port map( A => n1049, ZN => n1007);
   U707 : NAND2_X1 port map( A1 => n1046, A2 => n1007, ZN => n1018);
   U708 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => OP_B_22_port, ZN => 
                           n1123);
   U709 : OAI21_X1 port map( B1 => OP_A_22_port, B2 => OP_B_22_port, A => n1123
                           , ZN => n1124);
   U710 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => OP_B_24_port, ZN => 
                           n1192);
   U711 : NOR2_X1 port map( A1 => OP_A_24_port, A2 => OP_B_24_port, ZN => n1194
                           );
   U712 : INV_X1 port map( A => n1194, ZN => n1141);
   U713 : NAND2_X1 port map( A1 => n1192, A2 => n1141, ZN => n1128);
   U714 : NAND4_X1 port map( A1 => n308, A2 => n1018, A3 => n1124, A4 => n1128,
                           ZN => n311);
   U715 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => OP_B_10_port, ZN => n755
                           );
   U716 : OAI21_X1 port map( B1 => OP_A_10_port, B2 => OP_B_10_port, A => n755,
                           ZN => n719);
   U717 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => OP_B_12_port, ZN => n827
                           );
   U718 : NOR2_X1 port map( A1 => OP_A_12_port, A2 => OP_B_12_port, ZN => n830)
                           ;
   U719 : INV_X1 port map( A => n830, ZN => n780);
   U720 : NAND2_X1 port map( A1 => n827, A2 => n780, ZN => n779);
   U721 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => OP_B_14_port, ZN => n870
                           );
   U722 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => OP_B_14_port, A => n870,
                           ZN => n835);
   U723 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => OP_B_16_port, ZN => n949
                           );
   U724 : NOR2_X1 port map( A1 => OP_A_16_port, A2 => OP_B_16_port, ZN => n952)
                           ;
   U725 : INV_X1 port map( A => n952, ZN => n309);
   U726 : NAND2_X1 port map( A1 => n949, A2 => n309, ZN => n904);
   U727 : NAND4_X1 port map( A1 => n719, A2 => n779, A3 => n835, A4 => n904, ZN
                           => n310);
   U728 : NOR4_X1 port map( A1 => n313, A2 => n312, A3 => n311, A4 => n310, ZN 
                           => n314);
   U729 : AOI211_X1 port map( C1 => n315, C2 => n314, A => OP_COMPARE_1_port, B
                           => OP_COMPARE_2_port, ZN => n471);
   U730 : OAI22_X1 port map( A1 => OP_B_0_port, A2 => n316, B1 => OP_B_1_port, 
                           B2 => n578, ZN => n319);
   U731 : OAI21_X1 port map( B1 => OP_B_2_port, B2 => n576, A => n317, ZN => 
                           n368);
   U732 : AOI22_X1 port map( A1 => n365, A2 => n319, B1 => n318, B2 => n368, ZN
                           => n322);
   U733 : OAI21_X1 port map( B1 => n322, B2 => n321, A => n320, ZN => n324);
   U734 : AOI21_X1 port map( B1 => n325, B2 => n324, A => n323, ZN => n362);
   U735 : AOI221_X1 port map( B1 => n362, B2 => n328, C1 => n327, C2 => n328, A
                           => n326, ZN => n329);
   U736 : INV_X1 port map( A => n329, ZN => n463);
   U737 : INV_X1 port map( A => OP_COMPARE_1_port, ZN => n461);
   U738 : OAI211_X1 port map( C1 => n331, C2 => n463, A => n461, B => n330, ZN 
                           => n332);
   U739 : INV_X1 port map( A => n332, ZN => n438);
   U740 : NAND2_X1 port map( A1 => OP_B_14_port, A2 => n333, ZN => n352);
   U741 : INV_X1 port map( A => OP_B_13_port, ZN => n335);
   U742 : AOI222_X1 port map( A1 => OP_A_13_port, A2 => n335, B1 => 
                           OP_A_13_port, B2 => n334, C1 => n335, C2 => n334, ZN
                           => n349);
   U743 : INV_X1 port map( A => n336, ZN => n355);
   U744 : NAND2_X1 port map( A1 => OP_B_10_port, A2 => n337, ZN => n345);
   U745 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n356);
   U746 : AOI211_X1 port map( C1 => n341, C2 => OP_A_9_port, A => n356, B => 
                           n340, ZN => n342);
   U747 : INV_X1 port map( A => n342, ZN => n343);
   U748 : OAI211_X1 port map( C1 => n346, C2 => n345, A => n344, B => n343, ZN 
                           => n348);
   U749 : NOR2_X1 port map( A1 => n353, A2 => n347, ZN => n354);
   U750 : OAI221_X1 port map( B1 => n349, B2 => n355, C1 => n349, C2 => n348, A
                           => n354, ZN => n351);
   U751 : OAI211_X1 port map( C1 => n353, C2 => n352, A => n351, B => n350, ZN 
                           => n389);
   U752 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n357);
   U753 : NOR3_X1 port map( A1 => n358, A2 => n357, A3 => n356, ZN => n383);
   U754 : AOI21_X1 port map( B1 => OP_A_22_port, B2 => n391, A => n410, ZN => 
                           n404);
   U755 : AND2_X1 port map( A1 => n405, A2 => n404, ZN => n360);
   U756 : AOI21_X1 port map( B1 => n359, B2 => OP_A_18_port, A => n399, ZN => 
                           n393);
   U757 : AND4_X1 port map( A1 => n394, A2 => n361, A3 => n360, A4 => n393, ZN 
                           => n387);
   U758 : OAI221_X1 port map( B1 => n389, B2 => n383, C1 => n389, C2 => n362, A
                           => n387, ZN => n445);
   U759 : OAI21_X1 port map( B1 => OP_B_26_port, B2 => n424, A => n423, ZN => 
                           n427);
   U760 : AOI211_X1 port map( C1 => OP_A_24_port, C2 => n418, A => n420, B => 
                           n427, ZN => n440);
   U761 : OAI21_X1 port map( B1 => OP_B_28_port, B2 => n413, A => n363, ZN => 
                           n417);
   U762 : NOR3_X1 port map( A1 => n429, A2 => n441, A3 => n417, ZN => n364);
   U763 : NAND2_X1 port map( A1 => n440, A2 => n364, ZN => n433);
   U764 : OAI21_X1 port map( B1 => n445, B2 => n433, A => OP_COMPARE_1_port, ZN
                           => n436);
   U765 : OAI22_X1 port map( A1 => n368, A2 => n367, B1 => n366, B2 => n365, ZN
                           => n378);
   U766 : NAND2_X1 port map( A1 => OP_B_4_port, A2 => n369, ZN => n371);
   U767 : OAI21_X1 port map( B1 => n372, B2 => n371, A => n370, ZN => n377);
   U768 : AOI21_X1 port map( B1 => OP_A_4_port, B2 => n1362, A => n372, ZN => 
                           n376);
   U769 : OAI21_X1 port map( B1 => OP_B_6_port, B2 => n373, A => n381, ZN => 
                           n374);
   U770 : INV_X1 port map( A => n374, ZN => n375);
   U771 : OAI221_X1 port map( B1 => n378, B2 => n377, C1 => n376, C2 => n377, A
                           => n375, ZN => n386);
   U772 : NOR2_X1 port map( A1 => OP_A_6_port, A2 => n379, ZN => n382);
   U773 : AOI21_X1 port map( B1 => n382, B2 => n381, A => n380, ZN => n385);
   U774 : INV_X1 port map( A => n383, ZN => n384);
   U775 : AOI21_X1 port map( B1 => n386, B2 => n385, A => n384, ZN => n388);
   U776 : OAI21_X1 port map( B1 => n389, B2 => n388, A => n387, ZN => n390);
   U777 : INV_X1 port map( A => n390, ZN => n444);
   U778 : OR2_X1 port map( A1 => OP_A_22_port, A2 => n391, ZN => n411);
   U779 : NAND2_X1 port map( A1 => n392, A2 => OP_B_18_port, ZN => n400);
   U780 : OAI211_X1 port map( C1 => n396, C2 => n395, A => n394, B => n393, ZN 
                           => n397);
   U781 : OAI211_X1 port map( C1 => n400, C2 => n399, A => n398, B => n397, ZN 
                           => n407);
   U782 : INV_X1 port map( A => n401, ZN => n402);
   U783 : OAI222_X1 port map( A1 => n403, A2 => n402, B1 => n403, B2 => 
                           OP_A_21_port, C1 => n402, C2 => OP_A_21_port, ZN => 
                           n406);
   U784 : OAI221_X1 port map( B1 => n407, B2 => n406, C1 => n405, C2 => n406, A
                           => n404, ZN => n408);
   U785 : OAI211_X1 port map( C1 => n411, C2 => n410, A => n409, B => n408, ZN 
                           => n456);
   U786 : INV_X1 port map( A => n456, ZN => n434);
   U787 : AOI21_X1 port map( B1 => n412, B2 => n451, A => n454, ZN => n432);
   U788 : NAND2_X1 port map( A1 => OP_B_28_port, A2 => n413, ZN => n415);
   U789 : OAI21_X1 port map( B1 => n416, B2 => n415, A => n414, ZN => n450);
   U790 : INV_X1 port map( A => n417, ZN => n449);
   U791 : OR2_X1 port map( A1 => OP_A_24_port, A2 => n418, ZN => n421);
   U792 : OAI21_X1 port map( B1 => n421, B2 => n420, A => n419, ZN => n422);
   U793 : INV_X1 port map( A => n422, ZN => n428);
   U794 : NAND3_X1 port map( A1 => OP_B_26_port, A2 => n424, A3 => n423, ZN => 
                           n425);
   U795 : OAI211_X1 port map( C1 => n428, C2 => n427, A => n426, B => n425, ZN 
                           => n448);
   U796 : NOR2_X1 port map( A1 => n429, A2 => n441, ZN => n430);
   U797 : OAI221_X1 port map( B1 => n450, B2 => n449, C1 => n450, C2 => n448, A
                           => n430, ZN => n431);
   U798 : OAI211_X1 port map( C1 => n434, C2 => n433, A => n432, B => n431, ZN 
                           => n435);
   U799 : AOI221_X1 port map( B1 => OP_COMPARE_2_port, B2 => n436, C1 => n444, 
                           C2 => n436, A => n435, ZN => n437);
   U800 : OAI21_X1 port map( B1 => n438, B2 => n437, A => OP_COMPARE_0_port, ZN
                           => n470);
   U801 : INV_X1 port map( A => n439, ZN => n468);
   U802 : INV_X1 port map( A => n440, ZN => n443);
   U803 : NOR2_X1 port map( A1 => n454, A2 => n441, ZN => n447);
   U804 : NAND2_X1 port map( A1 => n449, A2 => n447, ZN => n442);
   U805 : NOR2_X1 port map( A1 => n443, A2 => n442, ZN => n457);
   U806 : AOI21_X1 port map( B1 => n444, B2 => n457, A => OP_COMPARE_2_port, ZN
                           => n460);
   U807 : INV_X1 port map( A => n445, ZN => n446);
   U808 : AOI21_X1 port map( B1 => n446, B2 => n457, A => n461, ZN => n459);
   U809 : OAI221_X1 port map( B1 => n450, B2 => n449, C1 => n450, C2 => n448, A
                           => n447, ZN => n452);
   U810 : OAI211_X1 port map( C1 => n454, C2 => n453, A => n452, B => n451, ZN 
                           => n455);
   U811 : AOI21_X1 port map( B1 => n457, B2 => n456, A => n455, ZN => n458);
   U812 : OAI21_X1 port map( B1 => n460, B2 => n459, A => n458, ZN => n466);
   U813 : OAI211_X1 port map( C1 => n464, C2 => n463, A => n462, B => n461, ZN 
                           => n465);
   U814 : AOI21_X1 port map( B1 => n466, B2 => n465, A => OP_COMPARE_0_port, ZN
                           => n467);
   U815 : OAI21_X1 port map( B1 => n471, B2 => n468, A => n467, ZN => n469);
   U816 : OAI21_X1 port map( B1 => n471, B2 => n470, A => n469, ZN => n473);
   U817 : INV_X1 port map( A => N285, ZN => n472);
   U818 : AOI221_X1 port map( B1 => OP_COMPARE_3_port, B2 => n475, C1 => n474, 
                           C2 => n473, A => n472, ZN => n480);
   U819 : INV_X1 port map( A => N279, ZN => n1397);
   U820 : XOR2_X1 port map( A => n477, B => OP_Ci, Z => n478);
   U821 : NAND2_X1 port map( A1 => OP_LOGIC_1_port, A2 => n476, ZN => n1371);
   U822 : OAI22_X1 port map( A1 => n1397, A2 => n478, B1 => n1371, B2 => n477, 
                           ZN => n479);
   U823 : AOI211_X1 port map( C1 => n1366, C2 => n489, A => n480, B => n479, ZN
                           => n481);
   U824 : OAI211_X1 port map( C1 => n1158, C2 => n483, A => n482, B => n481, ZN
                           => Y(0));
   U825 : INV_X1 port map( A => n508, ZN => n484);
   U826 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_1, A => n484, 
                           ZN => n486);
   U827 : OAI22_X1 port map( A1 => n1395, A2 => n486, B1 => n1138, B2 => n485, 
                           ZN => n488);
   U828 : AOI22_X1 port map( A1 => n56, A2 => OP_A_0_port, B1 => OP_A_1_port, 
                           B2 => n57, ZN => n920);
   U829 : OAI22_X1 port map( A1 => n920, A2 => n1061, B1 => n520, B2 => n1368, 
                           ZN => n487);
   U830 : AOI211_X1 port map( C1 => n1329, C2 => OP1(1), A => n488, B => n487, 
                           ZN => n505);
   U831 : AOI22_X1 port map( A1 => OP_B_0_port, A2 => OP_A_0_port, B1 => OP_Ci,
                           B2 => n489, ZN => n522);
   U832 : INV_X1 port map( A => n522, ZN => n491);
   U833 : INV_X1 port map( A => n506, ZN => n490);
   U834 : AOI221_X1 port map( B1 => n522, B2 => n506, C1 => n491, C2 => n490, A
                           => n1397, ZN => n502);
   U835 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n55, ZN => n1352);
   U836 : NAND2_X1 port map( A1 => n56, A2 => OP_A_26_port, ZN => n1225);
   U837 : NAND2_X1 port map( A1 => OP_A_27_port, A2 => n553, ZN => n1288);
   U838 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => n57, ZN => n1165);
   U839 : NAND4_X1 port map( A1 => n1352, A2 => n1225, A3 => n1288, A4 => n1165
                           , ZN => n791);
   U840 : NAND2_X1 port map( A1 => n56, A2 => OP_A_30_port, ZN => n1353);
   U841 : NAND2_X1 port map( A1 => OP_A_29_port, A2 => n57, ZN => n1289);
   U842 : OAI211_X1 port map( C1 => n575, C2 => n1369, A => n1353, B => n1289, 
                           ZN => n492);
   U843 : AOI21_X1 port map( B1 => OP_SHIFT, B2 => n55, A => n492, ZN => n1297)
                           ;
   U844 : INV_X1 port map( A => n1297, ZN => n797);
   U845 : AOI22_X1 port map( A1 => n855, A2 => n791, B1 => n511, B2 => n797, ZN
                           => n494);
   U846 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => n55, ZN => n1224);
   U847 : NAND2_X1 port map( A1 => n56, A2 => OP_A_22_port, ZN => n1097);
   U848 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => n553, ZN => n1168);
   U849 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => n57, ZN => n1033);
   U850 : NAND4_X1 port map( A1 => n1224, A2 => n1097, A3 => n1168, A4 => n1033
                           , ZN => n792);
   U851 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => n55, ZN => n1096);
   U852 : NAND2_X1 port map( A1 => n56, A2 => OP_A_18_port, ZN => n971);
   U853 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => n553, ZN => n1036);
   U854 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n57, ZN => n912);
   U855 : NAND4_X1 port map( A1 => n1096, A2 => n971, A3 => n1036, A4 => n912, 
                           ZN => n794);
   U856 : AOI22_X1 port map( A1 => n66, A2 => n792, B1 => n894, B2 => n794, ZN 
                           => n493);
   U857 : NAND2_X1 port map( A1 => n494, A2 => n493, ZN => n922);
   U858 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => n55, ZN => n738);
   U859 : NAND2_X1 port map( A1 => OP_A_7_port, A2 => n553, ZN => n693);
   U860 : NAND2_X1 port map( A1 => OP_A_5_port, A2 => n57, ZN => n495);
   U861 : NAND4_X1 port map( A1 => n738, A2 => n658, A3 => n693, A4 => n495, ZN
                           => n596);
   U862 : AOI22_X1 port map( A1 => OP_B_4_port, A2 => n922, B1 => n1357, B2 => 
                           n596, ZN => n500);
   U863 : NAND2_X1 port map( A1 => OP_A_4_port, A2 => n55, ZN => n656);
   U864 : NAND2_X1 port map( A1 => OP_A_1_port, A2 => n57, ZN => n496);
   U865 : OAI211_X1 port map( C1 => n575, C2 => n550, A => n656, B => n496, ZN 
                           => n498);
   U866 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n55, ZN => n970);
   U867 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => n57, ZN => n802);
   U868 : NAND2_X1 port map( A1 => OP_A_15_port, A2 => n553, ZN => n915);
   U869 : NAND4_X1 port map( A1 => n852, A2 => n970, A3 => n802, A4 => n915, ZN
                           => n609);
   U870 : INV_X1 port map( A => n609, ZN => n795);
   U871 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => n55, ZN => n850);
   U872 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => n553, ZN => n803);
   U873 : NAND2_X1 port map( A1 => OP_A_9_port, A2 => n57, ZN => n694);
   U874 : AND4_X1 port map( A1 => n850, A2 => n740, A3 => n803, A4 => n694, ZN 
                           => n699);
   U875 : OAI22_X1 port map( A1 => n795, A2 => n891, B1 => n699, B2 => n566, ZN
                           => n497);
   U876 : AOI221_X1 port map( B1 => n552, B2 => n1359, C1 => n498, C2 => n1359,
                           A => n497, ZN => n499);
   U877 : AOI21_X1 port map( B1 => n500, B2 => n499, A => n1158, ZN => n501);
   U878 : AOI211_X1 port map( C1 => n1366, C2 => n503, A => n502, B => n501, ZN
                           => n504);
   U879 : OAI211_X1 port map( C1 => n1371, C2 => n506, A => n505, B => n504, ZN
                           => Y(1));
   U880 : INV_X1 port map( A => n1371, ZN => n1343);
   U881 : INV_X1 port map( A => n524, ZN => n523);
   U882 : AOI22_X1 port map( A1 => n507, A2 => n1244, B1 => n1343, B2 => n523, 
                           ZN => n534);
   U883 : INV_X1 port map( A => n1138, ZN => n1347);
   U884 : NAND2_X1 port map( A1 => OP_A_2_port, A2 => n57, ZN => n516);
   U885 : OAI211_X1 port map( C1 => n575, C2 => n549, A => n508, B => n516, ZN 
                           => n820);
   U886 : AOI22_X1 port map( A1 => n1347, A2 => OP2(2), B1 => n1227, B2 => n820
                           , ZN => n533);
   U887 : AOI22_X1 port map( A1 => OP1(2), A2 => n1329, B1 => n1366, B2 => n546
                           , ZN => n532);
   U888 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => n57, ZN => n816);
   U889 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n603, ZN => n938);
   U890 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n55, ZN => n1003);
   U891 : NAND4_X1 port map( A1 => n890, A2 => n816, A3 => n938, A4 => n1003, 
                           ZN => n841);
   U892 : INV_X1 port map( A => n841, ZN => n728);
   U893 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => n603, ZN => n723);
   U894 : NAND2_X1 port map( A1 => OP_A_6_port, A2 => n57, ZN => n625);
   U895 : NAND2_X1 port map( A1 => OP_A_9_port, A2 => n55, ZN => n766);
   U896 : NAND4_X1 port map( A1 => n723, A2 => n625, A3 => n766, A4 => n675, ZN
                           => n618);
   U897 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => n603, ZN => n818);
   U898 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => n57, ZN => n724);
   U899 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => n55, ZN => n888);
   U900 : NAND4_X1 port map( A1 => n818, A2 => n724, A3 => n769, A4 => n888, ZN
                           => n721);
   U901 : AOI22_X1 port map( A1 => n1357, A2 => n618, B1 => n1349, B2 => n721, 
                           ZN => n519);
   U902 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => n603, ZN => n1205);
   U903 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => n57, ZN => n1056);
   U904 : NAND2_X1 port map( A1 => n56, A2 => OP_A_23_port, ZN => n1131);
   U905 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => n55, ZN => n1269);
   U906 : AND4_X1 port map( A1 => n1205, A2 => n1056, A3 => n1131, A4 => n1269,
                           ZN => n824);
   U907 : AOI22_X1 port map( A1 => OP_B_1_port, A2 => OP_SHIFT, B1 => 
                           OP_A_30_port, B2 => n57, ZN => n509);
   U908 : OAI21_X1 port map( B1 => n510, B2 => n1369, A => n509, ZN => n1327);
   U909 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => n603, ZN => n1059);
   U910 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => n57, ZN => n935);
   U911 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => n55, ZN => n1130);
   U912 : NAND2_X1 port map( A1 => n56, A2 => OP_A_19_port, ZN => n1004);
   U913 : NAND4_X1 port map( A1 => n1059, A2 => n935, A3 => n1130, A4 => n1004,
                           ZN => n826);
   U914 : AOI22_X1 port map( A1 => n511, A2 => n1327, B1 => n894, B2 => n826, 
                           ZN => n514);
   U915 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => n57, ZN => n1202);
   U916 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n553, ZN => n1319);
   U917 : NAND2_X1 port map( A1 => n56, A2 => OP_A_27_port, ZN => n1270);
   U918 : NAND2_X1 port map( A1 => OP_A_29_port, A2 => n55, ZN => n512);
   U919 : NAND4_X1 port map( A1 => n1202, A2 => n1319, A3 => n1270, A4 => n512,
                           ZN => n837);
   U920 : NAND2_X1 port map( A1 => n855, A2 => n837, ZN => n513);
   U921 : OAI211_X1 port map( C1 => n824, C2 => n742, A => n514, B => n513, ZN 
                           => n934);
   U922 : NAND2_X1 port map( A1 => OP_A_4_port, A2 => n553, ZN => n627);
   U923 : INV_X1 port map( A => n580, ZN => n515);
   U924 : NAND2_X1 port map( A1 => OP_A_5_port, A2 => n55, ZN => n673);
   U925 : NAND4_X1 port map( A1 => n627, A2 => n516, A3 => n515, A4 => n673, ZN
                           => n517);
   U926 : AOI22_X1 port map( A1 => OP_B_4_port, A2 => n934, B1 => n1359, B2 => 
                           n517, ZN => n518);
   U927 : OAI211_X1 port map( C1 => n728, C2 => n891, A => n519, B => n518, ZN 
                           => n530);
   U928 : OAI21_X1 port map( B1 => n522, B2 => n521, A => n520, ZN => n547);
   U929 : INV_X1 port map( A => n547, ZN => n525);
   U930 : AOI221_X1 port map( B1 => n525, B2 => n524, C1 => n547, C2 => n523, A
                           => n1397, ZN => n529);
   U931 : AOI211_X1 port map( C1 => n527, C2 => n526, A => n538, B => n1395, ZN
                           => n528);
   U932 : AOI211_X1 port map( C1 => N284, C2 => n530, A => n529, B => n528, ZN 
                           => n531);
   U933 : NAND4_X1 port map( A1 => n534, A2 => n533, A3 => n532, A4 => n531, ZN
                           => Y(2));
   U934 : XNOR2_X1 port map( A => n536, B => n535, ZN => n537);
   U935 : XNOR2_X1 port map( A => n538, B => n537, ZN => n563);
   U936 : INV_X1 port map( A => n1395, ZN => n986);
   U937 : INV_X1 port map( A => n986, ZN => n1283);
   U938 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => n553, ZN => n1226);
   U939 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => n57, ZN => n1095);
   U940 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => n55, ZN => n1286);
   U941 : NAND2_X1 port map( A1 => n56, A2 => OP_A_24_port, ZN => n1167);
   U942 : NAND4_X1 port map( A1 => n1226, A2 => n1095, A3 => n1286, A4 => n1167
                           , ZN => n863);
   U943 : NAND2_X1 port map( A1 => OP_A_29_port, A2 => n553, ZN => n1354);
   U944 : NAND2_X1 port map( A1 => OP_A_27_port, A2 => n57, ZN => n1223);
   U945 : NAND2_X1 port map( A1 => n56, A2 => OP_A_28_port, ZN => n1287);
   U946 : NAND3_X1 port map( A1 => n1354, A2 => n1223, A3 => n1287, ZN => n539)
                           ;
   U947 : AOI21_X1 port map( B1 => OP_A_30_port, B2 => n55, A => n539, ZN => 
                           n869);
   U948 : NOR2_X1 port map( A1 => n869, A2 => n741, ZN => n541);
   U949 : AOI22_X1 port map( A1 => n57, A2 => OP_A_31_port, B1 => OP_SHIFT, B2 
                           => n607, ZN => n1373);
   U950 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => n553, ZN => n1098);
   U951 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => n57, ZN => n969);
   U952 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => n55, ZN => n1166);
   U953 : NAND2_X1 port map( A1 => n56, A2 => OP_A_20_port, ZN => n1035);
   U954 : NAND4_X1 port map( A1 => n1098, A2 => n969, A3 => n1166, A4 => n1035,
                           ZN => n865);
   U955 : INV_X1 port map( A => n865, ZN => n748);
   U956 : OAI22_X1 port map( A1 => n1373, A2 => n857, B1 => n748, B2 => n765, 
                           ZN => n540);
   U957 : NAND2_X1 port map( A1 => OP_A_9_port, A2 => n553, ZN => n737);
   U958 : NAND2_X1 port map( A1 => OP_A_7_port, A2 => n57, ZN => n655);
   U959 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => n55, ZN => n801);
   U960 : NAND4_X1 port map( A1 => n737, A2 => n655, A3 => n801, A4 => n696, ZN
                           => n648);
   U961 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => n553, ZN => n851);
   U962 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => n57, ZN => n739);
   U963 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => n55, ZN => n913);
   U964 : NAND4_X1 port map( A1 => n851, A2 => n739, A3 => n804, A4 => n913, ZN
                           => n644);
   U965 : AOI22_X1 port map( A1 => n1357, A2 => n648, B1 => n1349, B2 => n644, 
                           ZN => n545);
   U966 : NAND2_X1 port map( A1 => OP_A_5_port, A2 => n553, ZN => n657);
   U967 : NAND2_X1 port map( A1 => OP_A_3_port, A2 => n57, ZN => n542);
   U968 : NAND2_X1 port map( A1 => OP_A_6_port, A2 => n55, ZN => n695);
   U969 : NAND4_X1 port map( A1 => n657, A2 => n542, A3 => n695, A4 => n604, ZN
                           => n543);
   U970 : NAND2_X1 port map( A1 => OP_A_15_port, A2 => n57, ZN => n849);
   U971 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n553, ZN => n972);
   U972 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => n55, ZN => n1034);
   U973 : NAND2_X1 port map( A1 => n56, A2 => OP_A_16_port, ZN => n914);
   U974 : NAND4_X1 port map( A1 => n849, A2 => n972, A3 => n1034, A4 => n914, 
                           ZN => n874);
   U975 : AOI22_X1 port map( A1 => n1359, A2 => n543, B1 => n1351, B2 => n874, 
                           ZN => n544);
   U976 : OAI211_X1 port map( C1 => n964, C2 => n1362, A => n545, B => n544, ZN
                           => n560);
   U977 : AOI22_X1 port map( A1 => OP_B_2_port, A2 => OP_A_2_port, B1 => n547, 
                           B2 => n546, ZN => n548);
   U978 : NOR2_X1 port map( A1 => n557, A2 => n548, ZN => n571);
   U979 : AOI211_X1 port map( C1 => n557, C2 => n548, A => n1397, B => n571, ZN
                           => n559);
   U980 : AOI22_X1 port map( A1 => n1347, A2 => OP2(3), B1 => n1346, B2 => 
                           OP1(3), ZN => n556);
   U981 : OAI22_X1 port map( A1 => n550, A2 => n607, B1 => n549, B2 => n577, ZN
                           => n551);
   U982 : AOI211_X1 port map( C1 => n553, C2 => OP_A_1_port, A => n552, B => 
                           n551, ZN => n966);
   U983 : INV_X1 port map( A => n966, ZN => n554);
   U984 : AOI22_X1 port map( A1 => OP_B_3_port, A2 => n1366, B1 => n1227, B2 =>
                           n554, ZN => n555);
   U985 : OAI211_X1 port map( C1 => n557, C2 => n1371, A => n556, B => n555, ZN
                           => n558);
   U986 : AOI211_X1 port map( C1 => N284, C2 => n560, A => n559, B => n558, ZN 
                           => n562);
   U987 : OAI221_X1 port map( B1 => n1366, B2 => OP_B_3_port, C1 => n1366, C2 
                           => n1244, A => OP_A_3_port, ZN => n561);
   U988 : OAI211_X1 port map( C1 => n563, C2 => n1283, A => n562, B => n561, ZN
                           => Y(3));
   U989 : NAND2_X1 port map( A1 => n1351, A2 => N284, ZN => n868);
   U990 : INV_X1 port map( A => n868, ZN => n838);
   U991 : AOI211_X1 port map( C1 => n565, C2 => intadd_0_SUM_0_port, A => n564,
                           B => n1395, ZN => n568);
   U992 : NOR2_X1 port map( A1 => n1158, A2 => n566, ZN => n864);
   U993 : INV_X1 port map( A => n864, ZN => n823);
   U994 : NOR2_X1 port map( A1 => n1158, A2 => n899, ZN => n866);
   U995 : INV_X1 port map( A => n866, ZN => n727);
   U996 : OAI22_X1 port map( A1 => n771, A2 => n823, B1 => n681, B2 => n727, ZN
                           => n567);
   U997 : AOI211_X1 port map( C1 => n838, C2 => n777, A => n568, B => n567, ZN 
                           => n589);
   U998 : INV_X1 port map( A => n573, ZN => n572);
   U999 : NAND2_X1 port map( A1 => OP_B_4_port, A2 => N284, ZN => n764);
   U1000 : INV_X1 port map( A => n764, ZN => n744);
   U1001 : AOI22_X1 port map( A1 => n855, A2 => n1264, B1 => n65, B2 => n781, 
                           ZN => n569);
   U1002 : INV_X1 port map( A => OP_SHIFT, ZN => n1157);
   U1003 : NOR2_X1 port map( A1 => n857, A2 => n1157, ZN => n660);
   U1004 : INV_X1 port map( A => n660, ZN => n623);
   U1005 : OAI211_X1 port map( C1 => n784, C2 => n765, A => n569, B => n623, ZN
                           => n1008);
   U1006 : AOI22_X1 port map( A1 => n1343, A2 => n572, B1 => n744, B2 => n1008,
                           ZN => n588);
   U1007 : INV_X1 port map( A => n570, ZN => n598);
   U1008 : AOI22_X1 port map( A1 => n1244, A2 => n598, B1 => n1366, B2 => n597,
                           ZN => n587);
   U1009 : AOI21_X1 port map( B1 => OP_A_3_port, B2 => OP_B_3_port, A => n571, 
                           ZN => n574);
   U1010 : INV_X1 port map( A => n574, ZN => n599);
   U1011 : AOI221_X1 port map( B1 => n574, B2 => n573, C1 => n599, C2 => n572, 
                           A => n1397, ZN => n585);
   U1012 : OAI22_X1 port map( A1 => n578, A2 => n577, B1 => n576, B2 => n575, 
                           ZN => n579);
   U1013 : AOI211_X1 port map( C1 => n57, C2 => OP_A_4_port, A => n580, B => 
                           n579, ZN => n892);
   U1014 : AOI22_X1 port map( A1 => OP_B_2_port, A2 => n895, B1 => n892, B2 => 
                           n581, ZN => n770);
   U1015 : NAND2_X1 port map( A1 => n770, A2 => n1159, ZN => n1011);
   U1016 : NAND2_X1 port map( A1 => n1362, A2 => n1365, ZN => n885);
   U1017 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n1158, ZN => n1251);
   U1018 : NAND2_X1 port map( A1 => n894, A2 => n1251, ZN => n1372);
   U1019 : INV_X1 port map( A => n1372, ZN => n1328);
   U1020 : AOI22_X1 port map( A1 => n1329, A2 => OP1(4), B1 => n1328, B2 => 
                           n582, ZN => n583);
   U1021 : OAI21_X1 port map( B1 => n1011, B2 => n885, A => n583, ZN => n584);
   U1022 : AOI211_X1 port map( C1 => n1347, C2 => OP2(4), A => n585, B => n584,
                           ZN => n586);
   U1023 : NAND4_X1 port map( A1 => n589, A2 => n588, A3 => n587, A4 => n586, 
                           ZN => Y(4));
   U1024 : XNOR2_X1 port map( A => n591, B => n590, ZN => n592);
   U1025 : XNOR2_X1 port map( A => intadd_0_SUM_1_port, B => n592, ZN => n617);
   U1026 : INV_X1 port map( A => n794, ZN => n703);
   U1027 : OAI22_X1 port map( A1 => n703, A2 => n868, B1 => n699, B2 => n727, 
                           ZN => n595);
   U1028 : OAI22_X1 port map( A1 => n593, A2 => n1368, B1 => n1371, B2 => n600,
                           ZN => n594);
   U1029 : AOI211_X1 port map( C1 => n1328, C2 => n596, A => n595, B => n594, 
                           ZN => n616);
   U1030 : OAI21_X1 port map( B1 => n599, B2 => n598, A => n597, ZN => n601);
   U1031 : INV_X1 port map( A => n601, ZN => n633);
   U1032 : INV_X1 port map( A => n600, ZN => n602);
   U1033 : AOI221_X1 port map( B1 => n633, B2 => n602, C1 => n601, C2 => n600, 
                           A => n1397, ZN => n614);
   U1034 : INV_X1 port map( A => n885, ZN => n743);
   U1035 : AOI22_X1 port map( A1 => OP_A_3_port, A2 => n603, B1 => OP_A_2_port,
                           B2 => n55, ZN => n605);
   U1036 : OAI211_X1 port map( C1 => n607, C2 => n606, A => n605, B => n604, ZN
                           => n919);
   U1037 : INV_X1 port map( A => n919, ZN => n697);
   U1038 : OAI22_X1 port map( A1 => n697, A2 => n765, B1 => n920, B2 => n742, 
                           ZN => n1029);
   U1039 : AOI22_X1 port map( A1 => n1329, A2 => OP1(5), B1 => n743, B2 => 
                           n1029, ZN => n611);
   U1040 : AOI22_X1 port map( A1 => n853, A2 => n791, B1 => n894, B2 => n792, 
                           ZN => n608);
   U1041 : OAI211_X1 port map( C1 => n1297, C2 => n741, A => n608, B => n623, 
                           ZN => n1038);
   U1042 : AOI22_X1 port map( A1 => n744, A2 => n1038, B1 => n864, B2 => n609, 
                           ZN => n610);
   U1043 : OAI211_X1 port map( C1 => n1138, C2 => n612, A => n611, B => n610, 
                           ZN => n613);
   U1044 : AOI211_X1 port map( C1 => n1366, C2 => n632, A => n614, B => n613, 
                           ZN => n615);
   U1045 : OAI211_X1 port map( C1 => n1283, C2 => n617, A => n616, B => n615, 
                           ZN => Y(5));
   U1046 : INV_X1 port map( A => n636, ZN => n634);
   U1047 : AOI22_X1 port map( A1 => n1328, A2 => n618, B1 => n1343, B2 => n634,
                           ZN => n640);
   U1048 : AOI211_X1 port map( C1 => n620, C2 => intadd_1_SUM_0_port, A => n619
                           , B => n1395, ZN => n622);
   U1049 : OAI22_X1 port map( A1 => n651, A2 => n1367, B1 => n728, B2 => n823, 
                           ZN => n621);
   U1050 : AOI211_X1 port map( C1 => n866, C2 => n721, A => n622, B => n621, ZN
                           => n639);
   U1051 : AOI22_X1 port map( A1 => n855, A2 => n1327, B1 => n66, B2 => n837, 
                           ZN => n624);
   U1052 : OAI211_X1 port map( C1 => n824, C2 => n765, A => n624, B => n623, ZN
                           => n1065);
   U1053 : NAND4_X1 port map( A1 => n628, A2 => n627, A3 => n626, A4 => n625, 
                           ZN => n940);
   U1054 : AOI22_X1 port map( A1 => n65, A2 => n820, B1 => n894, B2 => n940, ZN
                           => n1062);
   U1055 : AOI22_X1 port map( A1 => n1347, A2 => OP2(6), B1 => n1329, B2 => 
                           OP1(6), ZN => n629);
   U1056 : OAI21_X1 port map( B1 => n1062, B2 => n885, A => n629, ZN => n631);
   U1057 : INV_X1 port map( A => n826, ZN => n729);
   U1058 : OAI22_X1 port map( A1 => n729, A2 => n868, B1 => n649, B2 => n1368, 
                           ZN => n630);
   U1059 : AOI211_X1 port map( C1 => n744, C2 => n1065, A => n631, B => n630, 
                           ZN => n638);
   U1060 : AOI22_X1 port map( A1 => OP_B_5_port, A2 => OP_A_5_port, B1 => n633,
                           B2 => n632, ZN => n650);
   U1061 : INV_X1 port map( A => n650, ZN => n635);
   U1062 : OAI221_X1 port map( B1 => n650, B2 => n636, C1 => n635, C2 => n634, 
                           A => N279, ZN => n637);
   U1063 : NAND4_X1 port map( A1 => n640, A2 => n639, A3 => n638, A4 => n637, 
                           ZN => Y(6));
   U1064 : XNOR2_X1 port map( A => n642, B => n641, ZN => n643);
   U1065 : XNOR2_X1 port map( A => intadd_1_SUM_1_port, B => n643, ZN => n669);
   U1066 : INV_X1 port map( A => n644, ZN => n747);
   U1067 : OAI22_X1 port map( A1 => n748, A2 => n868, B1 => n747, B2 => n727, 
                           ZN => n647);
   U1068 : OAI22_X1 port map( A1 => n645, A2 => n1368, B1 => n1371, B2 => n653,
                           ZN => n646);
   U1069 : AOI211_X1 port map( C1 => n1328, C2 => n648, A => n647, B => n646, 
                           ZN => n668);
   U1070 : OAI21_X1 port map( B1 => n651, B2 => n650, A => n649, ZN => n677);
   U1071 : INV_X1 port map( A => n677, ZN => n654);
   U1072 : INV_X1 port map( A => n653, ZN => n652);
   U1073 : AOI221_X1 port map( B1 => n654, B2 => n653, C1 => n677, C2 => n652, 
                           A => n1397, ZN => n666);
   U1074 : NAND4_X1 port map( A1 => n658, A2 => n657, A3 => n656, A4 => n655, 
                           ZN => n854);
   U1075 : INV_X1 port map( A => n854, ZN => n963);
   U1076 : OAI22_X1 port map( A1 => n963, A2 => n765, B1 => n966, B2 => n742, 
                           ZN => n1099);
   U1077 : AOI22_X1 port map( A1 => n1329, A2 => OP1(7), B1 => n743, B2 => 
                           n1099, ZN => n663);
   U1078 : OAI22_X1 port map( A1 => n1373, A2 => n741, B1 => n869, B2 => n742, 
                           ZN => n659);
   U1079 : AOI211_X1 port map( C1 => n894, C2 => n863, A => n660, B => n659, ZN
                           => n1106);
   U1080 : INV_X1 port map( A => n1106, ZN => n661);
   U1081 : AOI22_X1 port map( A1 => n744, A2 => n661, B1 => n864, B2 => n874, 
                           ZN => n662);
   U1082 : OAI211_X1 port map( C1 => n1138, C2 => n664, A => n663, B => n662, 
                           ZN => n665);
   U1083 : AOI211_X1 port map( C1 => n1366, C2 => n678, A => n666, B => n665, 
                           ZN => n667);
   U1084 : OAI211_X1 port map( C1 => n1283, C2 => n669, A => n668, B => n667, 
                           ZN => Y(7));
   U1085 : AOI22_X1 port map( A1 => n66, A2 => n1264, B1 => n894, B2 => n781, 
                           ZN => n670);
   U1086 : OAI21_X1 port map( B1 => n1159, B2 => n1157, A => n670, ZN => n1134)
                           ;
   U1087 : AOI22_X1 port map( A1 => n744, A2 => n1134, B1 => n1366, B2 => n671,
                           ZN => n690);
   U1088 : INV_X1 port map( A => n711, ZN => n676);
   U1089 : NAND4_X1 port map( A1 => n675, A2 => n674, A3 => n673, A4 => n672, 
                           ZN => n1006);
   U1090 : INV_X1 port map( A => n1006, ZN => n905);
   U1091 : OAI222_X1 port map( A1 => n895, A2 => n741, B1 => n765, B2 => n905, 
                           C1 => n742, C2 => n892, ZN => n1133);
   U1092 : AOI22_X1 port map( A1 => n676, A2 => n1244, B1 => n743, B2 => n1133,
                           ZN => n689);
   U1093 : AOI22_X1 port map( A1 => OP_B_7_port, A2 => OP_A_7_port, B1 => n678,
                           B2 => n677, ZN => n712);
   U1094 : NOR2_X1 port map( A1 => n712, A2 => n680, ZN => n679);
   U1095 : AOI211_X1 port map( C1 => n712, C2 => n680, A => n1397, B => n679, 
                           ZN => n687);
   U1096 : OAI22_X1 port map( A1 => n681, A2 => n1372, B1 => n680, B2 => n1371,
                           ZN => n686);
   U1097 : AOI22_X1 port map( A1 => n1347, A2 => OP2(8), B1 => n1329, B2 => 
                           OP1(8), ZN => n684);
   U1098 : OAI22_X1 port map( A1 => n784, A2 => n868, B1 => n771, B2 => n727, 
                           ZN => n682);
   U1099 : AOI21_X1 port map( B1 => n864, B2 => n777, A => n682, ZN => n683);
   U1100 : OAI211_X1 port map( C1 => intadd_2_SUM_0_port, C2 => n1283, A => 
                           n684, B => n683, ZN => n685);
   U1101 : NOR3_X1 port map( A1 => n687, A2 => n686, A3 => n685, ZN => n688);
   U1102 : NAND3_X1 port map( A1 => n690, A2 => n689, A3 => n688, ZN => Y(8));
   U1103 : OAI22_X1 port map( A1 => intadd_2_SUM_1_port, A2 => n1283, B1 => 
                           n1138, B2 => n691, ZN => n692);
   U1104 : AOI21_X1 port map( B1 => n702, B2 => n1343, A => n692, ZN => n710);
   U1105 : NAND4_X1 port map( A1 => n696, A2 => n695, A3 => n694, A4 => n693, 
                           ZN => n1037);
   U1106 : INV_X1 port map( A => n1037, ZN => n931);
   U1107 : OAI222_X1 port map( A1 => n742, A2 => n697, B1 => n765, B2 => n931, 
                           C1 => n741, C2 => n920, ZN => n1160);
   U1108 : AOI22_X1 port map( A1 => n1329, A2 => OP1(9), B1 => n743, B2 => 
                           n1160, ZN => n709);
   U1109 : NOR2_X1 port map( A1 => n1157, A2 => n764, ZN => n1120);
   U1110 : INV_X1 port map( A => n1120, ZN => n1108);
   U1111 : NOR2_X1 port map( A1 => n1159, A2 => n1108, ZN => n753);
   U1112 : INV_X1 port map( A => n698, ZN => n713);
   U1113 : OAI22_X1 port map( A1 => n699, A2 => n1372, B1 => n713, B2 => n1368,
                           ZN => n700);
   U1114 : AOI211_X1 port map( C1 => n838, C2 => n792, A => n753, B => n700, ZN
                           => n708);
   U1115 : AOI21_X1 port map( B1 => n712, B2 => n711, A => n715, ZN => n701);
   U1116 : XOR2_X1 port map( A => n702, B => n701, Z => n706);
   U1117 : OAI22_X1 port map( A1 => n703, A2 => n823, B1 => n714, B2 => n1367, 
                           ZN => n705);
   U1118 : AOI22_X1 port map( A1 => n853, A2 => n797, B1 => n894, B2 => n791, 
                           ZN => n1173);
   U1119 : OAI22_X1 port map( A1 => n1173, A2 => n764, B1 => n795, B2 => n727, 
                           ZN => n704);
   U1120 : AOI211_X1 port map( C1 => n706, C2 => N279, A => n705, B => n704, ZN
                           => n707);
   U1121 : NAND4_X1 port map( A1 => n710, A2 => n709, A3 => n708, A4 => n707, 
                           ZN => Y(9));
   U1122 : NAND2_X1 port map( A1 => n713, A2 => n711, ZN => n718);
   U1123 : INV_X1 port map( A => n712, ZN => n717);
   U1124 : OAI21_X1 port map( B1 => n715, B2 => n714, A => n713, ZN => n716);
   U1125 : OAI21_X1 port map( B1 => n718, B2 => n717, A => n716, ZN => n756);
   U1126 : XNOR2_X1 port map( A => n719, B => n756, ZN => n736);
   U1127 : NOR2_X1 port map( A1 => OP_A_10_port, A2 => OP_B_10_port, ZN => n757
                           );
   U1128 : OAI22_X1 port map( A1 => n757, A2 => n1367, B1 => n1371, B2 => n719,
                           ZN => n720);
   U1129 : AOI211_X1 port map( C1 => n1328, C2 => n721, A => n753, B => n720, 
                           ZN => n735);
   U1130 : AOI22_X1 port map( A1 => n1347, A2 => OP2(10), B1 => n1346, B2 => 
                           OP1(10), ZN => n722);
   U1131 : OAI21_X1 port map( B1 => n755, B2 => n1368, A => n722, ZN => n733);
   U1132 : OAI22_X1 port map( A1 => n824, A2 => n868, B1 => intadd_2_SUM_2_port
                           , B2 => n1283, ZN => n732);
   U1133 : NAND4_X1 port map( A1 => n726, A2 => n725, A3 => n724, A4 => n723, 
                           ZN => n939);
   U1134 : AOI222_X1 port map( A1 => n820, A2 => n855, B1 => n940, B2 => n853, 
                           C1 => n939, C2 => n894, ZN => n1211);
   U1135 : AOI22_X1 port map( A1 => n65, A2 => n1327, B1 => n894, B2 => n837, 
                           ZN => n1181);
   U1136 : OAI22_X1 port map( A1 => n1211, A2 => n885, B1 => n1181, B2 => n764,
                           ZN => n731);
   U1137 : OAI22_X1 port map( A1 => n729, A2 => n823, B1 => n728, B2 => n727, 
                           ZN => n730);
   U1138 : NOR4_X1 port map( A1 => n733, A2 => n732, A3 => n731, A4 => n730, ZN
                           => n734);
   U1139 : OAI211_X1 port map( C1 => n1397, C2 => n736, A => n735, B => n734, 
                           ZN => Y(10));
   U1140 : AOI22_X1 port map( A1 => n866, A2 => n874, B1 => n838, B2 => n863, 
                           ZN => n763);
   U1141 : OAI22_X1 port map( A1 => n1373, A2 => n742, B1 => n869, B2 => n765, 
                           ZN => n1250);
   U1142 : NAND4_X1 port map( A1 => n740, A2 => n739, A3 => n738, A4 => n737, 
                           ZN => n973);
   U1143 : INV_X1 port map( A => n973, ZN => n1111);
   U1144 : OAI222_X1 port map( A1 => n742, A2 => n963, B1 => n765, B2 => n1111,
                           C1 => n741, C2 => n966, ZN => n1242);
   U1145 : AOI22_X1 port map( A1 => n744, A2 => n1250, B1 => n743, B2 => n1242,
                           ZN => n762);
   U1146 : AOI22_X1 port map( A1 => OP1(11), A2 => n1329, B1 => n1366, B2 => 
                           n773, ZN => n746);
   U1147 : NAND2_X1 port map( A1 => n1347, A2 => OP2(11), ZN => n745);
   U1148 : OAI211_X1 port map( C1 => intadd_2_SUM_3_port, C2 => n1283, A => 
                           n746, B => n745, ZN => n752);
   U1149 : OAI22_X1 port map( A1 => n748, A2 => n823, B1 => n747, B2 => n1372, 
                           ZN => n751);
   U1150 : OAI22_X1 port map( A1 => n749, A2 => n1368, B1 => n1371, B2 => n754,
                           ZN => n750);
   U1151 : NOR4_X1 port map( A1 => n753, A2 => n752, A3 => n751, A4 => n750, ZN
                           => n761);
   U1152 : INV_X1 port map( A => n754, ZN => n759);
   U1153 : OAI21_X1 port map( B1 => n757, B2 => n756, A => n755, ZN => n774);
   U1154 : AOI21_X1 port map( B1 => n759, B2 => n774, A => n1397, ZN => n758);
   U1155 : OAI21_X1 port map( B1 => n759, B2 => n774, A => n758, ZN => n760);
   U1156 : NAND4_X1 port map( A1 => n763, A2 => n762, A3 => n761, A4 => n760, 
                           ZN => Y(11));
   U1157 : NOR2_X1 port map( A1 => n765, A2 => n764, ZN => n876);
   U1158 : NAND4_X1 port map( A1 => n769, A2 => n768, A3 => n767, A4 => n766, 
                           ZN => n1118);
   U1159 : AOI222_X1 port map( A1 => n1006, A2 => n65, B1 => OP_B_3_port, B2 =>
                           n770, C1 => n1118, C2 => n894, ZN => n1277);
   U1160 : OAI22_X1 port map( A1 => n1277, A2 => n885, B1 => n771, B2 => n1372,
                           ZN => n772);
   U1161 : AOI21_X1 port map( B1 => n876, B2 => n1264, A => n772, ZN => n790);
   U1162 : AOI22_X1 port map( A1 => OP_A_11_port, A2 => OP_B_11_port, B1 => 
                           n774, B2 => n773, ZN => n828);
   U1163 : NOR2_X1 port map( A1 => n828, A2 => n779, ZN => n775);
   U1164 : AOI211_X1 port map( C1 => n828, C2 => n779, A => n1397, B => n775, 
                           ZN => n788);
   U1165 : OAI22_X1 port map( A1 => intadd_2_SUM_4_port, A2 => n1283, B1 => 
                           n1138, B2 => n776, ZN => n787);
   U1166 : AOI22_X1 port map( A1 => n1329, A2 => OP1(12), B1 => n866, B2 => 
                           n777, ZN => n778);
   U1167 : OAI21_X1 port map( B1 => n779, B2 => n1371, A => n778, ZN => n786);
   U1168 : AOI22_X1 port map( A1 => n838, A2 => n781, B1 => n1366, B2 => n780, 
                           ZN => n783);
   U1169 : NOR2_X1 port map( A1 => n894, A2 => n1108, ZN => n861);
   U1170 : INV_X1 port map( A => n861, ZN => n782);
   U1171 : OAI211_X1 port map( C1 => n784, C2 => n823, A => n783, B => n782, ZN
                           => n785);
   U1172 : NOR4_X1 port map( A1 => n788, A2 => n787, A3 => n786, A4 => n785, ZN
                           => n789);
   U1173 : OAI211_X1 port map( C1 => n827, C2 => n1368, A => n790, B => n789, 
                           ZN => Y(12));
   U1174 : AOI22_X1 port map( A1 => n864, A2 => n792, B1 => n838, B2 => n791, 
                           ZN => n815);
   U1175 : AOI22_X1 port map( A1 => n866, A2 => n794, B1 => n1366, B2 => n793, 
                           ZN => n814);
   U1176 : OAI22_X1 port map( A1 => n795, A2 => n1372, B1 => n829, B2 => n1368,
                           ZN => n796);
   U1177 : AOI211_X1 port map( C1 => n876, C2 => n797, A => n861, B => n796, ZN
                           => n813);
   U1178 : INV_X1 port map( A => n798, ZN => n807);
   U1179 : AOI21_X1 port map( B1 => n828, B2 => n827, A => n830, ZN => n799);
   U1180 : XOR2_X1 port map( A => n807, B => n799, Z => n811);
   U1181 : OAI22_X1 port map( A1 => intadd_2_SUM_5_port, A2 => n1283, B1 => 
                           n1138, B2 => n800, ZN => n810);
   U1182 : NAND4_X1 port map( A1 => n804, A2 => n803, A3 => n802, A4 => n801, 
                           ZN => n1169);
   U1183 : AOI22_X1 port map( A1 => n855, A2 => n919, B1 => n853, B2 => n1037, 
                           ZN => n805);
   U1184 : OAI21_X1 port map( B1 => n920, B2 => n857, A => n805, ZN => n806);
   U1185 : AOI21_X1 port map( B1 => n894, B2 => n1169, A => n806, ZN => n1294);
   U1186 : AOI22_X1 port map( A1 => n807, A2 => n1343, B1 => n1346, B2 => 
                           OP1(13), ZN => n808);
   U1187 : OAI21_X1 port map( B1 => n1294, B2 => n885, A => n808, ZN => n809);
   U1188 : AOI211_X1 port map( C1 => n811, C2 => N279, A => n810, B => n809, ZN
                           => n812);
   U1189 : NAND4_X1 port map( A1 => n815, A2 => n814, A3 => n813, A4 => n812, 
                           ZN => Y(13));
   U1190 : NOR2_X1 port map( A1 => OP_A_14_port, A2 => OP_B_14_port, ZN => n872
                           );
   U1191 : NAND4_X1 port map( A1 => n819, A2 => n818, A3 => n817, A4 => n816, 
                           ZN => n1206);
   U1192 : INV_X1 port map( A => n820, ZN => n932);
   U1193 : AOI22_X1 port map( A1 => n855, A2 => n940, B1 => n65, B2 => n939, ZN
                           => n821);
   U1194 : OAI21_X1 port map( B1 => n932, B2 => n857, A => n821, ZN => n822);
   U1195 : AOI21_X1 port map( B1 => n894, B2 => n1206, A => n822, ZN => n1325);
   U1196 : OAI22_X1 port map( A1 => n824, A2 => n823, B1 => n1325, B2 => n885, 
                           ZN => n825);
   U1197 : AOI21_X1 port map( B1 => n866, B2 => n826, A => n825, ZN => n848);
   U1198 : INV_X1 port map( A => n835, ZN => n842);
   U1199 : NAND2_X1 port map( A1 => n829, A2 => n827, ZN => n834);
   U1200 : INV_X1 port map( A => n828, ZN => n833);
   U1201 : OAI21_X1 port map( B1 => n831, B2 => n830, A => n829, ZN => n832);
   U1202 : OAI21_X1 port map( B1 => n834, B2 => n833, A => n832, ZN => n871);
   U1203 : INV_X1 port map( A => n871, ZN => n836);
   U1204 : AOI221_X1 port map( B1 => n842, B2 => n836, C1 => n835, C2 => n871, 
                           A => n1397, ZN => n846);
   U1205 : AOI22_X1 port map( A1 => n1347, A2 => OP2(14), B1 => n1346, B2 => 
                           OP1(14), ZN => n840);
   U1206 : AOI22_X1 port map( A1 => n838, A2 => n837, B1 => n876, B2 => n1327, 
                           ZN => n839);
   U1207 : OAI211_X1 port map( C1 => intadd_2_SUM_6_port, C2 => n1283, A => 
                           n840, B => n839, ZN => n845);
   U1208 : AOI22_X1 port map( A1 => n842, A2 => n1343, B1 => n1328, B2 => n841,
                           ZN => n843);
   U1209 : OAI21_X1 port map( B1 => n870, B2 => n1368, A => n843, ZN => n844);
   U1210 : NOR4_X1 port map( A1 => n861, A2 => n846, A3 => n845, A4 => n844, ZN
                           => n847);
   U1211 : OAI211_X1 port map( C1 => n872, C2 => n1367, A => n848, B => n847, 
                           ZN => Y(14));
   U1212 : NAND4_X1 port map( A1 => n852, A2 => n851, A3 => n850, A4 => n849, 
                           ZN => n1228);
   U1213 : AOI22_X1 port map( A1 => n855, A2 => n854, B1 => n66, B2 => n973, ZN
                           => n856);
   U1214 : OAI21_X1 port map( B1 => n966, B2 => n857, A => n856, ZN => n858);
   U1215 : AOI21_X1 port map( B1 => n894, B2 => n1228, A => n858, ZN => n1363);
   U1216 : OAI22_X1 port map( A1 => intadd_2_SUM_7_port, A2 => n1283, B1 => 
                           n1138, B2 => n859, ZN => n860);
   U1217 : AOI211_X1 port map( C1 => n1329, C2 => OP1(15), A => n861, B => n860
                           , ZN => n884);
   U1218 : INV_X1 port map( A => n862, ZN => n901);
   U1219 : AOI22_X1 port map( A1 => n866, A2 => n865, B1 => n864, B2 => n863, 
                           ZN => n867);
   U1220 : OAI21_X1 port map( B1 => n869, B2 => n868, A => n867, ZN => n882);
   U1221 : OAI21_X1 port map( B1 => n872, B2 => n871, A => n870, ZN => n902);
   U1222 : XNOR2_X1 port map( A => n873, B => n902, ZN => n880);
   U1223 : AOI22_X1 port map( A1 => n1328, A2 => n874, B1 => n1343, B2 => n873,
                           ZN => n879);
   U1224 : INV_X1 port map( A => n1373, ZN => n875);
   U1225 : AOI22_X1 port map( A1 => n877, A2 => n1244, B1 => n876, B2 => n875, 
                           ZN => n878);
   U1226 : OAI211_X1 port map( C1 => n1397, C2 => n880, A => n879, B => n878, 
                           ZN => n881);
   U1227 : AOI211_X1 port map( C1 => n1366, C2 => n901, A => n882, B => n881, 
                           ZN => n883);
   U1228 : OAI211_X1 port map( C1 => n1363, C2 => n885, A => n884, B => n883, 
                           ZN => Y(15));
   U1229 : AOI22_X1 port map( A1 => n1347, A2 => OP2(16), B1 => n1346, B2 => 
                           OP1(16), ZN => n911);
   U1230 : OAI22_X1 port map( A1 => intadd_2_SUM_8_port, A2 => n1283, B1 => 
                           n949, B2 => n1368, ZN => n886);
   U1231 : NOR2_X1 port map( A1 => n1120, A2 => n886, ZN => n910);
   U1232 : NAND4_X1 port map( A1 => n890, A2 => n889, A3 => n888, A4 => n887, 
                           ZN => n1267);
   U1233 : INV_X1 port map( A => n1267, ZN => n893);
   U1234 : NOR2_X1 port map( A1 => n900, A2 => n891, ZN => n1229);
   U1235 : INV_X1 port map( A => n1229, ZN => n1110);
   U1236 : OAI22_X1 port map( A1 => n893, A2 => n1061, B1 => n892, B2 => n1110,
                           ZN => n897);
   U1237 : NOR2_X1 port map( A1 => n900, A2 => n1362, ZN => n1243);
   U1238 : NAND2_X1 port map( A1 => n894, A2 => n1243, ZN => n965);
   U1239 : OAI22_X1 port map( A1 => n952, A2 => n1367, B1 => n965, B2 => n895, 
                           ZN => n896);
   U1240 : AOI211_X1 port map( C1 => n1251, C2 => n898, A => n897, B => n896, 
                           ZN => n909);
   U1241 : NOR2_X1 port map( A1 => n900, A2 => n899, ZN => n1241);
   U1242 : AOI22_X1 port map( A1 => OP_A_15_port, A2 => OP_B_15_port, B1 => 
                           n902, B2 => n901, ZN => n950);
   U1243 : NOR2_X1 port map( A1 => n950, A2 => n904, ZN => n903);
   U1244 : AOI211_X1 port map( C1 => n950, C2 => n904, A => n1397, B => n903, 
                           ZN => n907);
   U1245 : NAND2_X1 port map( A1 => n1349, A2 => n1365, ZN => n1232);
   U1246 : OAI22_X1 port map( A1 => n905, A2 => n1232, B1 => n904, B2 => n1371,
                           ZN => n906);
   U1247 : AOI211_X1 port map( C1 => n1241, C2 => n1118, A => n907, B => n906, 
                           ZN => n908);
   U1248 : NAND4_X1 port map( A1 => n911, A2 => n910, A3 => n909, A4 => n908, 
                           ZN => Y(16));
   U1249 : NAND4_X1 port map( A1 => n915, A2 => n914, A3 => n913, A4 => n912, 
                           ZN => n1284);
   U1250 : AOI22_X1 port map( A1 => n918, A2 => n1343, B1 => n1227, B2 => n1284
                           , ZN => n930);
   U1251 : AOI22_X1 port map( A1 => n1347, A2 => OP2(17), B1 => n1346, B2 => 
                           OP1(17), ZN => n916);
   U1252 : OAI211_X1 port map( C1 => intadd_2_SUM_9_port, C2 => n1283, A => 
                           n916, B => n1108, ZN => n927);
   U1253 : AOI21_X1 port map( B1 => n950, B2 => n949, A => n952, ZN => n917);
   U1254 : XNOR2_X1 port map( A => n918, B => n917, ZN => n925);
   U1255 : AOI22_X1 port map( A1 => n1229, A2 => n919, B1 => n1241, B2 => n1169
                           , ZN => n924);
   U1256 : OAI22_X1 port map( A1 => n920, A2 => n965, B1 => n953, B2 => n1367, 
                           ZN => n921);
   U1257 : AOI21_X1 port map( B1 => n1251, B2 => n922, A => n921, ZN => n923);
   U1258 : OAI211_X1 port map( C1 => n1397, C2 => n925, A => n924, B => n923, 
                           ZN => n926);
   U1259 : AOI211_X1 port map( C1 => n928, C2 => n1244, A => n927, B => n926, 
                           ZN => n929);
   U1260 : OAI211_X1 port map( C1 => n931, C2 => n1232, A => n930, B => n929, 
                           ZN => Y(17));
   U1261 : OAI22_X1 port map( A1 => n932, A2 => n965, B1 => n982, B2 => n1367, 
                           ZN => n933);
   U1262 : AOI211_X1 port map( C1 => n1251, C2 => n934, A => n1120, B => n933, 
                           ZN => n961);
   U1263 : NAND4_X1 port map( A1 => n938, A2 => n937, A3 => n936, A4 => n935, 
                           ZN => n1315);
   U1264 : INV_X1 port map( A => n1315, ZN => n1209);
   U1265 : INV_X1 port map( A => n939, ZN => n1068);
   U1266 : OAI22_X1 port map( A1 => n1209, A2 => n1061, B1 => n1068, B2 => 
                           n1232, ZN => n947);
   U1267 : INV_X1 port map( A => n940, ZN => n945);
   U1268 : AOI222_X1 port map( A1 => n1413, A2 => C429_DATA4_18, B1 => 
                           OP_A_12_port, B2 => n63, C1 => OP_A_11_port, C2 => 
                           n1027, ZN => n978);
   U1269 : XOR2_X1 port map( A => n978, B => intadd_1_SUM_12_port, Z => n941);
   U1270 : XNOR2_X1 port map( A => intadd_2_n1, B => n941, ZN => n942);
   U1271 : AOI22_X1 port map( A1 => n986, A2 => n942, B1 => n1241, B2 => n1206,
                           ZN => n944);
   U1272 : AOI22_X1 port map( A1 => n1347, A2 => OP2(18), B1 => n1346, B2 => 
                           OP1(18), ZN => n943);
   U1273 : OAI211_X1 port map( C1 => n945, C2 => n1110, A => n944, B => n943, 
                           ZN => n946);
   U1274 : AOI211_X1 port map( C1 => n948, C2 => n1244, A => n947, B => n946, 
                           ZN => n960);
   U1275 : NAND2_X1 port map( A1 => n951, A2 => n949, ZN => n956);
   U1276 : INV_X1 port map( A => n950, ZN => n955);
   U1277 : OAI21_X1 port map( B1 => n953, B2 => n952, A => n951, ZN => n954);
   U1278 : OAI21_X1 port map( B1 => n956, B2 => n955, A => n954, ZN => n981);
   U1279 : XNOR2_X1 port map( A => n958, B => n981, ZN => n957);
   U1280 : AOI22_X1 port map( A1 => n958, A2 => n1343, B1 => N279, B2 => n957, 
                           ZN => n959);
   U1281 : NAND3_X1 port map( A1 => n961, A2 => n960, A3 => n959, ZN => Y(18));
   U1282 : AOI22_X1 port map( A1 => n1347, A2 => OP2(19), B1 => n1346, B2 => 
                           OP1(19), ZN => n962);
   U1283 : OAI21_X1 port map( B1 => n963, B2 => n1110, A => n962, ZN => n968);
   U1284 : INV_X1 port map( A => n1251, ZN => n1180);
   U1285 : OAI22_X1 port map( A1 => n966, A2 => n965, B1 => n964, B2 => n1180, 
                           ZN => n967);
   U1286 : AOI211_X1 port map( C1 => n1366, C2 => n991, A => n968, B => n967, 
                           ZN => n990);
   U1287 : NAND4_X1 port map( A1 => n972, A2 => n971, A3 => n970, A4 => n969, 
                           ZN => n1350);
   U1288 : INV_X1 port map( A => n1232, ZN => n1121);
   U1289 : AOI22_X1 port map( A1 => n1227, A2 => n1350, B1 => n1121, B2 => n973
                           , ZN => n989);
   U1290 : OAI22_X1 port map( A1 => n975, A2 => n1368, B1 => n1371, B2 => n974,
                           ZN => n976);
   U1291 : AOI211_X1 port map( C1 => n1241, C2 => n1228, A => n1120, B => n976,
                           ZN => n988);
   U1292 : AND2_X1 port map( A1 => intadd_1_SUM_12_port, A2 => intadd_2_n1, ZN 
                           => n977);
   U1293 : OAI22_X1 port map( A1 => n978, A2 => n977, B1 => 
                           intadd_1_SUM_12_port, B2 => intadd_2_n1, ZN => n994)
                           ;
   U1294 : AOI222_X1 port map( A1 => n1413, A2 => C429_DATA4_19, B1 => 
                           OP_A_12_port, B2 => n1027, C1 => n63, C2 => 
                           OP_A_13_port, ZN => n997);
   U1295 : XNOR2_X1 port map( A => intadd_1_SUM_13_port, B => n997, ZN => n979)
                           ;
   U1296 : XNOR2_X1 port map( A => n994, B => n979, ZN => n985);
   U1297 : OAI21_X1 port map( B1 => n982, B2 => n981, A => n980, ZN => n992);
   U1298 : XOR2_X1 port map( A => n983, B => n992, Z => n984);
   U1299 : AOI22_X1 port map( A1 => n986, A2 => n985, B1 => n984, B2 => N279, 
                           ZN => n987);
   U1300 : NAND4_X1 port map( A1 => n990, A2 => n989, A3 => n988, A4 => n987, 
                           ZN => Y(19));
   U1301 : AOI22_X1 port map( A1 => n1241, A2 => n1267, B1 => n1121, B2 => 
                           n1118, ZN => n1017);
   U1302 : AOI22_X1 port map( A1 => OP_A_19_port, A2 => OP_B_19_port, B1 => 
                           n992, B2 => n991, ZN => n1047);
   U1303 : NOR2_X1 port map( A1 => n1047, A2 => n1018, ZN => n993);
   U1304 : AOI211_X1 port map( C1 => n1047, C2 => n1018, A => n1397, B => n993,
                           ZN => n1015);
   U1305 : INV_X1 port map( A => n994, ZN => n998);
   U1306 : INV_X1 port map( A => intadd_1_SUM_13_port, ZN => n995);
   U1307 : NAND2_X1 port map( A1 => n995, A2 => n994, ZN => n996);
   U1308 : AOI22_X1 port map( A1 => intadd_1_SUM_13_port, A2 => n998, B1 => 
                           n997, B2 => n996, ZN => n1026);
   U1309 : AOI222_X1 port map( A1 => n1413, A2 => C429_DATA4_20, B1 => n63, B2 
                           => OP_A_14_port, C1 => n1027, C2 => OP_A_13_port, ZN
                           => n1022);
   U1310 : INV_X1 port map( A => intadd_1_SUM_14_port, ZN => n1025);
   U1311 : XNOR2_X1 port map( A => n1022, B => n1025, ZN => n999);
   U1312 : XNOR2_X1 port map( A => n1026, B => n999, ZN => n1000);
   U1313 : NOR2_X1 port map( A1 => n1000, A2 => n1283, ZN => n1014);
   U1314 : AOI22_X1 port map( A1 => n1347, A2 => OP2(20), B1 => n1346, B2 => 
                           OP1(20), ZN => n1001);
   U1315 : OAI211_X1 port map( C1 => n1368, C2 => n1046, A => n1001, B => n1108
                           , ZN => n1013);
   U1316 : INV_X1 port map( A => n1243, ZN => n1210);
   U1317 : NAND4_X1 port map( A1 => n1005, A2 => n1004, A3 => n1003, A4 => 
                           n1002, ZN => n1268);
   U1318 : AOI22_X1 port map( A1 => n1227, A2 => n1268, B1 => n1229, B2 => 
                           n1006, ZN => n1010);
   U1319 : AOI22_X1 port map( A1 => n1251, A2 => n1008, B1 => n1366, B2 => 
                           n1007, ZN => n1009);
   U1320 : OAI211_X1 port map( C1 => n1210, C2 => n1011, A => n1010, B => n1009
                           , ZN => n1012);
   U1321 : NOR4_X1 port map( A1 => n1015, A2 => n1014, A3 => n1013, A4 => n1012
                           , ZN => n1016);
   U1322 : OAI211_X1 port map( C1 => n1018, C2 => n1371, A => n1017, B => n1016
                           , ZN => Y(20));
   U1323 : AOI21_X1 port map( B1 => n1047, B2 => n1046, A => n1049, ZN => n1019
                           );
   U1324 : XNOR2_X1 port map( A => n1020, B => n1019, ZN => n1045);
   U1325 : AOI22_X1 port map( A1 => n1021, A2 => n1244, B1 => n1020, B2 => 
                           n1343, ZN => n1044);
   U1326 : INV_X1 port map( A => n1026, ZN => n1023);
   U1327 : OAI21_X1 port map( B1 => intadd_1_SUM_14_port, B2 => n1023, A => 
                           n1022, ZN => n1024);
   U1328 : OAI21_X1 port map( B1 => n1026, B2 => n1025, A => n1024, ZN => n1076
                           );
   U1329 : INV_X1 port map( A => n1076, ZN => n1073);
   U1330 : AOI222_X1 port map( A1 => OP_A_15_port, A2 => n63, B1 => n1413, B2 
                           => C429_DATA4_21, C1 => n1027, C2 => OP_A_14_port, 
                           ZN => n1075);
   U1331 : INV_X1 port map( A => intadd_1_SUM_15_port, ZN => n1072);
   U1332 : XNOR2_X1 port map( A => n1075, B => n1072, ZN => n1028);
   U1333 : XNOR2_X1 port map( A => n1073, B => n1028, ZN => n1032);
   U1334 : AOI22_X1 port map( A1 => n1347, A2 => OP2(21), B1 => n1329, B2 => 
                           OP1(21), ZN => n1031);
   U1335 : AOI22_X1 port map( A1 => n1243, A2 => n1029, B1 => n1241, B2 => 
                           n1284, ZN => n1030);
   U1336 : OAI211_X1 port map( C1 => n1032, C2 => n1283, A => n1031, B => n1030
                           , ZN => n1042);
   U1337 : NAND4_X1 port map( A1 => n1036, A2 => n1035, A3 => n1034, A4 => 
                           n1033, ZN => n1285);
   U1338 : AOI22_X1 port map( A1 => n1227, A2 => n1285, B1 => n1229, B2 => 
                           n1037, ZN => n1040);
   U1339 : AOI21_X1 port map( B1 => n1251, B2 => n1038, A => n1120, ZN => n1039
                           );
   U1340 : OAI211_X1 port map( C1 => n1050, C2 => n1367, A => n1040, B => n1039
                           , ZN => n1041);
   U1341 : AOI211_X1 port map( C1 => n1121, C2 => n1169, A => n1042, B => n1041
                           , ZN => n1043);
   U1342 : OAI211_X1 port map( C1 => n1397, C2 => n1045, A => n1044, B => n1043
                           , ZN => Y(21));
   U1343 : INV_X1 port map( A => n1124, ZN => n1055);
   U1344 : NAND2_X1 port map( A1 => n1048, A2 => n1046, ZN => n1053);
   U1345 : INV_X1 port map( A => n1047, ZN => n1052);
   U1346 : OAI21_X1 port map( B1 => n1050, B2 => n1049, A => n1048, ZN => n1051
                           );
   U1347 : OAI21_X1 port map( B1 => n1053, B2 => n1052, A => n1051, ZN => n1125
                           );
   U1348 : INV_X1 port map( A => n1125, ZN => n1054);
   U1349 : AOI221_X1 port map( B1 => n1055, B2 => n1054, C1 => n1124, C2 => 
                           n1125, A => n1397, ZN => n1071);
   U1350 : NOR2_X1 port map( A1 => OP_A_22_port, A2 => OP_B_22_port, ZN => 
                           n1103);
   U1351 : OAI22_X1 port map( A1 => n1103, A2 => n1367, B1 => n1123, B2 => 
                           n1368, ZN => n1070);
   U1352 : AOI22_X1 port map( A1 => n1347, A2 => OP2(22), B1 => n1329, B2 => 
                           OP1(22), ZN => n1067);
   U1353 : NAND4_X1 port map( A1 => n1059, A2 => n1058, A3 => n1057, A4 => 
                           n1056, ZN => n1316);
   U1354 : INV_X1 port map( A => n1316, ZN => n1183);
   U1355 : INV_X1 port map( A => n1206, ZN => n1060);
   U1356 : OAI22_X1 port map( A1 => n1183, A2 => n1061, B1 => n1060, B2 => 
                           n1232, ZN => n1064);
   U1357 : INV_X1 port map( A => n1241, ZN => n1182);
   U1358 : OAI22_X1 port map( A1 => n1209, A2 => n1182, B1 => n1062, B2 => 
                           n1210, ZN => n1063);
   U1359 : AOI211_X1 port map( C1 => n1251, C2 => n1065, A => n1064, B => n1063
                           , ZN => n1066);
   U1360 : OAI211_X1 port map( C1 => n1068, C2 => n1110, A => n1067, B => n1066
                           , ZN => n1069);
   U1361 : NOR4_X1 port map( A1 => n1120, A2 => n1071, A3 => n1070, A4 => n1069
                           , ZN => n1087);
   U1362 : NAND2_X1 port map( A1 => n1073, A2 => n1072, ZN => n1074);
   U1363 : AOI22_X1 port map( A1 => intadd_1_SUM_15_port, A2 => n1076, B1 => 
                           n1075, B2 => n1074, ZN => n1090);
   U1364 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n1078, A => n1077, ZN 
                           => n1079);
   U1365 : INV_X1 port map( A => n1079, ZN => n1091);
   U1366 : XNOR2_X1 port map( A => DP_OP_446J3_125_4819_n12, B => n1091, ZN => 
                           n1082);
   U1367 : AOI21_X1 port map( B1 => n1413, B2 => n1082, A => n1379, ZN => n1083
                           );
   U1368 : INV_X1 port map( A => n1083, ZN => n1089);
   U1369 : XNOR2_X1 port map( A => n1090, B => n1089, ZN => n1085);
   U1370 : AOI21_X1 port map( B1 => intadd_1_SUM_16_port, B2 => n1085, A => 
                           n1283, ZN => n1084);
   U1371 : OAI21_X1 port map( B1 => intadd_1_SUM_16_port, B2 => n1085, A => 
                           n1084, ZN => n1086);
   U1372 : OAI211_X1 port map( C1 => n1371, C2 => n1124, A => n1087, B => n1086
                           , ZN => Y(22));
   U1373 : INV_X1 port map( A => intadd_1_SUM_16_port, ZN => n1088);
   U1374 : FA_X1 port map( A => n1090, B => n1089, CI => n1088, CO => n1092, S 
                           => n_1170);
   U1375 : NOR3_X1 port map( A1 => n1092, A2 => n59, A3 => n1379, ZN => n1142);
   U1376 : INV_X1 port map( A => n1142, ZN => n1093);
   U1377 : OAI21_X1 port map( B1 => n1379, B2 => n59, A => n1092, ZN => n1143);
   U1378 : NAND2_X1 port map( A1 => n1093, A2 => n1143, ZN => n1094);
   U1379 : XNOR2_X1 port map( A => intadd_1_SUM_17_port, B => n1094, ZN => 
                           n1117);
   U1380 : NAND4_X1 port map( A1 => n1098, A2 => n1097, A3 => n1096, A4 => 
                           n1095, ZN => n1348);
   U1381 : AOI22_X1 port map( A1 => n1227, A2 => n1348, B1 => n1121, B2 => 
                           n1228, ZN => n1101);
   U1382 : AOI22_X1 port map( A1 => n1243, A2 => n1099, B1 => n1241, B2 => 
                           n1350, ZN => n1100);
   U1383 : OAI211_X1 port map( C1 => n1122, C2 => n1368, A => n1101, B => n1100
                           , ZN => n1102);
   U1384 : AOI21_X1 port map( B1 => n1343, B2 => n1105, A => n1102, ZN => n1116
                           );
   U1385 : OAI21_X1 port map( B1 => n1103, B2 => n1125, A => n1123, ZN => n1104
                           );
   U1386 : XOR2_X1 port map( A => n1105, B => n1104, Z => n1114);
   U1387 : OAI22_X1 port map( A1 => n1107, A2 => n1367, B1 => n1106, B2 => 
                           n1180, ZN => n1113);
   U1388 : AOI22_X1 port map( A1 => n1347, A2 => OP2(23), B1 => n1329, B2 => 
                           OP1(23), ZN => n1109);
   U1389 : OAI211_X1 port map( C1 => n1111, C2 => n1110, A => n1109, B => n1108
                           , ZN => n1112);
   U1390 : AOI211_X1 port map( C1 => n1114, C2 => N279, A => n1113, B => n1112,
                           ZN => n1115);
   U1391 : OAI211_X1 port map( C1 => n1283, C2 => n1117, A => n1116, B => n1115
                           , ZN => Y(23));
   U1392 : AOI22_X1 port map( A1 => n1241, A2 => n1268, B1 => n1229, B2 => 
                           n1118, ZN => n1151);
   U1393 : OAI22_X1 port map( A1 => n1192, A2 => n1368, B1 => n1128, B2 => 
                           n1371, ZN => n1119);
   U1394 : AOI211_X1 port map( C1 => n1121, C2 => n1267, A => n1120, B => n1119
                           , ZN => n1150);
   U1395 : OAI211_X1 port map( C1 => n1125, C2 => n1124, A => n1123, B => n1122
                           , ZN => n1126);
   U1396 : OAI21_X1 port map( B1 => OP_A_23_port, B2 => OP_B_23_port, A => 
                           n1126, ZN => n1191);
   U1397 : NOR2_X1 port map( A1 => n1191, A2 => n1128, ZN => n1127);
   U1398 : AOI211_X1 port map( C1 => n1191, C2 => n1128, A => n1397, B => n1127
                           , ZN => n1140);
   U1399 : NAND4_X1 port map( A1 => n1132, A2 => n1131, A3 => n1130, A4 => 
                           n1129, ZN => n1273);
   U1400 : AOI22_X1 port map( A1 => n1329, A2 => OP1(24), B1 => n1227, B2 => 
                           n1273, ZN => n1136);
   U1401 : AOI22_X1 port map( A1 => n1251, A2 => n1134, B1 => n1243, B2 => 
                           n1133, ZN => n1135);
   U1402 : OAI211_X1 port map( C1 => n1138, C2 => n1137, A => n1136, B => n1135
                           , ZN => n1139);
   U1403 : AOI211_X1 port map( C1 => n1366, C2 => n1141, A => n1140, B => n1139
                           , ZN => n1149);
   U1404 : AOI21_X1 port map( B1 => intadd_1_SUM_17_port, B2 => n1143, A => 
                           n1142, ZN => n1144);
   U1405 : NOR3_X1 port map( A1 => n1144, A2 => n59, A3 => n1379, ZN => n1152);
   U1406 : INV_X1 port map( A => n1152, ZN => n1145);
   U1407 : OAI21_X1 port map( B1 => n1379, B2 => n59, A => n1144, ZN => n1153);
   U1408 : NAND2_X1 port map( A1 => n1145, A2 => n1153, ZN => n1147);
   U1409 : AOI21_X1 port map( B1 => intadd_1_SUM_18_port, B2 => n1147, A => 
                           n1283, ZN => n1146);
   U1410 : OAI21_X1 port map( B1 => intadd_1_SUM_18_port, B2 => n1147, A => 
                           n1146, ZN => n1148);
   U1411 : NAND4_X1 port map( A1 => n1151, A2 => n1150, A3 => n1149, A4 => 
                           n1148, ZN => Y(24));
   U1412 : AOI21_X1 port map( B1 => intadd_1_SUM_18_port, B2 => n1153, A => 
                           n1152, ZN => n1154);
   U1413 : NOR3_X1 port map( A1 => n1154, A2 => n59, A3 => n1379, ZN => n1185);
   U1414 : INV_X1 port map( A => n1185, ZN => n1155);
   U1415 : OAI21_X1 port map( B1 => n1379, B2 => n59, A => n1154, ZN => n1186);
   U1416 : NAND2_X1 port map( A1 => n1155, A2 => n1186, ZN => n1156);
   U1417 : XNOR2_X1 port map( A => intadd_1_SUM_19_port, B => n1156, ZN => 
                           n1179);
   U1418 : AOI211_X1 port map( C1 => n1159, C2 => n1362, A => n1158, B => n1157
                           , ZN => n1235);
   U1419 : AOI22_X1 port map( A1 => n1243, A2 => n1160, B1 => n1241, B2 => 
                           n1285, ZN => n1161);
   U1420 : OAI21_X1 port map( B1 => n1193, B2 => n1368, A => n1161, ZN => n1162
                           );
   U1421 : AOI211_X1 port map( C1 => n1164, C2 => n1343, A => n1235, B => n1162
                           , ZN => n1178);
   U1422 : AOI21_X1 port map( B1 => n1191, B2 => n1192, A => n1194, ZN => n1163
                           );
   U1423 : XOR2_X1 port map( A => n1164, B => n1163, Z => n1176);
   U1424 : INV_X1 port map( A => n1284, ZN => n1172);
   U1425 : NAND4_X1 port map( A1 => n1168, A2 => n1167, A3 => n1166, A4 => 
                           n1165, ZN => n1290);
   U1426 : AOI22_X1 port map( A1 => n1229, A2 => n1169, B1 => n1227, B2 => 
                           n1290, ZN => n1171);
   U1427 : AOI22_X1 port map( A1 => n1347, A2 => OP2(25), B1 => n1329, B2 => 
                           OP1(25), ZN => n1170);
   U1428 : OAI211_X1 port map( C1 => n1172, C2 => n1232, A => n1171, B => n1170
                           , ZN => n1175);
   U1429 : OAI22_X1 port map( A1 => n1195, A2 => n1367, B1 => n1173, B2 => 
                           n1180, ZN => n1174);
   U1430 : AOI211_X1 port map( C1 => n1176, C2 => N279, A => n1175, B => n1174,
                           ZN => n1177);
   U1431 : OAI211_X1 port map( C1 => n1283, C2 => n1179, A => n1178, B => n1177
                           , ZN => Y(25));
   U1432 : INV_X1 port map( A => n1199, ZN => n1201);
   U1433 : OAI22_X1 port map( A1 => n1183, A2 => n1182, B1 => n1181, B2 => 
                           n1180, ZN => n1184);
   U1434 : AOI211_X1 port map( C1 => n1201, C2 => n1343, A => n1235, B => n1184
                           , ZN => n1217);
   U1435 : AOI21_X1 port map( B1 => intadd_1_SUM_19_port, B2 => n1186, A => 
                           n1185, ZN => n1187);
   U1436 : NOR3_X1 port map( A1 => n1187, A2 => n59, A3 => n1379, ZN => n1218);
   U1437 : INV_X1 port map( A => n1218, ZN => n1188);
   U1438 : OAI21_X1 port map( B1 => n1379, B2 => n59, A => n1187, ZN => n1219);
   U1439 : NAND2_X1 port map( A1 => n1188, A2 => n1219, ZN => n1190);
   U1440 : NOR2_X1 port map( A1 => intadd_1_SUM_20_port, A2 => n1190, ZN => 
                           n1189);
   U1441 : AOI211_X1 port map( C1 => intadd_1_SUM_20_port, C2 => n1190, A => 
                           n1283, B => n1189, ZN => n1215);
   U1442 : INV_X1 port map( A => n1191, ZN => n1198);
   U1443 : NAND2_X1 port map( A1 => n1193, A2 => n1192, ZN => n1197);
   U1444 : OAI21_X1 port map( B1 => n1195, B2 => n1194, A => n1193, ZN => n1196
                           );
   U1445 : OAI21_X1 port map( B1 => n1198, B2 => n1197, A => n1196, ZN => n1237
                           );
   U1446 : INV_X1 port map( A => n1237, ZN => n1200);
   U1447 : AOI221_X1 port map( B1 => n1201, B2 => n1200, C1 => n1199, C2 => 
                           n1237, A => n1397, ZN => n1214);
   U1448 : NAND4_X1 port map( A1 => n1205, A2 => n1204, A3 => n1203, A4 => 
                           n1202, ZN => n1321);
   U1449 : AOI22_X1 port map( A1 => n1229, A2 => n1206, B1 => n1227, B2 => 
                           n1321, ZN => n1208);
   U1450 : AOI22_X1 port map( A1 => n1347, A2 => OP2(26), B1 => n1329, B2 => 
                           OP1(26), ZN => n1207);
   U1451 : OAI211_X1 port map( C1 => n1209, C2 => n1232, A => n1208, B => n1207
                           , ZN => n1213);
   U1452 : NOR2_X1 port map( A1 => OP_A_26_port, A2 => OP_B_26_port, ZN => 
                           n1238);
   U1453 : OAI22_X1 port map( A1 => n1238, A2 => n1367, B1 => n1211, B2 => 
                           n1210, ZN => n1212);
   U1454 : NOR4_X1 port map( A1 => n1215, A2 => n1214, A3 => n1213, A4 => n1212
                           , ZN => n1216);
   U1455 : OAI211_X1 port map( C1 => n1236, C2 => n1368, A => n1217, B => n1216
                           , ZN => Y(26));
   U1456 : AOI21_X1 port map( B1 => intadd_1_SUM_20_port, B2 => n1219, A => 
                           n1218, ZN => n1220);
   U1457 : NOR3_X1 port map( A1 => n1220, A2 => n59, A3 => n1379, ZN => n1255);
   U1458 : INV_X1 port map( A => n1255, ZN => n1221);
   U1459 : OAI21_X1 port map( B1 => n1379, B2 => n59, A => n1220, ZN => n1256);
   U1460 : NAND2_X1 port map( A1 => n1221, A2 => n1256, ZN => n1222);
   U1461 : XNOR2_X1 port map( A => intadd_1_SUM_21_port, B => n1222, ZN => 
                           n1254);
   U1462 : INV_X1 port map( A => n1350, ZN => n1233);
   U1463 : NAND4_X1 port map( A1 => n1226, A2 => n1225, A3 => n1224, A4 => 
                           n1223, ZN => n1356);
   U1464 : AOI22_X1 port map( A1 => n1229, A2 => n1228, B1 => n1227, B2 => 
                           n1356, ZN => n1231);
   U1465 : AOI22_X1 port map( A1 => n1347, A2 => OP2(27), B1 => n1329, B2 => 
                           OP1(27), ZN => n1230);
   U1466 : OAI211_X1 port map( C1 => n1233, C2 => n1232, A => n1231, B => n1230
                           , ZN => n1234);
   U1467 : AOI211_X1 port map( C1 => n1343, C2 => n1240, A => n1235, B => n1234
                           , ZN => n1253);
   U1468 : OAI21_X1 port map( B1 => n1238, B2 => n1237, A => n1236, ZN => n1265
                           );
   U1469 : OAI21_X1 port map( B1 => n1240, B2 => n1265, A => N279, ZN => n1239)
                           ;
   U1470 : AOI21_X1 port map( B1 => n1240, B2 => n1265, A => n1239, ZN => n1249
                           );
   U1471 : AOI22_X1 port map( A1 => n1243, A2 => n1242, B1 => n1241, B2 => 
                           n1348, ZN => n1246);
   U1472 : OAI221_X1 port map( B1 => n1366, B2 => n1244, C1 => n1366, C2 => 
                           OP_A_27_port, A => OP_B_27_port, ZN => n1245);
   U1473 : OAI211_X1 port map( C1 => n1367, C2 => n1247, A => n1246, B => n1245
                           , ZN => n1248);
   U1474 : AOI211_X1 port map( C1 => n1251, C2 => n1250, A => n1249, B => n1248
                           , ZN => n1252);
   U1475 : OAI211_X1 port map( C1 => n1283, C2 => n1254, A => n1253, B => n1252
                           , ZN => Y(27));
   U1476 : AOI21_X1 port map( B1 => intadd_1_SUM_21_port, B2 => n1256, A => 
                           n1255, ZN => n1257);
   U1477 : NOR3_X1 port map( A1 => n1257, A2 => n59, A3 => n1379, ZN => n1302);
   U1478 : INV_X1 port map( A => n1302, ZN => n1258);
   U1479 : OAI21_X1 port map( B1 => n1379, B2 => n59, A => n1257, ZN => n1303);
   U1480 : NAND2_X1 port map( A1 => n1258, A2 => n1303, ZN => n1259);
   U1481 : XNOR2_X1 port map( A => intadd_1_SUM_22_port, B => n1259, ZN => 
                           n1282);
   U1482 : AOI22_X1 port map( A1 => n1347, A2 => OP2(28), B1 => n1329, B2 => 
                           OP1(28), ZN => n1261);
   U1483 : NAND3_X1 port map( A1 => OP_SHIFT, A2 => N284, A3 => n1260, ZN => 
                           n1401);
   U1484 : OAI211_X1 port map( C1 => n1298, C2 => n1367, A => n1261, B => n1401
                           , ZN => n1263);
   U1485 : OAI22_X1 port map( A1 => n1300, A2 => n1368, B1 => n1371, B2 => 
                           n1266, ZN => n1262);
   U1486 : AOI211_X1 port map( C1 => n1328, C2 => n1264, A => n1263, B => n1262
                           , ZN => n1281);
   U1487 : AOI222_X1 port map( A1 => OP_A_27_port, A2 => OP_B_27_port, B1 => 
                           OP_A_27_port, B2 => n1265, C1 => OP_B_27_port, C2 =>
                           n1265, ZN => n1299);
   U1488 : XOR2_X1 port map( A => n1266, B => n1299, Z => n1279);
   U1489 : AOI22_X1 port map( A1 => n1349, A2 => n1268, B1 => n1351, B2 => 
                           n1267, ZN => n1276);
   U1490 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n57, ZN => n1272);
   U1491 : NAND4_X1 port map( A1 => n1272, A2 => n1271, A3 => n1270, A4 => 
                           n1269, ZN => n1274);
   U1492 : AOI22_X1 port map( A1 => n1359, A2 => n1274, B1 => n1357, B2 => 
                           n1273, ZN => n1275);
   U1493 : OAI211_X1 port map( C1 => n1277, C2 => n1362, A => n1276, B => n1275
                           , ZN => n1278);
   U1494 : AOI22_X1 port map( A1 => n1279, A2 => N279, B1 => n1365, B2 => n1278
                           , ZN => n1280);
   U1495 : OAI211_X1 port map( C1 => n1283, C2 => n1282, A => n1281, B => n1280
                           , ZN => Y(28));
   U1496 : AOI22_X1 port map( A1 => n1347, A2 => OP2(29), B1 => n1329, B2 => 
                           OP1(29), ZN => n1314);
   U1497 : AOI22_X1 port map( A1 => n1349, A2 => n1285, B1 => n1351, B2 => 
                           n1284, ZN => n1293);
   U1498 : NAND4_X1 port map( A1 => n1289, A2 => n1288, A3 => n1287, A4 => 
                           n1286, ZN => n1291);
   U1499 : AOI22_X1 port map( A1 => n1359, A2 => n1291, B1 => n1357, B2 => 
                           n1290, ZN => n1292);
   U1500 : OAI211_X1 port map( C1 => n1294, C2 => n1362, A => n1293, B => n1292
                           , ZN => n1295);
   U1501 : AOI22_X1 port map( A1 => OP_A_29_port, A2 => n1366, B1 => n1365, B2 
                           => n1295, ZN => n1313);
   U1502 : OAI21_X1 port map( B1 => n1296, B2 => n1368, A => n1367, ZN => n1311
                           );
   U1503 : OAI22_X1 port map( A1 => n1301, A2 => n1371, B1 => n1297, B2 => 
                           n1372, ZN => n1310);
   U1504 : AOI21_X1 port map( B1 => n1300, B2 => n1299, A => n1298, ZN => n1331
                           );
   U1505 : XOR2_X1 port map( A => n1331, B => n1301, Z => n1308);
   U1506 : AOI21_X1 port map( B1 => intadd_1_SUM_22_port, B2 => n1303, A => 
                           n1302, ZN => n1304);
   U1507 : NOR3_X1 port map( A1 => n1304, A2 => n59, A3 => n1379, ZN => n1333);
   U1508 : INV_X1 port map( A => n1333, ZN => n1305);
   U1509 : OAI21_X1 port map( B1 => n1379, B2 => n59, A => n1304, ZN => n1334);
   U1510 : NAND2_X1 port map( A1 => n1305, A2 => n1334, ZN => n1306);
   U1511 : XNOR2_X1 port map( A => intadd_1_SUM_23_port, B => n1306, ZN => 
                           n1307);
   U1512 : OAI22_X1 port map( A1 => n1397, A2 => n1308, B1 => n1395, B2 => 
                           n1307, ZN => n1309);
   U1513 : AOI211_X1 port map( C1 => OP_B_29_port, C2 => n1311, A => n1310, B 
                           => n1309, ZN => n1312);
   U1514 : NAND4_X1 port map( A1 => n1314, A2 => n1313, A3 => n1312, A4 => 
                           n1401, ZN => Y(29));
   U1515 : AOI22_X1 port map( A1 => n1349, A2 => n1316, B1 => n1351, B2 => 
                           n1315, ZN => n1324);
   U1516 : NAND2_X1 port map( A1 => OP_A_30_port, A2 => n57, ZN => n1320);
   U1517 : NAND4_X1 port map( A1 => n1320, A2 => n1319, A3 => n1318, A4 => 
                           n1317, ZN => n1322);
   U1518 : AOI22_X1 port map( A1 => n1359, A2 => n1322, B1 => n1357, B2 => 
                           n1321, ZN => n1323);
   U1519 : OAI211_X1 port map( C1 => n1325, C2 => n1362, A => n1324, B => n1323
                           , ZN => n1326);
   U1520 : AOI22_X1 port map( A1 => n1328, A2 => n1327, B1 => n1365, B2 => 
                           n1326, ZN => n1345);
   U1521 : AOI22_X1 port map( A1 => n1347, A2 => OP2(30), B1 => n1329, B2 => 
                           OP1(30), ZN => n1330);
   U1522 : OAI211_X1 port map( C1 => n1374, C2 => n1367, A => n1330, B => n1401
                           , ZN => n1341);
   U1523 : AOI222_X1 port map( A1 => OP_B_29_port, A2 => OP_A_29_port, B1 => 
                           OP_B_29_port, B2 => n1331, C1 => OP_A_29_port, C2 =>
                           n1331, ZN => n1375);
   U1524 : XNOR2_X1 port map( A => n1375, B => n1332, ZN => n1339);
   U1525 : AOI21_X1 port map( B1 => intadd_1_SUM_23_port, B2 => n1334, A => 
                           n1333, ZN => n1335);
   U1526 : NOR3_X1 port map( A1 => n1335, A2 => n59, A3 => n1379, ZN => n1385);
   U1527 : INV_X1 port map( A => n1385, ZN => n1336);
   U1528 : OAI21_X1 port map( B1 => n1379, B2 => n59, A => n1335, ZN => n1386);
   U1529 : NAND2_X1 port map( A1 => n1336, A2 => n1386, ZN => n1337);
   U1530 : XNOR2_X1 port map( A => intadd_1_SUM_24_port, B => n1337, ZN => 
                           n1338);
   U1531 : OAI22_X1 port map( A1 => n1397, A2 => n1339, B1 => n1395, B2 => 
                           n1338, ZN => n1340);
   U1532 : AOI211_X1 port map( C1 => n1343, C2 => n1342, A => n1341, B => n1340
                           , ZN => n1344);
   U1533 : OAI211_X1 port map( C1 => n1376, C2 => n1368, A => n1345, B => n1344
                           , ZN => Y(30));
   U1534 : AOI22_X1 port map( A1 => n1347, A2 => OP2(31), B1 => OP1(31), B2 => 
                           n1346, ZN => n1404);
   U1535 : AOI22_X1 port map( A1 => n1351, A2 => n1350, B1 => n1349, B2 => 
                           n1348, ZN => n1361);
   U1536 : NAND2_X1 port map( A1 => OP_A_31_port, A2 => n57, ZN => n1355);
   U1537 : NAND4_X1 port map( A1 => n1355, A2 => n1354, A3 => n1353, A4 => 
                           n1352, ZN => n1358);
   U1538 : AOI22_X1 port map( A1 => n1359, A2 => n1358, B1 => n1357, B2 => 
                           n1356, ZN => n1360);
   U1539 : OAI211_X1 port map( C1 => n1363, C2 => n1362, A => n1361, B => n1360
                           , ZN => n1364);
   U1540 : AOI22_X1 port map( A1 => OP_A_31_port, A2 => n1366, B1 => n1365, B2 
                           => n1364, ZN => n1403);
   U1541 : OAI21_X1 port map( B1 => n1369, B2 => n1368, A => n1367, ZN => n1400
                           );
   U1542 : INV_X1 port map( A => n1370, ZN => n1377);
   U1543 : OAI22_X1 port map( A1 => n1373, A2 => n1372, B1 => n1377, B2 => 
                           n1371, ZN => n1399);
   U1544 : AOI21_X1 port map( B1 => n1376, B2 => n1375, A => n1374, ZN => n1378
                           );
   U1545 : XOR2_X1 port map( A => n1378, B => n1377, Z => n1396);
   U1546 : NOR2_X1 port map( A1 => n59, A2 => n1379, ZN => n1384);
   U1547 : INV_X1 port map( A => n1380, ZN => n1381);
   U1548 : AOI21_X1 port map( B1 => n1382, B2 => n1381, A => n1384, ZN => n1383
                           );
   U1549 : AOI21_X1 port map( B1 => n1384, B2 => intadd_1_B_18_port, A => n1383
                           , ZN => n1388);
   U1550 : AOI21_X1 port map( B1 => intadd_1_SUM_24_port, B2 => n1386, A => 
                           n1385, ZN => n1387);
   U1551 : XOR2_X1 port map( A => n1388, B => n1387, Z => n1389);
   U1552 : MUX2_X1 port map( A => n64, B => n60, S => n1389, Z => n1393);
   U1553 : INV_X1 port map( A => intadd_0_A_16_port, ZN => n1390);
   U1554 : MUX2_X1 port map( A => intadd_0_A_16_port, B => n1390, S => 
                           intadd_0_n1, Z => n1391);
   U1555 : XOR2_X1 port map( A => intadd_1_n1, B => n1391, Z => n1392);
   U1556 : XNOR2_X1 port map( A => n1393, B => n1392, ZN => n1394);
   U1557 : OAI22_X1 port map( A1 => n1397, A2 => n1396, B1 => n1395, B2 => 
                           n1394, ZN => n1398);
   U1558 : AOI211_X1 port map( C1 => OP_B_31_port, C2 => n1400, A => n1399, B 
                           => n1398, ZN => n1402);
   U1559 : NAND4_X1 port map( A1 => n1404, A2 => n1403, A3 => n1402, A4 => 
                           n1401, ZN => Y(31));
   U1560 : OAI22_X1 port map( A1 => OPC(6), A2 => n1406, B1 => n1405, B2 => 
                           n1410, ZN => N282);
   U1561 : OAI22_X1 port map( A1 => n1410, A2 => n1409, B1 => n1408, B2 => 
                           n1407, ZN => N283);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( CLK, RST : in std_logic);

end DLX;

architecture SYN_DLX_RTL of DLX is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component RF_N32_NA5
      port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
            ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component ALU_N32_NB8
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
            std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);
            Z : out std_logic);
   end component;
   
   component DLX_DRAM_N256_NW32
      port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector 
            (31 downto 0);  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component DLX_IRAM_RAM_DEPTH256_I_SIZE32
      port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  
            DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, 
      IR_26_port, IR_10_port, IR_9_port, IR_8_port, IR_7_port, IR_6_port, 
      IR_5_port, IR_4_port, IR_3_port, IR_2_port, IR_1_port, IR_0_port, 
      ALU_OPCODE_i_0_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_4_port, ALU_OPCODE_i_5_port, 
      ALU_OPCODE_i_6_port, IR_BUS_31_port, IR_BUS_30_port, IR_BUS_29_port, 
      IR_BUS_28_port, IR_BUS_27_port, IR_BUS_26_port, IR_BUS_25_port, 
      IR_BUS_24_port, IR_BUS_23_port, IR_BUS_22_port, IR_BUS_21_port, 
      IR_BUS_20_port, IR_BUS_19_port, IR_BUS_18_port, IR_BUS_17_port, 
      IR_BUS_16_port, IR_BUS_15_port, IR_BUS_14_port, IR_BUS_13_port, 
      IR_BUS_12_port, IR_BUS_11_port, IR_BUS_10_port, IR_BUS_9_port, 
      IR_BUS_8_port, IR_BUS_7_port, IR_BUS_6_port, IR_BUS_5_port, IR_BUS_4_port
      , IR_BUS_3_port, IR_BUS_2_port, IR_BUS_1_port, IR_BUS_0_port, 
      DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, DATA_OUT_28_port, 
      DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, DATA_OUT_24_port, 
      DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, 
      DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, 
      DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, 
      DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, 
      DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, 
      DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port, 
      DATA_ADDR_31_port, DATA_ADDR_30_port, DATA_ADDR_29_port, 
      DATA_ADDR_28_port, DATA_ADDR_27_port, DATA_ADDR_26_port, 
      DATA_ADDR_25_port, DATA_ADDR_24_port, DATA_ADDR_23_port, 
      DATA_ADDR_22_port, DATA_ADDR_21_port, DATA_ADDR_20_port, 
      DATA_ADDR_19_port, DATA_ADDR_18_port, DATA_ADDR_17_port, 
      DATA_ADDR_16_port, DATA_ADDR_15_port, DATA_ADDR_14_port, 
      DATA_ADDR_13_port, DATA_ADDR_12_port, DATA_ADDR_11_port, 
      DATA_ADDR_10_port, DATA_ADDR_9_port, DATA_ADDR_8_port, DATA_ADDR_7_port, 
      DATA_ADDR_6_port, DATA_ADDR_5_port, DATA_ADDR_4_port, DATA_ADDR_3_port, 
      DATA_ADDR_2_port, DATA_ADDR_1_port, DATA_ADDR_0_port, DATA_IN_31_port, 
      DATA_IN_30_port, DATA_IN_29_port, DATA_IN_28_port, DATA_IN_27_port, 
      DATA_IN_26_port, DATA_IN_25_port, DATA_IN_24_port, DATA_IN_23_port, 
      DATA_IN_22_port, DATA_IN_21_port, DATA_IN_20_port, DATA_IN_19_port, 
      DATA_IN_18_port, DATA_IN_17_port, DATA_IN_16_port, DATA_IN_15_port, 
      DATA_IN_14_port, DATA_IN_13_port, DATA_IN_12_port, DATA_IN_11_port, 
      DATA_IN_10_port, DATA_IN_9_port, DATA_IN_8_port, DATA_IN_7_port, 
      DATA_IN_6_port, DATA_IN_5_port, DATA_IN_4_port, DATA_IN_3_port, 
      DATA_IN_2_port, DATA_IN_1_port, DATA_IN_0_port, CU_I_aluOpcode2_0_port, 
      CU_I_aluOpcode2_1_port, CU_I_aluOpcode2_2_port, CU_I_aluOpcode2_3_port, 
      CU_I_aluOpcode2_4_port, CU_I_aluOpcode2_5_port, CU_I_aluOpcode2_6_port, 
      CU_I_aluOpcode1_0_port, CU_I_aluOpcode1_1_port, CU_I_aluOpcode1_2_port, 
      CU_I_aluOpcode1_3_port, CU_I_aluOpcode1_4_port, CU_I_aluOpcode1_5_port, 
      CU_I_aluOpcode1_6_port, DATAPATH_I_ALU_OUTPUT_0_port, 
      DATAPATH_I_ALU_OUTPUT_1_port, DATAPATH_I_ALU_OUTPUT_2_port, 
      DATAPATH_I_ALU_OUTPUT_3_port, DATAPATH_I_ALU_OUTPUT_4_port, 
      DATAPATH_I_ALU_OUTPUT_5_port, DATAPATH_I_ALU_OUTPUT_6_port, 
      DATAPATH_I_ALU_OUTPUT_7_port, DATAPATH_I_ALU_OUTPUT_8_port, 
      DATAPATH_I_ALU_OUTPUT_9_port, DATAPATH_I_ALU_OUTPUT_10_port, 
      DATAPATH_I_ALU_OUTPUT_11_port, DATAPATH_I_ALU_OUTPUT_12_port, 
      DATAPATH_I_ALU_OUTPUT_13_port, DATAPATH_I_ALU_OUTPUT_14_port, 
      DATAPATH_I_ALU_OUTPUT_15_port, DATAPATH_I_ALU_OUTPUT_16_port, 
      DATAPATH_I_ALU_OUTPUT_17_port, DATAPATH_I_ALU_OUTPUT_18_port, 
      DATAPATH_I_ALU_OUTPUT_19_port, DATAPATH_I_ALU_OUTPUT_20_port, 
      DATAPATH_I_ALU_OUTPUT_21_port, DATAPATH_I_ALU_OUTPUT_22_port, 
      DATAPATH_I_ALU_OUTPUT_23_port, DATAPATH_I_ALU_OUTPUT_24_port, 
      DATAPATH_I_ALU_OUTPUT_25_port, DATAPATH_I_ALU_OUTPUT_26_port, 
      DATAPATH_I_ALU_OUTPUT_27_port, DATAPATH_I_ALU_OUTPUT_28_port, 
      DATAPATH_I_ALU_OUTPUT_29_port, DATAPATH_I_ALU_OUTPUT_30_port, 
      DATAPATH_I_ALU_OUTPUT_31_port, DATAPATH_I_RF_OUT2_0_port, 
      DATAPATH_I_RF_OUT2_1_port, DATAPATH_I_RF_OUT2_2_port, 
      DATAPATH_I_RF_OUT2_3_port, DATAPATH_I_RF_OUT2_4_port, 
      DATAPATH_I_RF_OUT2_5_port, DATAPATH_I_RF_OUT2_6_port, 
      DATAPATH_I_RF_OUT2_7_port, DATAPATH_I_RF_OUT2_8_port, 
      DATAPATH_I_RF_OUT2_9_port, DATAPATH_I_RF_OUT2_10_port, 
      DATAPATH_I_RF_OUT2_11_port, DATAPATH_I_RF_OUT2_12_port, 
      DATAPATH_I_RF_OUT2_13_port, DATAPATH_I_RF_OUT2_14_port, 
      DATAPATH_I_RF_OUT2_15_port, DATAPATH_I_RF_OUT2_16_port, 
      DATAPATH_I_RF_OUT2_17_port, DATAPATH_I_RF_OUT2_18_port, 
      DATAPATH_I_RF_OUT2_19_port, DATAPATH_I_RF_OUT2_20_port, 
      DATAPATH_I_RF_OUT2_21_port, DATAPATH_I_RF_OUT2_22_port, 
      DATAPATH_I_RF_OUT2_23_port, DATAPATH_I_RF_OUT2_24_port, 
      DATAPATH_I_RF_OUT2_25_port, DATAPATH_I_RF_OUT2_26_port, 
      DATAPATH_I_RF_OUT2_27_port, DATAPATH_I_RF_OUT2_28_port, 
      DATAPATH_I_RF_OUT2_29_port, DATAPATH_I_RF_OUT2_30_port, 
      DATAPATH_I_RF_OUT2_31_port, DATAPATH_I_RF_OUT1_0_port, 
      DATAPATH_I_RF_OUT1_1_port, DATAPATH_I_RF_OUT1_2_port, 
      DATAPATH_I_RF_OUT1_3_port, DATAPATH_I_RF_OUT1_4_port, 
      DATAPATH_I_RF_OUT1_5_port, DATAPATH_I_RF_OUT1_6_port, 
      DATAPATH_I_RF_OUT1_7_port, DATAPATH_I_RF_OUT1_8_port, 
      DATAPATH_I_RF_OUT1_9_port, DATAPATH_I_RF_OUT1_10_port, 
      DATAPATH_I_RF_OUT1_11_port, DATAPATH_I_RF_OUT1_12_port, 
      DATAPATH_I_RF_OUT1_13_port, DATAPATH_I_RF_OUT1_14_port, 
      DATAPATH_I_RF_OUT1_15_port, DATAPATH_I_RF_OUT1_16_port, 
      DATAPATH_I_RF_OUT1_17_port, DATAPATH_I_RF_OUT1_18_port, 
      DATAPATH_I_RF_OUT1_19_port, DATAPATH_I_RF_OUT1_20_port, 
      DATAPATH_I_RF_OUT1_21_port, DATAPATH_I_RF_OUT1_22_port, 
      DATAPATH_I_RF_OUT1_23_port, DATAPATH_I_RF_OUT1_24_port, 
      DATAPATH_I_RF_OUT1_25_port, DATAPATH_I_RF_OUT1_26_port, 
      DATAPATH_I_RF_OUT1_27_port, DATAPATH_I_RF_OUT1_28_port, 
      DATAPATH_I_RF_OUT1_29_port, DATAPATH_I_RF_OUT1_30_port, 
      DATAPATH_I_RF_OUT1_31_port, DATAPATH_I_N414, DATAPATH_I_N413, 
      DATAPATH_I_N412, DATAPATH_I_N411, DATAPATH_I_N410, DATAPATH_I_N409, 
      DATAPATH_I_N408, DATAPATH_I_N407, DATAPATH_I_N406, DATAPATH_I_N405, 
      DATAPATH_I_N404, DATAPATH_I_N403, DATAPATH_I_N402, DATAPATH_I_N401, 
      DATAPATH_I_N400, DATAPATH_I_N399, DATAPATH_I_N398, DATAPATH_I_N397, 
      DATAPATH_I_N396, DATAPATH_I_N395, DATAPATH_I_N394, DATAPATH_I_N393, 
      DATAPATH_I_N392, DATAPATH_I_N391, DATAPATH_I_N390, DATAPATH_I_N389, 
      DATAPATH_I_N388, DATAPATH_I_N387, DATAPATH_I_N386, DATAPATH_I_N385, 
      DATAPATH_I_N384, DATAPATH_I_N383, DATAPATH_I_N382, DATAPATH_I_N381, 
      DATAPATH_I_N380, DATAPATH_I_N379, DATAPATH_I_N378, DATAPATH_I_N312, 
      DATAPATH_I_N311, DATAPATH_I_N310, DATAPATH_I_N309, DATAPATH_I_N308, 
      DATAPATH_I_N306, DATAPATH_I_N305, DATAPATH_I_N304, DATAPATH_I_N303, 
      DATAPATH_I_N302, DATAPATH_I_N301, DATAPATH_I_N300, DATAPATH_I_N299, 
      DATAPATH_I_N298, DATAPATH_I_N297, DATAPATH_I_N296, DATAPATH_I_N295, 
      DATAPATH_I_N294, DATAPATH_I_N293, DATAPATH_I_N292, DATAPATH_I_N291, 
      DATAPATH_I_N290, DATAPATH_I_N289, DATAPATH_I_N288, DATAPATH_I_N287, 
      DATAPATH_I_N286, DATAPATH_I_N285, DATAPATH_I_N284, DATAPATH_I_N283, 
      DATAPATH_I_N282, DATAPATH_I_N281, DATAPATH_I_N280, DATAPATH_I_N279, 
      DATAPATH_I_N278, DATAPATH_I_N277, DATAPATH_I_N276, DATAPATH_I_N275, 
      DATAPATH_I_N274, DATAPATH_I_N273, DATAPATH_I_N272, DATAPATH_I_N271, 
      DATAPATH_I_N270, DATAPATH_I_N269, DATAPATH_I_N268, DATAPATH_I_N267, 
      DATAPATH_I_N266, DATAPATH_I_N265, DATAPATH_I_N264, DATAPATH_I_N263, 
      DATAPATH_I_N262, DATAPATH_I_N261, DATAPATH_I_N260, DATAPATH_I_N259, 
      DATAPATH_I_N258, DATAPATH_I_N257, DATAPATH_I_N256, DATAPATH_I_N255, 
      DATAPATH_I_N254, DATAPATH_I_N253, DATAPATH_I_N252, DATAPATH_I_N251, 
      DATAPATH_I_N250, DATAPATH_I_N249, DATAPATH_I_N248, DATAPATH_I_N247, 
      DATAPATH_I_N246, DATAPATH_I_N245, DATAPATH_I_N244, DATAPATH_I_N243, 
      DATAPATH_I_N177, DATAPATH_I_N176, DATAPATH_I_N175, DATAPATH_I_N174, 
      DATAPATH_I_N173, DATAPATH_I_N172, DATAPATH_I_N171, DATAPATH_I_N170, 
      DATAPATH_I_N169, DATAPATH_I_N168, DATAPATH_I_N167, DATAPATH_I_N166, 
      DATAPATH_I_N165, DATAPATH_I_N164, DATAPATH_I_N163, DATAPATH_I_N162, 
      DATAPATH_I_N161, DATAPATH_I_N160, DATAPATH_I_N159, DATAPATH_I_N158, 
      DATAPATH_I_N157, DATAPATH_I_N156, DATAPATH_I_N155, DATAPATH_I_N154, 
      DATAPATH_I_N153, DATAPATH_I_N152, DATAPATH_I_N151, DATAPATH_I_N150, 
      DATAPATH_I_N149, DATAPATH_I_N148, DATAPATH_I_N147, DATAPATH_I_N146, 
      DATAPATH_I_N145, DATAPATH_I_N144, DATAPATH_I_N143, DATAPATH_I_N142, 
      DATAPATH_I_N141, DATAPATH_I_N140, DATAPATH_I_N139, DATAPATH_I_N138, 
      DATAPATH_I_N137, DATAPATH_I_N136, DATAPATH_I_N135, DATAPATH_I_N134, 
      DATAPATH_I_N133, DATAPATH_I_N132, DATAPATH_I_N131, DATAPATH_I_N130, 
      DATAPATH_I_N129, DATAPATH_I_N128, DATAPATH_I_N127, DATAPATH_I_N126, 
      DATAPATH_I_N125, DATAPATH_I_N124, DATAPATH_I_N123, DATAPATH_I_N122, 
      DATAPATH_I_N121, DATAPATH_I_N120, DATAPATH_I_N119, DATAPATH_I_N118, 
      DATAPATH_I_N117, DATAPATH_I_N116, DATAPATH_I_N115, DATAPATH_I_N114, 
      DATAPATH_I_N113, DATAPATH_I_N112, DATAPATH_I_N111, DATAPATH_I_N110, 
      DATAPATH_I_N109, DATAPATH_I_N65, DATAPATH_I_N64, DATAPATH_I_N63, 
      DATAPATH_I_N62, DATAPATH_I_N61, DATAPATH_I_N60, DATAPATH_I_N59, 
      DATAPATH_I_N58, DATAPATH_I_N57, DATAPATH_I_N56, DATAPATH_I_N55, 
      DATAPATH_I_N54, DATAPATH_I_N53, DATAPATH_I_N52, DATAPATH_I_N51, 
      DATAPATH_I_N50, DATAPATH_I_N49, DATAPATH_I_N48, DATAPATH_I_N47, 
      DATAPATH_I_N46, DATAPATH_I_N45, DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_0_port
      , DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_1_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_2_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_3_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_4_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_5_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_6_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_7_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_8_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_9_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_10_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_11_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_12_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_13_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_14_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_15_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_16_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_17_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_18_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_19_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_20_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_21_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_22_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_23_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_24_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_25_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_26_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_27_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_28_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_29_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_30_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_31_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_0_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_1_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_2_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_3_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_4_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_5_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_6_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_7_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_8_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_9_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_10_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_11_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_12_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_13_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_14_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_15_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_16_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_17_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_18_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_19_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_20_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_21_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_22_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_23_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_24_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_25_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_26_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_27_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_28_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_29_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_30_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_31_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_0_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_1_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_2_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_3_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_4_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_5_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_6_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_7_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_8_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_9_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_10_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_11_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_12_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_13_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_14_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_15_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_16_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_17_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_18_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_19_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_20_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_21_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_22_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_23_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_24_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_25_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_26_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_27_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_28_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_29_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_30_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_31_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_0_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_1_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_2_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_3_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_4_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_5_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_6_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_7_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_8_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_9_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_10_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_11_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_12_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_13_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_14_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_15_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_16_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_17_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_18_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_19_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_20_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_21_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_22_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_23_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_24_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_25_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_26_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_27_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_28_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_29_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_30_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_31_port, DATAPATH_I_ID_EX_RS1_NEXT_0_port, 
      DATAPATH_I_ID_EX_RS1_NEXT_1_port, DATAPATH_I_ID_EX_RS1_NEXT_2_port, 
      DATAPATH_I_ID_EX_RS1_NEXT_3_port, DATAPATH_I_ID_EX_RS1_NEXT_4_port, 
      DATAPATH_I_MEM_WB_RD_0_port, DATAPATH_I_MEM_WB_RD_1_port, 
      DATAPATH_I_MEM_WB_RD_2_port, DATAPATH_I_MEM_WB_RD_3_port, 
      DATAPATH_I_MEM_WB_RD_4_port, DATAPATH_I_MEM_WB_DRAM_OUTPUT_0_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_1_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_2_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_3_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_4_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_5_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_6_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_7_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_8_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_9_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_10_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_11_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_12_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_13_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_14_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_15_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_16_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_17_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_18_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_19_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_20_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_21_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_22_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_23_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_24_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_25_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_26_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_27_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_28_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_29_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_30_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_31_port, DATAPATH_I_MEM_WB_RF_WE, 
      DATAPATH_I_EX_MEM_RD_0_port, DATAPATH_I_EX_MEM_RD_1_port, 
      DATAPATH_I_EX_MEM_RD_2_port, DATAPATH_I_EX_MEM_RD_3_port, 
      DATAPATH_I_EX_MEM_RD_4_port, DATAPATH_I_ID_EX_RF_OUT2_0_port, 
      DATAPATH_I_ID_EX_RF_OUT2_1_port, DATAPATH_I_ID_EX_RF_OUT2_2_port, 
      DATAPATH_I_ID_EX_RF_OUT2_3_port, DATAPATH_I_ID_EX_RF_OUT2_4_port, 
      DATAPATH_I_ID_EX_RF_OUT2_5_port, DATAPATH_I_ID_EX_RF_OUT2_6_port, 
      DATAPATH_I_ID_EX_RF_OUT2_7_port, DATAPATH_I_ID_EX_RF_OUT2_8_port, 
      DATAPATH_I_ID_EX_RF_OUT2_9_port, DATAPATH_I_ID_EX_RF_OUT2_10_port, 
      DATAPATH_I_ID_EX_RF_OUT2_11_port, DATAPATH_I_ID_EX_RF_OUT2_12_port, 
      DATAPATH_I_ID_EX_RF_OUT2_13_port, DATAPATH_I_ID_EX_RF_OUT2_14_port, 
      DATAPATH_I_ID_EX_RF_OUT2_15_port, DATAPATH_I_ID_EX_RF_OUT2_16_port, 
      DATAPATH_I_ID_EX_RF_OUT2_17_port, DATAPATH_I_ID_EX_RF_OUT2_18_port, 
      DATAPATH_I_ID_EX_RF_OUT2_19_port, DATAPATH_I_ID_EX_RF_OUT2_20_port, 
      DATAPATH_I_ID_EX_RF_OUT2_21_port, DATAPATH_I_ID_EX_RF_OUT2_22_port, 
      DATAPATH_I_ID_EX_RF_OUT2_23_port, DATAPATH_I_ID_EX_RF_OUT2_24_port, 
      DATAPATH_I_ID_EX_RF_OUT2_25_port, DATAPATH_I_ID_EX_RF_OUT2_26_port, 
      DATAPATH_I_ID_EX_RF_OUT2_27_port, DATAPATH_I_ID_EX_RF_OUT2_28_port, 
      DATAPATH_I_ID_EX_RF_OUT2_29_port, DATAPATH_I_ID_EX_RF_OUT2_30_port, 
      DATAPATH_I_ID_EX_RF_OUT2_31_port, DATAPATH_I_ID_EX_RF_OUT1_0_port, 
      DATAPATH_I_ID_EX_RF_OUT1_1_port, DATAPATH_I_ID_EX_RF_OUT1_2_port, 
      DATAPATH_I_ID_EX_RF_OUT1_3_port, DATAPATH_I_ID_EX_RF_OUT1_4_port, 
      DATAPATH_I_ID_EX_RF_OUT1_5_port, DATAPATH_I_ID_EX_RF_OUT1_6_port, 
      DATAPATH_I_ID_EX_RF_OUT1_7_port, DATAPATH_I_ID_EX_RF_OUT1_8_port, 
      DATAPATH_I_ID_EX_RF_OUT1_9_port, DATAPATH_I_ID_EX_RF_OUT1_10_port, 
      DATAPATH_I_ID_EX_RF_OUT1_11_port, DATAPATH_I_ID_EX_RF_OUT1_12_port, 
      DATAPATH_I_ID_EX_RF_OUT1_13_port, DATAPATH_I_ID_EX_RF_OUT1_14_port, 
      DATAPATH_I_ID_EX_RF_OUT1_15_port, DATAPATH_I_ID_EX_RF_OUT1_16_port, 
      DATAPATH_I_ID_EX_RF_OUT1_17_port, DATAPATH_I_ID_EX_RF_OUT1_18_port, 
      DATAPATH_I_ID_EX_RF_OUT1_19_port, DATAPATH_I_ID_EX_RF_OUT1_20_port, 
      DATAPATH_I_ID_EX_RF_OUT1_21_port, DATAPATH_I_ID_EX_RF_OUT1_22_port, 
      DATAPATH_I_ID_EX_RF_OUT1_23_port, DATAPATH_I_ID_EX_RF_OUT1_24_port, 
      DATAPATH_I_ID_EX_RF_OUT1_25_port, DATAPATH_I_ID_EX_RF_OUT1_26_port, 
      DATAPATH_I_ID_EX_RF_OUT1_27_port, DATAPATH_I_ID_EX_RF_OUT1_28_port, 
      DATAPATH_I_ID_EX_RF_OUT1_29_port, DATAPATH_I_ID_EX_RF_OUT1_30_port, 
      DATAPATH_I_ID_EX_RF_OUT1_31_port, DATAPATH_I_ID_EX_RD_0_port, 
      DATAPATH_I_ID_EX_RD_1_port, DATAPATH_I_ID_EX_RD_2_port, 
      DATAPATH_I_ID_EX_RD_3_port, DATAPATH_I_ID_EX_RD_4_port, 
      DATAPATH_I_IF_ID_IR_11_port, DATAPATH_I_IF_ID_IR_12_port, 
      DATAPATH_I_IF_ID_IR_13_port, DATAPATH_I_IF_ID_IR_14_port, 
      DATAPATH_I_IF_ID_IR_15_port, DATAPATH_I_IF_ID_IR_16_port, 
      DATAPATH_I_IF_ID_IR_17_port, DATAPATH_I_IF_ID_IR_18_port, 
      DATAPATH_I_IF_ID_IR_19_port, DATAPATH_I_IF_ID_IR_20_port, 
      DATAPATH_I_IF_ID_IR_21_port, DATAPATH_I_IF_ID_IR_22_port, 
      DATAPATH_I_IF_ID_IR_23_port, DATAPATH_I_IF_ID_IR_24_port, 
      DATAPATH_I_IF_ID_IR_25_port, DATAPATH_I_IF_ID_IR_26_port, 
      DATAPATH_I_IF_ID_IR_27_port, DATAPATH_I_IF_ID_IR_28_port, 
      DATAPATH_I_IF_ID_IR_29_port, DATAPATH_I_IF_ID_IR_30_port, 
      DATAPATH_I_IF_ID_IR_31_port, DATAPATH_I_n29, DATAPATH_I_n28, 
      DATAPATH_I_n27, DATAPATH_I_n26, DATAPATH_I_n25, DATAPATH_I_n24, 
      DATAPATH_I_n23, DATAPATH_I_n22, DATAPATH_I_n21, DATAPATH_I_n20, 
      DATAPATH_I_n19, DATAPATH_I_n18, DATAPATH_I_n17, DATAPATH_I_n16, 
      DATAPATH_I_n15, DATAPATH_I_LATCH_LMD_LDI_0_N3, 
      DATAPATH_I_LATCH_LMD_LDI_1_N3, DATAPATH_I_LATCH_LMD_LDI_2_N3, 
      DATAPATH_I_LATCH_LMD_LDI_3_N3, DATAPATH_I_LATCH_LMD_LDI_4_N3, 
      DATAPATH_I_LATCH_LMD_LDI_5_N3, DATAPATH_I_LATCH_LMD_LDI_6_N3, 
      DATAPATH_I_LATCH_LMD_LDI_7_N3, DATAPATH_I_LATCH_LMD_LDI_8_N3, 
      DATAPATH_I_LATCH_LMD_LDI_9_N3, DATAPATH_I_LATCH_LMD_LDI_10_N3, 
      DATAPATH_I_LATCH_LMD_LDI_11_N3, DATAPATH_I_LATCH_LMD_LDI_12_N3, 
      DATAPATH_I_LATCH_LMD_LDI_13_N3, DATAPATH_I_LATCH_LMD_LDI_14_N3, 
      DATAPATH_I_LATCH_LMD_LDI_15_N3, DATAPATH_I_LATCH_LMD_LDI_16_N3, 
      DATAPATH_I_LATCH_LMD_LDI_17_N3, DATAPATH_I_LATCH_LMD_LDI_18_N3, 
      DATAPATH_I_LATCH_LMD_LDI_19_N3, DATAPATH_I_LATCH_LMD_LDI_20_N3, 
      DATAPATH_I_LATCH_LMD_LDI_21_N3, DATAPATH_I_LATCH_LMD_LDI_22_N3, 
      DATAPATH_I_LATCH_LMD_LDI_23_N3, DATAPATH_I_LATCH_LMD_LDI_24_N3, 
      DATAPATH_I_LATCH_LMD_LDI_25_N3, DATAPATH_I_LATCH_LMD_LDI_26_N3, 
      DATAPATH_I_LATCH_LMD_LDI_27_N3, DATAPATH_I_LATCH_LMD_LDI_28_N3, 
      DATAPATH_I_LATCH_LMD_LDI_29_N3, DATAPATH_I_LATCH_LMD_LDI_30_N3, 
      DATAPATH_I_LATCH_LMD_LDI_31_N3, DATAPATH_I_LATCH_ALUOUT_LDI_0_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_1_N3, DATAPATH_I_LATCH_ALUOUT_LDI_2_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_3_N3, DATAPATH_I_LATCH_ALUOUT_LDI_4_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_5_N3, DATAPATH_I_LATCH_ALUOUT_LDI_6_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_7_N3, DATAPATH_I_LATCH_ALUOUT_LDI_8_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_9_N3, DATAPATH_I_LATCH_ALUOUT_LDI_10_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_11_N3, DATAPATH_I_LATCH_ALUOUT_LDI_12_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_13_N3, DATAPATH_I_LATCH_ALUOUT_LDI_14_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_15_N3, DATAPATH_I_LATCH_ALUOUT_LDI_16_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_17_N3, DATAPATH_I_LATCH_ALUOUT_LDI_18_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_19_N3, DATAPATH_I_LATCH_ALUOUT_LDI_20_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_21_N3, DATAPATH_I_LATCH_ALUOUT_LDI_22_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_23_N3, DATAPATH_I_LATCH_ALUOUT_LDI_24_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_25_N3, DATAPATH_I_LATCH_ALUOUT_LDI_26_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_27_N3, DATAPATH_I_LATCH_ALUOUT_LDI_28_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_29_N3, DATAPATH_I_LATCH_ALUOUT_LDI_30_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_31_N3, DATAPATH_I_LATCH_RF2_LDI_0_N3, 
      DATAPATH_I_LATCH_RF2_LDI_1_N3, DATAPATH_I_LATCH_RF2_LDI_2_N3, 
      DATAPATH_I_LATCH_RF2_LDI_3_N3, DATAPATH_I_LATCH_RF2_LDI_4_N3, 
      DATAPATH_I_LATCH_RF2_LDI_5_N3, DATAPATH_I_LATCH_RF2_LDI_6_N3, 
      DATAPATH_I_LATCH_RF2_LDI_7_N3, DATAPATH_I_LATCH_RF2_LDI_8_N3, 
      DATAPATH_I_LATCH_RF2_LDI_9_N3, DATAPATH_I_LATCH_RF2_LDI_10_N3, 
      DATAPATH_I_LATCH_RF2_LDI_11_N3, DATAPATH_I_LATCH_RF2_LDI_12_N3, 
      DATAPATH_I_LATCH_RF2_LDI_13_N3, DATAPATH_I_LATCH_RF2_LDI_14_N3, 
      DATAPATH_I_LATCH_RF2_LDI_15_N3, DATAPATH_I_LATCH_RF2_LDI_16_N3, 
      DATAPATH_I_LATCH_RF2_LDI_17_N3, DATAPATH_I_LATCH_RF2_LDI_18_N3, 
      DATAPATH_I_LATCH_RF2_LDI_19_N3, DATAPATH_I_LATCH_RF2_LDI_20_N3, 
      DATAPATH_I_LATCH_RF2_LDI_21_N3, DATAPATH_I_LATCH_RF2_LDI_22_N3, 
      DATAPATH_I_LATCH_RF2_LDI_23_N3, DATAPATH_I_LATCH_RF2_LDI_24_N3, 
      DATAPATH_I_LATCH_RF2_LDI_25_N3, DATAPATH_I_LATCH_RF2_LDI_26_N3, 
      DATAPATH_I_LATCH_RF2_LDI_27_N3, DATAPATH_I_LATCH_RF2_LDI_28_N3, 
      DATAPATH_I_LATCH_RF2_LDI_29_N3, DATAPATH_I_LATCH_RF2_LDI_30_N3, 
      DATAPATH_I_LATCH_RF2_LDI_31_N3, DATAPATH_I_LATCH_RF1_LDI_0_N3, 
      DATAPATH_I_LATCH_RF1_LDI_1_N3, DATAPATH_I_LATCH_RF1_LDI_2_N3, 
      DATAPATH_I_LATCH_RF1_LDI_3_N3, DATAPATH_I_LATCH_RF1_LDI_4_N3, 
      DATAPATH_I_LATCH_RF1_LDI_5_N3, DATAPATH_I_LATCH_RF1_LDI_6_N3, 
      DATAPATH_I_LATCH_RF1_LDI_7_N3, DATAPATH_I_LATCH_RF1_LDI_8_N3, 
      DATAPATH_I_LATCH_RF1_LDI_9_N3, DATAPATH_I_LATCH_RF1_LDI_10_N3, 
      DATAPATH_I_LATCH_RF1_LDI_11_N3, DATAPATH_I_LATCH_RF1_LDI_12_N3, 
      DATAPATH_I_LATCH_RF1_LDI_13_N3, DATAPATH_I_LATCH_RF1_LDI_14_N3, 
      DATAPATH_I_LATCH_RF1_LDI_15_N3, DATAPATH_I_LATCH_RF1_LDI_16_N3, 
      DATAPATH_I_LATCH_RF1_LDI_17_N3, DATAPATH_I_LATCH_RF1_LDI_18_N3, 
      DATAPATH_I_LATCH_RF1_LDI_19_N3, DATAPATH_I_LATCH_RF1_LDI_20_N3, 
      DATAPATH_I_LATCH_RF1_LDI_21_N3, DATAPATH_I_LATCH_RF1_LDI_22_N3, 
      DATAPATH_I_LATCH_RF1_LDI_23_N3, DATAPATH_I_LATCH_RF1_LDI_24_N3, 
      DATAPATH_I_LATCH_RF1_LDI_25_N3, DATAPATH_I_LATCH_RF1_LDI_26_N3, 
      DATAPATH_I_LATCH_RF1_LDI_27_N3, DATAPATH_I_LATCH_RF1_LDI_28_N3, 
      DATAPATH_I_LATCH_RF1_LDI_29_N3, DATAPATH_I_LATCH_RF1_LDI_30_N3, 
      DATAPATH_I_LATCH_RF1_LDI_31_N3, DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_N3,
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_N3, n285, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, 
      n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, 
      n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
      n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, 
      n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, 
      n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, 
      n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, 
      n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, 
      n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, 
      n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, 
      n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, 
      n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, 
      n_1370 : std_logic;

begin
   
   IRAM_I : DLX_IRAM_RAM_DEPTH256_I_SIZE32 port map( RST => n320, ADDR(31) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(30) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(29) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(28) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(27) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(26) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(25) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(24) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(23) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(22) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(21) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(20) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(19) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(18) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(17) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(16) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(15) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(14) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(13) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(12) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(11) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(10) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(9) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(8) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(7) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(6) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(5) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(4) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(3) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(2) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(1) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(0) => 
                           DATAPATH_I_MEM_WB_RF_WE, DOUT(31) => IR_BUS_31_port,
                           DOUT(30) => IR_BUS_30_port, DOUT(29) => 
                           IR_BUS_29_port, DOUT(28) => IR_BUS_28_port, DOUT(27)
                           => IR_BUS_27_port, DOUT(26) => IR_BUS_26_port, 
                           DOUT(25) => IR_BUS_25_port, DOUT(24) => 
                           IR_BUS_24_port, DOUT(23) => IR_BUS_23_port, DOUT(22)
                           => IR_BUS_22_port, DOUT(21) => IR_BUS_21_port, 
                           DOUT(20) => IR_BUS_20_port, DOUT(19) => 
                           IR_BUS_19_port, DOUT(18) => IR_BUS_18_port, DOUT(17)
                           => IR_BUS_17_port, DOUT(16) => IR_BUS_16_port, 
                           DOUT(15) => IR_BUS_15_port, DOUT(14) => 
                           IR_BUS_14_port, DOUT(13) => IR_BUS_13_port, DOUT(12)
                           => IR_BUS_12_port, DOUT(11) => IR_BUS_11_port, 
                           DOUT(10) => IR_BUS_10_port, DOUT(9) => IR_BUS_9_port
                           , DOUT(8) => IR_BUS_8_port, DOUT(7) => IR_BUS_7_port
                           , DOUT(6) => IR_BUS_6_port, DOUT(5) => IR_BUS_5_port
                           , DOUT(4) => IR_BUS_4_port, DOUT(3) => IR_BUS_3_port
                           , DOUT(2) => IR_BUS_2_port, DOUT(1) => IR_BUS_1_port
                           , DOUT(0) => IR_BUS_0_port);
   DRAM_I : DLX_DRAM_N256_NW32 port map( CLK => CLK, RST => n320, RE => 
                           DATAPATH_I_MEM_WB_RF_WE, WE => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(31) => 
                           DATA_ADDR_31_port, ADDR(30) => DATA_ADDR_30_port, 
                           ADDR(29) => DATA_ADDR_29_port, ADDR(28) => 
                           DATA_ADDR_28_port, ADDR(27) => DATA_ADDR_27_port, 
                           ADDR(26) => DATA_ADDR_26_port, ADDR(25) => 
                           DATA_ADDR_25_port, ADDR(24) => DATA_ADDR_24_port, 
                           ADDR(23) => DATA_ADDR_23_port, ADDR(22) => 
                           DATA_ADDR_22_port, ADDR(21) => DATA_ADDR_21_port, 
                           ADDR(20) => DATA_ADDR_20_port, ADDR(19) => 
                           DATA_ADDR_19_port, ADDR(18) => DATA_ADDR_18_port, 
                           ADDR(17) => DATA_ADDR_17_port, ADDR(16) => 
                           DATA_ADDR_16_port, ADDR(15) => DATA_ADDR_15_port, 
                           ADDR(14) => DATA_ADDR_14_port, ADDR(13) => 
                           DATA_ADDR_13_port, ADDR(12) => DATA_ADDR_12_port, 
                           ADDR(11) => DATA_ADDR_11_port, ADDR(10) => 
                           DATA_ADDR_10_port, ADDR(9) => DATA_ADDR_9_port, 
                           ADDR(8) => DATA_ADDR_8_port, ADDR(7) => 
                           DATA_ADDR_7_port, ADDR(6) => DATA_ADDR_6_port, 
                           ADDR(5) => DATA_ADDR_5_port, ADDR(4) => 
                           DATA_ADDR_4_port, ADDR(3) => DATA_ADDR_3_port, 
                           ADDR(2) => DATA_ADDR_2_port, ADDR(1) => 
                           DATA_ADDR_1_port, ADDR(0) => DATA_ADDR_0_port, 
                           DIN(31) => DATA_IN_31_port, DIN(30) => 
                           DATA_IN_30_port, DIN(29) => DATA_IN_29_port, DIN(28)
                           => DATA_IN_28_port, DIN(27) => DATA_IN_27_port, 
                           DIN(26) => DATA_IN_26_port, DIN(25) => 
                           DATA_IN_25_port, DIN(24) => DATA_IN_24_port, DIN(23)
                           => DATA_IN_23_port, DIN(22) => DATA_IN_22_port, 
                           DIN(21) => DATA_IN_21_port, DIN(20) => 
                           DATA_IN_20_port, DIN(19) => DATA_IN_19_port, DIN(18)
                           => DATA_IN_18_port, DIN(17) => DATA_IN_17_port, 
                           DIN(16) => DATA_IN_16_port, DIN(15) => 
                           DATA_IN_15_port, DIN(14) => DATA_IN_14_port, DIN(13)
                           => DATA_IN_13_port, DIN(12) => DATA_IN_12_port, 
                           DIN(11) => DATA_IN_11_port, DIN(10) => 
                           DATA_IN_10_port, DIN(9) => DATA_IN_9_port, DIN(8) =>
                           DATA_IN_8_port, DIN(7) => DATA_IN_7_port, DIN(6) => 
                           DATA_IN_6_port, DIN(5) => DATA_IN_5_port, DIN(4) => 
                           DATA_IN_4_port, DIN(3) => DATA_IN_3_port, DIN(2) => 
                           DATA_IN_2_port, DIN(1) => DATA_IN_1_port, DIN(0) => 
                           DATA_IN_0_port, DOUT(31) => DATA_OUT_31_port, 
                           DOUT(30) => DATA_OUT_30_port, DOUT(29) => 
                           DATA_OUT_29_port, DOUT(28) => DATA_OUT_28_port, 
                           DOUT(27) => DATA_OUT_27_port, DOUT(26) => 
                           DATA_OUT_26_port, DOUT(25) => DATA_OUT_25_port, 
                           DOUT(24) => DATA_OUT_24_port, DOUT(23) => 
                           DATA_OUT_23_port, DOUT(22) => DATA_OUT_22_port, 
                           DOUT(21) => DATA_OUT_21_port, DOUT(20) => 
                           DATA_OUT_20_port, DOUT(19) => DATA_OUT_19_port, 
                           DOUT(18) => DATA_OUT_18_port, DOUT(17) => 
                           DATA_OUT_17_port, DOUT(16) => DATA_OUT_16_port, 
                           DOUT(15) => DATA_OUT_15_port, DOUT(14) => 
                           DATA_OUT_14_port, DOUT(13) => DATA_OUT_13_port, 
                           DOUT(12) => DATA_OUT_12_port, DOUT(11) => 
                           DATA_OUT_11_port, DOUT(10) => DATA_OUT_10_port, 
                           DOUT(9) => DATA_OUT_9_port, DOUT(8) => 
                           DATA_OUT_8_port, DOUT(7) => DATA_OUT_7_port, DOUT(6)
                           => DATA_OUT_6_port, DOUT(5) => DATA_OUT_5_port, 
                           DOUT(4) => DATA_OUT_4_port, DOUT(3) => 
                           DATA_OUT_3_port, DOUT(2) => DATA_OUT_2_port, DOUT(1)
                           => DATA_OUT_1_port, DOUT(0) => DATA_OUT_0_port);
   DATAPATH_I_ARITHMETIC_LOGIC_UNIT : ALU_N32_NB8 port map( OP1(31) => 
                           DATAPATH_I_ID_EX_RF_OUT1_31_port, OP1(30) => 
                           DATAPATH_I_ID_EX_RF_OUT1_30_port, OP1(29) => 
                           DATAPATH_I_ID_EX_RF_OUT1_29_port, OP1(28) => 
                           DATAPATH_I_ID_EX_RF_OUT1_28_port, OP1(27) => 
                           DATAPATH_I_ID_EX_RF_OUT1_27_port, OP1(26) => 
                           DATAPATH_I_ID_EX_RF_OUT1_26_port, OP1(25) => 
                           DATAPATH_I_ID_EX_RF_OUT1_25_port, OP1(24) => 
                           DATAPATH_I_ID_EX_RF_OUT1_24_port, OP1(23) => 
                           DATAPATH_I_ID_EX_RF_OUT1_23_port, OP1(22) => 
                           DATAPATH_I_ID_EX_RF_OUT1_22_port, OP1(21) => 
                           DATAPATH_I_ID_EX_RF_OUT1_21_port, OP1(20) => 
                           DATAPATH_I_ID_EX_RF_OUT1_20_port, OP1(19) => 
                           DATAPATH_I_ID_EX_RF_OUT1_19_port, OP1(18) => 
                           DATAPATH_I_ID_EX_RF_OUT1_18_port, OP1(17) => 
                           DATAPATH_I_ID_EX_RF_OUT1_17_port, OP1(16) => 
                           DATAPATH_I_ID_EX_RF_OUT1_16_port, OP1(15) => 
                           DATAPATH_I_ID_EX_RF_OUT1_15_port, OP1(14) => 
                           DATAPATH_I_ID_EX_RF_OUT1_14_port, OP1(13) => 
                           DATAPATH_I_ID_EX_RF_OUT1_13_port, OP1(12) => 
                           DATAPATH_I_ID_EX_RF_OUT1_12_port, OP1(11) => 
                           DATAPATH_I_ID_EX_RF_OUT1_11_port, OP1(10) => 
                           DATAPATH_I_ID_EX_RF_OUT1_10_port, OP1(9) => 
                           DATAPATH_I_ID_EX_RF_OUT1_9_port, OP1(8) => 
                           DATAPATH_I_ID_EX_RF_OUT1_8_port, OP1(7) => 
                           DATAPATH_I_ID_EX_RF_OUT1_7_port, OP1(6) => 
                           DATAPATH_I_ID_EX_RF_OUT1_6_port, OP1(5) => 
                           DATAPATH_I_ID_EX_RF_OUT1_5_port, OP1(4) => 
                           DATAPATH_I_ID_EX_RF_OUT1_4_port, OP1(3) => 
                           DATAPATH_I_ID_EX_RF_OUT1_3_port, OP1(2) => 
                           DATAPATH_I_ID_EX_RF_OUT1_2_port, OP1(1) => 
                           DATAPATH_I_ID_EX_RF_OUT1_1_port, OP1(0) => 
                           DATAPATH_I_ID_EX_RF_OUT1_0_port, OP2(31) => 
                           DATAPATH_I_ID_EX_RF_OUT2_31_port, OP2(30) => 
                           DATAPATH_I_ID_EX_RF_OUT2_30_port, OP2(29) => 
                           DATAPATH_I_ID_EX_RF_OUT2_29_port, OP2(28) => 
                           DATAPATH_I_ID_EX_RF_OUT2_28_port, OP2(27) => 
                           DATAPATH_I_ID_EX_RF_OUT2_27_port, OP2(26) => 
                           DATAPATH_I_ID_EX_RF_OUT2_26_port, OP2(25) => 
                           DATAPATH_I_ID_EX_RF_OUT2_25_port, OP2(24) => 
                           DATAPATH_I_ID_EX_RF_OUT2_24_port, OP2(23) => 
                           DATAPATH_I_ID_EX_RF_OUT2_23_port, OP2(22) => 
                           DATAPATH_I_ID_EX_RF_OUT2_22_port, OP2(21) => 
                           DATAPATH_I_ID_EX_RF_OUT2_21_port, OP2(20) => 
                           DATAPATH_I_ID_EX_RF_OUT2_20_port, OP2(19) => 
                           DATAPATH_I_ID_EX_RF_OUT2_19_port, OP2(18) => 
                           DATAPATH_I_ID_EX_RF_OUT2_18_port, OP2(17) => 
                           DATAPATH_I_ID_EX_RF_OUT2_17_port, OP2(16) => 
                           DATAPATH_I_ID_EX_RF_OUT2_16_port, OP2(15) => 
                           DATAPATH_I_ID_EX_RF_OUT2_15_port, OP2(14) => 
                           DATAPATH_I_ID_EX_RF_OUT2_14_port, OP2(13) => 
                           DATAPATH_I_ID_EX_RF_OUT2_13_port, OP2(12) => 
                           DATAPATH_I_ID_EX_RF_OUT2_12_port, OP2(11) => 
                           DATAPATH_I_ID_EX_RF_OUT2_11_port, OP2(10) => 
                           DATAPATH_I_ID_EX_RF_OUT2_10_port, OP2(9) => 
                           DATAPATH_I_ID_EX_RF_OUT2_9_port, OP2(8) => 
                           DATAPATH_I_ID_EX_RF_OUT2_8_port, OP2(7) => 
                           DATAPATH_I_ID_EX_RF_OUT2_7_port, OP2(6) => 
                           DATAPATH_I_ID_EX_RF_OUT2_6_port, OP2(5) => 
                           DATAPATH_I_ID_EX_RF_OUT2_5_port, OP2(4) => 
                           DATAPATH_I_ID_EX_RF_OUT2_4_port, OP2(3) => 
                           DATAPATH_I_ID_EX_RF_OUT2_3_port, OP2(2) => 
                           DATAPATH_I_ID_EX_RF_OUT2_2_port, OP2(1) => 
                           DATAPATH_I_ID_EX_RF_OUT2_1_port, OP2(0) => 
                           DATAPATH_I_ID_EX_RF_OUT2_0_port, OPC(0) => 
                           ALU_OPCODE_i_0_port, OPC(1) => ALU_OPCODE_i_1_port, 
                           OPC(2) => ALU_OPCODE_i_2_port, OPC(3) => 
                           ALU_OPCODE_i_3_port, OPC(4) => ALU_OPCODE_i_4_port, 
                           OPC(5) => ALU_OPCODE_i_5_port, OPC(6) => 
                           ALU_OPCODE_i_6_port, Y(31) => 
                           DATAPATH_I_ALU_OUTPUT_31_port, Y(30) => 
                           DATAPATH_I_ALU_OUTPUT_30_port, Y(29) => 
                           DATAPATH_I_ALU_OUTPUT_29_port, Y(28) => 
                           DATAPATH_I_ALU_OUTPUT_28_port, Y(27) => 
                           DATAPATH_I_ALU_OUTPUT_27_port, Y(26) => 
                           DATAPATH_I_ALU_OUTPUT_26_port, Y(25) => 
                           DATAPATH_I_ALU_OUTPUT_25_port, Y(24) => 
                           DATAPATH_I_ALU_OUTPUT_24_port, Y(23) => 
                           DATAPATH_I_ALU_OUTPUT_23_port, Y(22) => 
                           DATAPATH_I_ALU_OUTPUT_22_port, Y(21) => 
                           DATAPATH_I_ALU_OUTPUT_21_port, Y(20) => 
                           DATAPATH_I_ALU_OUTPUT_20_port, Y(19) => 
                           DATAPATH_I_ALU_OUTPUT_19_port, Y(18) => 
                           DATAPATH_I_ALU_OUTPUT_18_port, Y(17) => 
                           DATAPATH_I_ALU_OUTPUT_17_port, Y(16) => 
                           DATAPATH_I_ALU_OUTPUT_16_port, Y(15) => 
                           DATAPATH_I_ALU_OUTPUT_15_port, Y(14) => 
                           DATAPATH_I_ALU_OUTPUT_14_port, Y(13) => 
                           DATAPATH_I_ALU_OUTPUT_13_port, Y(12) => 
                           DATAPATH_I_ALU_OUTPUT_12_port, Y(11) => 
                           DATAPATH_I_ALU_OUTPUT_11_port, Y(10) => 
                           DATAPATH_I_ALU_OUTPUT_10_port, Y(9) => 
                           DATAPATH_I_ALU_OUTPUT_9_port, Y(8) => 
                           DATAPATH_I_ALU_OUTPUT_8_port, Y(7) => 
                           DATAPATH_I_ALU_OUTPUT_7_port, Y(6) => 
                           DATAPATH_I_ALU_OUTPUT_6_port, Y(5) => 
                           DATAPATH_I_ALU_OUTPUT_5_port, Y(4) => 
                           DATAPATH_I_ALU_OUTPUT_4_port, Y(3) => 
                           DATAPATH_I_ALU_OUTPUT_3_port, Y(2) => 
                           DATAPATH_I_ALU_OUTPUT_2_port, Y(1) => 
                           DATAPATH_I_ALU_OUTPUT_1_port, Y(0) => 
                           DATAPATH_I_ALU_OUTPUT_0_port, Z => n_1171);
   DATAPATH_I_REGISTER_FILE : RF_N32_NA5 port map( RST => n317, EN => n285, 
                           EN_RD1 => n285, EN_RD2 => n285, EN_WR => 
                           DATAPATH_I_MEM_WB_RF_WE, ADD_RD1(4) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_4_port, ADD_RD1(3) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_3_port, ADD_RD1(2) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_2_port, ADD_RD1(1) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_1_port, ADD_RD1(0) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_0_port, ADD_RD2(4) => n335
                           , ADD_RD2(3) => n333, ADD_RD2(2) => n332, ADD_RD2(1)
                           => n334, ADD_RD2(0) => n331, ADD_WR(4) => 
                           DATAPATH_I_MEM_WB_RD_4_port, ADD_WR(3) => 
                           DATAPATH_I_MEM_WB_RD_3_port, ADD_WR(2) => 
                           DATAPATH_I_MEM_WB_RD_2_port, ADD_WR(1) => 
                           DATAPATH_I_MEM_WB_RD_1_port, ADD_WR(0) => 
                           DATAPATH_I_MEM_WB_RD_0_port, DATAIN(31) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_31_port, DATAIN(30) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_30_port, DATAIN(29) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_29_port, DATAIN(28) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_28_port, DATAIN(27) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_27_port, DATAIN(26) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_26_port, DATAIN(25) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_25_port, DATAIN(24) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_24_port, DATAIN(23) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_23_port, DATAIN(22) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_22_port, DATAIN(21) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_21_port, DATAIN(20) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_20_port, DATAIN(19) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_19_port, DATAIN(18) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_18_port, DATAIN(17) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_17_port, DATAIN(16) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_16_port, DATAIN(15) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_15_port, DATAIN(14) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_14_port, DATAIN(13) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_13_port, DATAIN(12) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_12_port, DATAIN(11) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_11_port, DATAIN(10) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_10_port, DATAIN(9) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_9_port, DATAIN(8) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_8_port, DATAIN(7) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_7_port, DATAIN(6) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_6_port, DATAIN(5) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_5_port, DATAIN(4) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_4_port, DATAIN(3) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_3_port, DATAIN(2) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_2_port, DATAIN(1) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_1_port, DATAIN(0) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_0_port, OUT1(31) => 
                           DATAPATH_I_RF_OUT1_31_port, OUT1(30) => 
                           DATAPATH_I_RF_OUT1_30_port, OUT1(29) => 
                           DATAPATH_I_RF_OUT1_29_port, OUT1(28) => 
                           DATAPATH_I_RF_OUT1_28_port, OUT1(27) => 
                           DATAPATH_I_RF_OUT1_27_port, OUT1(26) => 
                           DATAPATH_I_RF_OUT1_26_port, OUT1(25) => 
                           DATAPATH_I_RF_OUT1_25_port, OUT1(24) => 
                           DATAPATH_I_RF_OUT1_24_port, OUT1(23) => 
                           DATAPATH_I_RF_OUT1_23_port, OUT1(22) => 
                           DATAPATH_I_RF_OUT1_22_port, OUT1(21) => 
                           DATAPATH_I_RF_OUT1_21_port, OUT1(20) => 
                           DATAPATH_I_RF_OUT1_20_port, OUT1(19) => 
                           DATAPATH_I_RF_OUT1_19_port, OUT1(18) => 
                           DATAPATH_I_RF_OUT1_18_port, OUT1(17) => 
                           DATAPATH_I_RF_OUT1_17_port, OUT1(16) => 
                           DATAPATH_I_RF_OUT1_16_port, OUT1(15) => 
                           DATAPATH_I_RF_OUT1_15_port, OUT1(14) => 
                           DATAPATH_I_RF_OUT1_14_port, OUT1(13) => 
                           DATAPATH_I_RF_OUT1_13_port, OUT1(12) => 
                           DATAPATH_I_RF_OUT1_12_port, OUT1(11) => 
                           DATAPATH_I_RF_OUT1_11_port, OUT1(10) => 
                           DATAPATH_I_RF_OUT1_10_port, OUT1(9) => 
                           DATAPATH_I_RF_OUT1_9_port, OUT1(8) => 
                           DATAPATH_I_RF_OUT1_8_port, OUT1(7) => 
                           DATAPATH_I_RF_OUT1_7_port, OUT1(6) => 
                           DATAPATH_I_RF_OUT1_6_port, OUT1(5) => 
                           DATAPATH_I_RF_OUT1_5_port, OUT1(4) => 
                           DATAPATH_I_RF_OUT1_4_port, OUT1(3) => 
                           DATAPATH_I_RF_OUT1_3_port, OUT1(2) => 
                           DATAPATH_I_RF_OUT1_2_port, OUT1(1) => 
                           DATAPATH_I_RF_OUT1_1_port, OUT1(0) => 
                           DATAPATH_I_RF_OUT1_0_port, OUT2(31) => 
                           DATAPATH_I_RF_OUT2_31_port, OUT2(30) => 
                           DATAPATH_I_RF_OUT2_30_port, OUT2(29) => 
                           DATAPATH_I_RF_OUT2_29_port, OUT2(28) => 
                           DATAPATH_I_RF_OUT2_28_port, OUT2(27) => 
                           DATAPATH_I_RF_OUT2_27_port, OUT2(26) => 
                           DATAPATH_I_RF_OUT2_26_port, OUT2(25) => 
                           DATAPATH_I_RF_OUT2_25_port, OUT2(24) => 
                           DATAPATH_I_RF_OUT2_24_port, OUT2(23) => 
                           DATAPATH_I_RF_OUT2_23_port, OUT2(22) => 
                           DATAPATH_I_RF_OUT2_22_port, OUT2(21) => 
                           DATAPATH_I_RF_OUT2_21_port, OUT2(20) => 
                           DATAPATH_I_RF_OUT2_20_port, OUT2(19) => 
                           DATAPATH_I_RF_OUT2_19_port, OUT2(18) => 
                           DATAPATH_I_RF_OUT2_18_port, OUT2(17) => 
                           DATAPATH_I_RF_OUT2_17_port, OUT2(16) => 
                           DATAPATH_I_RF_OUT2_16_port, OUT2(15) => 
                           DATAPATH_I_RF_OUT2_15_port, OUT2(14) => 
                           DATAPATH_I_RF_OUT2_14_port, OUT2(13) => 
                           DATAPATH_I_RF_OUT2_13_port, OUT2(12) => 
                           DATAPATH_I_RF_OUT2_12_port, OUT2(11) => 
                           DATAPATH_I_RF_OUT2_11_port, OUT2(10) => 
                           DATAPATH_I_RF_OUT2_10_port, OUT2(9) => 
                           DATAPATH_I_RF_OUT2_9_port, OUT2(8) => 
                           DATAPATH_I_RF_OUT2_8_port, OUT2(7) => 
                           DATAPATH_I_RF_OUT2_7_port, OUT2(6) => 
                           DATAPATH_I_RF_OUT2_6_port, OUT2(5) => 
                           DATAPATH_I_RF_OUT2_5_port, OUT2(4) => 
                           DATAPATH_I_RF_OUT2_4_port, OUT2(3) => 
                           DATAPATH_I_RF_OUT2_3_port, OUT2(2) => 
                           DATAPATH_I_RF_OUT2_2_port, OUT2(1) => 
                           DATAPATH_I_RF_OUT2_1_port, OUT2(0) => 
                           DATAPATH_I_RF_OUT2_0_port);
   DATAPATH_I_IF_ID_IR_reg_11_inst : DFF_X1 port map( D => DATAPATH_I_N45, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_11_port, QN => 
                           n_1172);
   DATAPATH_I_IF_ID_IR_reg_12_inst : DFF_X1 port map( D => DATAPATH_I_N46, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_12_port, QN => 
                           n_1173);
   DATAPATH_I_IF_ID_IR_reg_13_inst : DFF_X1 port map( D => DATAPATH_I_N47, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_13_port, QN => 
                           n_1174);
   DATAPATH_I_IF_ID_IR_reg_14_inst : DFF_X1 port map( D => DATAPATH_I_N48, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_14_port, QN => 
                           n_1175);
   DATAPATH_I_IF_ID_IR_reg_15_inst : DFF_X1 port map( D => DATAPATH_I_N49, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_15_port, QN => 
                           n_1176);
   DATAPATH_I_IF_ID_IR_reg_16_inst : DFF_X1 port map( D => DATAPATH_I_N50, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_16_port, QN => n479
                           );
   DATAPATH_I_IF_ID_IR_reg_17_inst : DFF_X1 port map( D => DATAPATH_I_N51, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_17_port, QN => n478
                           );
   DATAPATH_I_IF_ID_IR_reg_18_inst : DFF_X1 port map( D => DATAPATH_I_N52, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_18_port, QN => n477
                           );
   DATAPATH_I_IF_ID_IR_reg_19_inst : DFF_X1 port map( D => DATAPATH_I_N53, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_19_port, QN => n476
                           );
   DATAPATH_I_IF_ID_IR_reg_20_inst : DFF_X1 port map( D => DATAPATH_I_N54, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_20_port, QN => n480
                           );
   DATAPATH_I_IF_ID_IR_reg_21_inst : DFF_X1 port map( D => DATAPATH_I_N55, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_21_port, QN => 
                           n_1177);
   DATAPATH_I_IF_ID_IR_reg_22_inst : DFF_X1 port map( D => DATAPATH_I_N56, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_22_port, QN => 
                           n_1178);
   DATAPATH_I_IF_ID_IR_reg_23_inst : DFF_X1 port map( D => DATAPATH_I_N57, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_23_port, QN => 
                           n_1179);
   DATAPATH_I_IF_ID_IR_reg_24_inst : DFF_X1 port map( D => DATAPATH_I_N58, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_24_port, QN => 
                           n_1180);
   DATAPATH_I_IF_ID_IR_reg_25_inst : DFF_X1 port map( D => DATAPATH_I_N59, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_25_port, QN => 
                           n_1181);
   DATAPATH_I_IF_ID_IR_reg_26_inst : DFF_X1 port map( D => DATAPATH_I_N60, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_26_port, QN => n481
                           );
   DATAPATH_I_IF_ID_IR_reg_27_inst : DFF_X1 port map( D => DATAPATH_I_N61, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_27_port, QN => n482
                           );
   DATAPATH_I_IF_ID_IR_reg_28_inst : DFF_X1 port map( D => DATAPATH_I_N62, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_28_port, QN => n483
                           );
   DATAPATH_I_IF_ID_IR_reg_29_inst : DFF_X1 port map( D => DATAPATH_I_N63, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_29_port, QN => n485
                           );
   DATAPATH_I_IF_ID_IR_reg_30_inst : DFF_X1 port map( D => DATAPATH_I_N64, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_30_port, QN => n484
                           );
   DATAPATH_I_IF_ID_IR_reg_31_inst : DFF_X1 port map( D => DATAPATH_I_N65, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_31_port, QN => n486
                           );
   DATAPATH_I_EX_MEM_RD_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N308, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_0_port, QN => 
                           n_1182);
   DATAPATH_I_MEM_WB_RD_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N410, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_0_port, QN => 
                           n_1183);
   DATAPATH_I_EX_MEM_RD_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N309, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_1_port, QN => 
                           n_1184);
   DATAPATH_I_MEM_WB_RD_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N411, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_1_port, QN => 
                           n_1185);
   DATAPATH_I_EX_MEM_RD_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N310, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_2_port, QN => 
                           n_1186);
   DATAPATH_I_MEM_WB_RD_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N412, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_2_port, QN => 
                           n_1187);
   DATAPATH_I_EX_MEM_RD_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N311, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_3_port, QN => 
                           n_1188);
   DATAPATH_I_MEM_WB_RD_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N413, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_3_port, QN => 
                           n_1189);
   DATAPATH_I_EX_MEM_RD_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N312, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_4_port, QN => 
                           n_1190);
   DATAPATH_I_MEM_WB_RD_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N414, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_4_port, QN => 
                           n_1191);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_0_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N275, CK => CLK, Q => DATA_ADDR_0_port, 
                           QN => n_1192);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_1_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N276, CK => CLK, Q => DATA_ADDR_1_port, 
                           QN => n_1193);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_2_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N277, CK => CLK, Q => DATA_ADDR_2_port, 
                           QN => n_1194);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_3_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N278, CK => CLK, Q => DATA_ADDR_3_port, 
                           QN => n_1195);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_4_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N279, CK => CLK, Q => DATA_ADDR_4_port, 
                           QN => n_1196);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_5_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N280, CK => CLK, Q => DATA_ADDR_5_port, 
                           QN => n_1197);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_6_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N281, CK => CLK, Q => DATA_ADDR_6_port, 
                           QN => n_1198);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_7_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N282, CK => CLK, Q => DATA_ADDR_7_port, 
                           QN => n_1199);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_8_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N283, CK => CLK, Q => DATA_ADDR_8_port, 
                           QN => n_1200);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_9_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N284, CK => CLK, Q => DATA_ADDR_9_port, 
                           QN => n_1201);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_10_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N285, CK => CLK, Q => DATA_ADDR_10_port, 
                           QN => n_1202);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_11_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N286, CK => CLK, Q => DATA_ADDR_11_port, 
                           QN => n_1203);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_12_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N287, CK => CLK, Q => DATA_ADDR_12_port, 
                           QN => n_1204);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_13_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N288, CK => CLK, Q => DATA_ADDR_13_port, 
                           QN => n_1205);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_14_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N289, CK => CLK, Q => DATA_ADDR_14_port, 
                           QN => n_1206);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_15_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N290, CK => CLK, Q => DATA_ADDR_15_port, 
                           QN => n_1207);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_16_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N291, CK => CLK, Q => DATA_ADDR_16_port, 
                           QN => n_1208);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_17_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N292, CK => CLK, Q => DATA_ADDR_17_port, 
                           QN => n_1209);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_18_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N293, CK => CLK, Q => DATA_ADDR_18_port, 
                           QN => n_1210);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_19_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N294, CK => CLK, Q => DATA_ADDR_19_port, 
                           QN => n_1211);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_20_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N295, CK => CLK, Q => DATA_ADDR_20_port, 
                           QN => n_1212);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_21_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N296, CK => CLK, Q => DATA_ADDR_21_port, 
                           QN => n_1213);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_22_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N297, CK => CLK, Q => DATA_ADDR_22_port, 
                           QN => n_1214);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_23_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N298, CK => CLK, Q => DATA_ADDR_23_port, 
                           QN => n_1215);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_24_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N299, CK => CLK, Q => DATA_ADDR_24_port, 
                           QN => n_1216);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_25_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N300, CK => CLK, Q => DATA_ADDR_25_port, 
                           QN => n_1217);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_26_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N301, CK => CLK, Q => DATA_ADDR_26_port, 
                           QN => n_1218);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_27_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N302, CK => CLK, Q => DATA_ADDR_27_port, 
                           QN => n_1219);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_28_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N303, CK => CLK, Q => DATA_ADDR_28_port, 
                           QN => n_1220);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_29_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N304, CK => CLK, Q => DATA_ADDR_29_port, 
                           QN => n_1221);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_30_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N305, CK => CLK, Q => DATA_ADDR_30_port, 
                           QN => n_1222);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_31_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N306, CK => CLK, Q => DATA_ADDR_31_port, 
                           QN => n_1223);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_0_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N378, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_0_port, QN => n_1224);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_1_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N379, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_1_port, QN => n_1225);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_2_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N380, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_2_port, QN => n_1226);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_3_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N381, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_3_port, QN => n_1227);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_4_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N382, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_4_port, QN => n_1228);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_5_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N383, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_5_port, QN => n_1229);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_6_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N384, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_6_port, QN => n_1230);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_7_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N385, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_7_port, QN => n_1231);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_8_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N386, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_8_port, QN => n_1232);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_9_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N387, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_9_port, QN => n_1233);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_10_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N388, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_10_port, QN => n_1234)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_11_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N389, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_11_port, QN => n_1235)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_12_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N390, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_12_port, QN => n_1236)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_13_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N391, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_13_port, QN => n_1237)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_14_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N392, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_14_port, QN => n_1238)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_15_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N393, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_15_port, QN => n_1239)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_16_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N394, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_16_port, QN => n_1240)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_17_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N395, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_17_port, QN => n_1241)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_18_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N396, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_18_port, QN => n_1242)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_19_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N397, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_19_port, QN => n_1243)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_20_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N398, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_20_port, QN => n_1244)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_21_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N399, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_21_port, QN => n_1245)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_22_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N400, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_22_port, QN => n_1246)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_23_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N401, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_23_port, QN => n_1247)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_24_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N402, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_24_port, QN => n_1248)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_25_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N403, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_25_port, QN => n_1249)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_26_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N404, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_26_port, QN => n_1250)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_27_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N405, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_27_port, QN => n_1251)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_28_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N406, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_28_port, QN => n_1252)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_29_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N407, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_29_port, QN => n_1253)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_30_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N408, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_30_port, QN => n_1254)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_31_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N409, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_31_port, QN => n_1255)
                           ;
   DATAPATH_I_ID_EX_RF_OUT2_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N146,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_0_port, QN 
                           => n_1256);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N243
                           , CK => CLK, Q => DATA_IN_0_port, QN => n_1257);
   DATAPATH_I_ID_EX_RF_OUT2_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N147,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_1_port, QN 
                           => n_1258);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N244
                           , CK => CLK, Q => DATA_IN_1_port, QN => n_1259);
   DATAPATH_I_ID_EX_RF_OUT2_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N148,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_2_port, QN 
                           => n_1260);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N245
                           , CK => CLK, Q => DATA_IN_2_port, QN => n_1261);
   DATAPATH_I_ID_EX_RF_OUT2_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N149,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_3_port, QN 
                           => n_1262);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N246
                           , CK => CLK, Q => DATA_IN_3_port, QN => n_1263);
   DATAPATH_I_ID_EX_RF_OUT2_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N150,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_4_port, QN 
                           => n_1264);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N247
                           , CK => CLK, Q => DATA_IN_4_port, QN => n_1265);
   DATAPATH_I_ID_EX_RF_OUT2_reg_5_inst : DFF_X1 port map( D => DATAPATH_I_N151,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_5_port, QN 
                           => n_1266);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_5_inst : DFF_X1 port map( D => DATAPATH_I_N248
                           , CK => CLK, Q => DATA_IN_5_port, QN => n_1267);
   DATAPATH_I_ID_EX_RF_OUT2_reg_6_inst : DFF_X1 port map( D => DATAPATH_I_N152,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_6_port, QN 
                           => n_1268);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_6_inst : DFF_X1 port map( D => DATAPATH_I_N249
                           , CK => CLK, Q => DATA_IN_6_port, QN => n_1269);
   DATAPATH_I_ID_EX_RF_OUT2_reg_7_inst : DFF_X1 port map( D => DATAPATH_I_N153,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_7_port, QN 
                           => n_1270);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_7_inst : DFF_X1 port map( D => DATAPATH_I_N250
                           , CK => CLK, Q => DATA_IN_7_port, QN => n_1271);
   DATAPATH_I_ID_EX_RF_OUT2_reg_8_inst : DFF_X1 port map( D => DATAPATH_I_N154,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_8_port, QN 
                           => n_1272);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_8_inst : DFF_X1 port map( D => DATAPATH_I_N251
                           , CK => CLK, Q => DATA_IN_8_port, QN => n_1273);
   DATAPATH_I_ID_EX_RF_OUT2_reg_9_inst : DFF_X1 port map( D => DATAPATH_I_N155,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_9_port, QN 
                           => n_1274);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_9_inst : DFF_X1 port map( D => DATAPATH_I_N252
                           , CK => CLK, Q => DATA_IN_9_port, QN => n_1275);
   DATAPATH_I_ID_EX_RF_OUT2_reg_10_inst : DFF_X1 port map( D => DATAPATH_I_N156
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_10_port, 
                           QN => n_1276);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_10_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N253, CK => CLK, Q => DATA_IN_10_port, QN
                           => n_1277);
   DATAPATH_I_ID_EX_RF_OUT2_reg_11_inst : DFF_X1 port map( D => DATAPATH_I_N157
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_11_port, 
                           QN => n_1278);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_11_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N254, CK => CLK, Q => DATA_IN_11_port, QN
                           => n_1279);
   DATAPATH_I_ID_EX_RF_OUT2_reg_12_inst : DFF_X1 port map( D => DATAPATH_I_N158
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_12_port, 
                           QN => n_1280);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_12_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N255, CK => CLK, Q => DATA_IN_12_port, QN
                           => n_1281);
   DATAPATH_I_ID_EX_RF_OUT2_reg_13_inst : DFF_X1 port map( D => DATAPATH_I_N159
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_13_port, 
                           QN => n_1282);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_13_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N256, CK => CLK, Q => DATA_IN_13_port, QN
                           => n_1283);
   DATAPATH_I_ID_EX_RF_OUT2_reg_14_inst : DFF_X1 port map( D => DATAPATH_I_N160
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_14_port, 
                           QN => n_1284);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_14_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N257, CK => CLK, Q => DATA_IN_14_port, QN
                           => n_1285);
   DATAPATH_I_ID_EX_RF_OUT2_reg_15_inst : DFF_X1 port map( D => DATAPATH_I_N161
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_15_port, 
                           QN => n_1286);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_15_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N258, CK => CLK, Q => DATA_IN_15_port, QN
                           => n_1287);
   DATAPATH_I_ID_EX_RF_OUT2_reg_16_inst : DFF_X1 port map( D => DATAPATH_I_N162
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_16_port, 
                           QN => n_1288);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_16_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N259, CK => CLK, Q => DATA_IN_16_port, QN
                           => n_1289);
   DATAPATH_I_ID_EX_RF_OUT2_reg_17_inst : DFF_X1 port map( D => DATAPATH_I_N163
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_17_port, 
                           QN => n_1290);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_17_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N260, CK => CLK, Q => DATA_IN_17_port, QN
                           => n_1291);
   DATAPATH_I_ID_EX_RF_OUT2_reg_18_inst : DFF_X1 port map( D => DATAPATH_I_N164
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_18_port, 
                           QN => n_1292);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_18_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N261, CK => CLK, Q => DATA_IN_18_port, QN
                           => n_1293);
   DATAPATH_I_ID_EX_RF_OUT2_reg_19_inst : DFF_X1 port map( D => DATAPATH_I_N165
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_19_port, 
                           QN => n_1294);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_19_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N262, CK => CLK, Q => DATA_IN_19_port, QN
                           => n_1295);
   DATAPATH_I_ID_EX_RF_OUT2_reg_20_inst : DFF_X1 port map( D => DATAPATH_I_N166
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_20_port, 
                           QN => n_1296);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_20_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N263, CK => CLK, Q => DATA_IN_20_port, QN
                           => n_1297);
   DATAPATH_I_ID_EX_RF_OUT2_reg_21_inst : DFF_X1 port map( D => DATAPATH_I_N167
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_21_port, 
                           QN => n_1298);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_21_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N264, CK => CLK, Q => DATA_IN_21_port, QN
                           => n_1299);
   DATAPATH_I_ID_EX_RF_OUT2_reg_22_inst : DFF_X1 port map( D => DATAPATH_I_N168
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_22_port, 
                           QN => n_1300);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_22_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N265, CK => CLK, Q => DATA_IN_22_port, QN
                           => n_1301);
   DATAPATH_I_ID_EX_RF_OUT2_reg_23_inst : DFF_X1 port map( D => DATAPATH_I_N169
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_23_port, 
                           QN => n_1302);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_23_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N266, CK => CLK, Q => DATA_IN_23_port, QN
                           => n_1303);
   DATAPATH_I_ID_EX_RF_OUT2_reg_24_inst : DFF_X1 port map( D => DATAPATH_I_N170
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_24_port, 
                           QN => n_1304);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_24_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N267, CK => CLK, Q => DATA_IN_24_port, QN
                           => n_1305);
   DATAPATH_I_ID_EX_RF_OUT2_reg_25_inst : DFF_X1 port map( D => DATAPATH_I_N171
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_25_port, 
                           QN => n_1306);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_25_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N268, CK => CLK, Q => DATA_IN_25_port, QN
                           => n_1307);
   DATAPATH_I_ID_EX_RF_OUT2_reg_26_inst : DFF_X1 port map( D => DATAPATH_I_N172
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_26_port, 
                           QN => n_1308);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_26_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N269, CK => CLK, Q => DATA_IN_26_port, QN
                           => n_1309);
   DATAPATH_I_ID_EX_RF_OUT2_reg_27_inst : DFF_X1 port map( D => DATAPATH_I_N173
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_27_port, 
                           QN => n_1310);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_27_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N270, CK => CLK, Q => DATA_IN_27_port, QN
                           => n_1311);
   DATAPATH_I_ID_EX_RF_OUT2_reg_28_inst : DFF_X1 port map( D => DATAPATH_I_N174
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_28_port, 
                           QN => n_1312);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_28_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N271, CK => CLK, Q => DATA_IN_28_port, QN
                           => n_1313);
   DATAPATH_I_ID_EX_RF_OUT2_reg_29_inst : DFF_X1 port map( D => DATAPATH_I_N175
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_29_port, 
                           QN => n_1314);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_29_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N272, CK => CLK, Q => DATA_IN_29_port, QN
                           => n_1315);
   DATAPATH_I_ID_EX_RF_OUT2_reg_30_inst : DFF_X1 port map( D => DATAPATH_I_N176
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_30_port, 
                           QN => n_1316);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_30_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N273, CK => CLK, Q => DATA_IN_30_port, QN
                           => n_1317);
   DATAPATH_I_ID_EX_RF_OUT2_reg_31_inst : DFF_X1 port map( D => DATAPATH_I_N177
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_31_port, 
                           QN => n_1318);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_31_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N274, CK => CLK, Q => DATA_IN_31_port, QN
                           => n_1319);
   DATAPATH_I_ID_EX_RF_OUT1_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N114,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_0_port, QN 
                           => n_1320);
   DATAPATH_I_ID_EX_RF_OUT1_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N115,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_1_port, QN 
                           => n_1321);
   DATAPATH_I_ID_EX_RF_OUT1_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N116,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_2_port, QN 
                           => n_1322);
   DATAPATH_I_ID_EX_RF_OUT1_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N117,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_3_port, QN 
                           => n_1323);
   DATAPATH_I_ID_EX_RF_OUT1_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N118,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_4_port, QN 
                           => n_1324);
   DATAPATH_I_ID_EX_RF_OUT1_reg_5_inst : DFF_X1 port map( D => DATAPATH_I_N119,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_5_port, QN 
                           => n_1325);
   DATAPATH_I_ID_EX_RF_OUT1_reg_6_inst : DFF_X1 port map( D => DATAPATH_I_N120,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_6_port, QN 
                           => n_1326);
   DATAPATH_I_ID_EX_RF_OUT1_reg_7_inst : DFF_X1 port map( D => DATAPATH_I_N121,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_7_port, QN 
                           => n_1327);
   DATAPATH_I_ID_EX_RF_OUT1_reg_8_inst : DFF_X1 port map( D => DATAPATH_I_N122,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_8_port, QN 
                           => n_1328);
   DATAPATH_I_ID_EX_RF_OUT1_reg_9_inst : DFF_X1 port map( D => DATAPATH_I_N123,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_9_port, QN 
                           => n_1329);
   DATAPATH_I_ID_EX_RF_OUT1_reg_10_inst : DFF_X1 port map( D => DATAPATH_I_N124
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_10_port, 
                           QN => n_1330);
   DATAPATH_I_ID_EX_RF_OUT1_reg_11_inst : DFF_X1 port map( D => DATAPATH_I_N125
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_11_port, 
                           QN => n_1331);
   DATAPATH_I_ID_EX_RF_OUT1_reg_12_inst : DFF_X1 port map( D => DATAPATH_I_N126
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_12_port, 
                           QN => n_1332);
   DATAPATH_I_ID_EX_RF_OUT1_reg_13_inst : DFF_X1 port map( D => DATAPATH_I_N127
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_13_port, 
                           QN => n_1333);
   DATAPATH_I_ID_EX_RF_OUT1_reg_14_inst : DFF_X1 port map( D => DATAPATH_I_N128
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_14_port, 
                           QN => n_1334);
   DATAPATH_I_ID_EX_RF_OUT1_reg_15_inst : DFF_X1 port map( D => DATAPATH_I_N129
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_15_port, 
                           QN => n_1335);
   DATAPATH_I_ID_EX_RF_OUT1_reg_16_inst : DFF_X1 port map( D => DATAPATH_I_N130
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_16_port, 
                           QN => n_1336);
   DATAPATH_I_ID_EX_RF_OUT1_reg_17_inst : DFF_X1 port map( D => DATAPATH_I_N131
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_17_port, 
                           QN => n_1337);
   DATAPATH_I_ID_EX_RF_OUT1_reg_18_inst : DFF_X1 port map( D => DATAPATH_I_N132
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_18_port, 
                           QN => n_1338);
   DATAPATH_I_ID_EX_RF_OUT1_reg_19_inst : DFF_X1 port map( D => DATAPATH_I_N133
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_19_port, 
                           QN => n_1339);
   DATAPATH_I_ID_EX_RF_OUT1_reg_20_inst : DFF_X1 port map( D => DATAPATH_I_N134
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_20_port, 
                           QN => n_1340);
   DATAPATH_I_ID_EX_RF_OUT1_reg_21_inst : DFF_X1 port map( D => DATAPATH_I_N135
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_21_port, 
                           QN => n_1341);
   DATAPATH_I_ID_EX_RF_OUT1_reg_22_inst : DFF_X1 port map( D => DATAPATH_I_N136
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_22_port, 
                           QN => n_1342);
   DATAPATH_I_ID_EX_RF_OUT1_reg_23_inst : DFF_X1 port map( D => DATAPATH_I_N137
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_23_port, 
                           QN => n_1343);
   DATAPATH_I_ID_EX_RF_OUT1_reg_24_inst : DFF_X1 port map( D => DATAPATH_I_N138
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_24_port, 
                           QN => n_1344);
   DATAPATH_I_ID_EX_RF_OUT1_reg_25_inst : DFF_X1 port map( D => DATAPATH_I_N139
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_25_port, 
                           QN => n_1345);
   DATAPATH_I_ID_EX_RF_OUT1_reg_26_inst : DFF_X1 port map( D => DATAPATH_I_N140
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_26_port, 
                           QN => n_1346);
   DATAPATH_I_ID_EX_RF_OUT1_reg_27_inst : DFF_X1 port map( D => DATAPATH_I_N141
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_27_port, 
                           QN => n_1347);
   DATAPATH_I_ID_EX_RF_OUT1_reg_28_inst : DFF_X1 port map( D => DATAPATH_I_N142
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_28_port, 
                           QN => n_1348);
   DATAPATH_I_ID_EX_RF_OUT1_reg_29_inst : DFF_X1 port map( D => DATAPATH_I_N143
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_29_port, 
                           QN => n_1349);
   DATAPATH_I_ID_EX_RF_OUT1_reg_30_inst : DFF_X1 port map( D => DATAPATH_I_N144
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_30_port, 
                           QN => n_1350);
   DATAPATH_I_ID_EX_RF_OUT1_reg_31_inst : DFF_X1 port map( D => DATAPATH_I_N145
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_31_port, 
                           QN => n_1351);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_N3, GN => n317
                           , Q => IR_0_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_N3, GN => n317
                           , Q => IR_1_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_N3, GN => n317
                           , Q => IR_2_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_N3, GN => n317
                           , Q => IR_3_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_N3, GN => n317
                           , Q => IR_4_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_N3, GN => n317
                           , Q => IR_5_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_N3, GN => n317
                           , Q => IR_6_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_N3, GN => n317
                           , Q => IR_7_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_N3, GN => n317
                           , Q => IR_8_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_N3, GN => n317
                           , Q => IR_9_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_N3, GN => 
                           n317, Q => IR_10_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_N3, GN => 
                           n317, Q => DATAPATH_I_n29);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_N3, GN => 
                           n317, Q => DATAPATH_I_n28);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_N3, GN => 
                           n317, Q => DATAPATH_I_n27);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_N3, GN => 
                           n317, Q => DATAPATH_I_n26);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_N3, GN => 
                           n317, Q => DATAPATH_I_n25);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_N3, GN => 
                           n317, Q => DATAPATH_I_n24);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_N3, GN => 
                           n317, Q => DATAPATH_I_n23);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_N3, GN => 
                           n317, Q => DATAPATH_I_n22);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_N3, GN => 
                           n317, Q => DATAPATH_I_n21);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_N3, GN => 
                           n317, Q => DATAPATH_I_n20);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_N3, GN => 
                           n317, Q => DATAPATH_I_n19);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_N3, GN => 
                           n317, Q => DATAPATH_I_n18);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_N3, GN => 
                           n317, Q => DATAPATH_I_n17);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_N3, GN => 
                           n317, Q => DATAPATH_I_n16);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_N3, GN => 
                           n317, Q => DATAPATH_I_n15);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_N3, GN => 
                           n317, Q => IR_26_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_N3, GN => 
                           n317, Q => IR_27_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_N3, GN => 
                           n317, Q => IR_28_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_N3, GN => 
                           n317, Q => IR_29_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_N3, GN => 
                           n317, Q => IR_30_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_N3, GN => 
                           n317, Q => IR_31_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_0_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_0_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_1_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_1_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_2_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_2_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_3_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_3_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_4_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_4_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_5_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_5_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_6_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_6_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_7_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_7_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_8_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_8_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_9_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_9_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_10_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_10_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_11_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_11_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_12_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_12_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_13_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_13_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_14_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_14_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_15_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_15_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_16_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_16_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_17_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_17_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_18_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_18_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_19_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_19_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_20_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_20_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_21_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_21_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_22_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_22_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_23_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_23_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_24_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_24_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_25_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_25_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_26_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_26_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_27_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_27_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_28_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_28_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_29_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_29_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_30_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_30_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_31_N3, GN => n317, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_31_port);
   DATAPATH_I_LATCH_LMD_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_0_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_0_port);
   DATAPATH_I_LATCH_LMD_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_1_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_1_port);
   DATAPATH_I_LATCH_LMD_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_2_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_2_port);
   DATAPATH_I_LATCH_LMD_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_3_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_3_port);
   DATAPATH_I_LATCH_LMD_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_4_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_4_port);
   DATAPATH_I_LATCH_LMD_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_5_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_5_port);
   DATAPATH_I_LATCH_LMD_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_6_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_6_port);
   DATAPATH_I_LATCH_LMD_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_7_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_7_port);
   DATAPATH_I_LATCH_LMD_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_8_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_8_port);
   DATAPATH_I_LATCH_LMD_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_9_N3, GN => n318, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_9_port);
   DATAPATH_I_LATCH_LMD_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_10_N3, GN => n318, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_10_port);
   DATAPATH_I_LATCH_LMD_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_11_N3, GN => n318, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_11_port);
   DATAPATH_I_LATCH_LMD_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_12_N3, GN => n318, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_12_port);
   DATAPATH_I_LATCH_LMD_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_13_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_13_port);
   DATAPATH_I_LATCH_LMD_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_14_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_14_port);
   DATAPATH_I_LATCH_LMD_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_15_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_15_port);
   DATAPATH_I_LATCH_LMD_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_16_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_16_port);
   DATAPATH_I_LATCH_LMD_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_17_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_17_port);
   DATAPATH_I_LATCH_LMD_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_18_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_18_port);
   DATAPATH_I_LATCH_LMD_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_19_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_19_port);
   DATAPATH_I_LATCH_LMD_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_20_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_20_port);
   DATAPATH_I_LATCH_LMD_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_21_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_21_port);
   DATAPATH_I_LATCH_LMD_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_22_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_22_port);
   DATAPATH_I_LATCH_LMD_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_23_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_23_port);
   DATAPATH_I_LATCH_LMD_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_24_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_24_port);
   DATAPATH_I_LATCH_LMD_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_25_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_25_port);
   DATAPATH_I_LATCH_LMD_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_26_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_26_port);
   DATAPATH_I_LATCH_LMD_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_27_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_27_port);
   DATAPATH_I_LATCH_LMD_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_28_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_28_port);
   DATAPATH_I_LATCH_LMD_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_29_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_29_port);
   DATAPATH_I_LATCH_LMD_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_30_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_30_port);
   DATAPATH_I_LATCH_LMD_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_31_N3, GN => n317, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_31_port);
   DATAPATH_I_LATCH_RF2_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_0_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_0_port);
   DATAPATH_I_LATCH_RF2_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_1_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_1_port);
   DATAPATH_I_LATCH_RF2_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_2_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_2_port);
   DATAPATH_I_LATCH_RF2_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_3_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_3_port);
   DATAPATH_I_LATCH_RF2_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_4_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_4_port);
   DATAPATH_I_LATCH_RF2_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_5_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_5_port);
   DATAPATH_I_LATCH_RF2_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_6_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_6_port);
   DATAPATH_I_LATCH_RF2_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_7_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_7_port);
   DATAPATH_I_LATCH_RF2_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_8_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_8_port);
   DATAPATH_I_LATCH_RF2_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_9_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_9_port);
   DATAPATH_I_LATCH_RF2_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_10_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_10_port);
   DATAPATH_I_LATCH_RF2_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_11_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_11_port);
   DATAPATH_I_LATCH_RF2_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_12_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_12_port);
   DATAPATH_I_LATCH_RF2_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_13_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_13_port);
   DATAPATH_I_LATCH_RF2_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_14_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_14_port);
   DATAPATH_I_LATCH_RF2_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_15_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_15_port);
   DATAPATH_I_LATCH_RF2_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_16_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_16_port);
   DATAPATH_I_LATCH_RF2_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_17_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_17_port);
   DATAPATH_I_LATCH_RF2_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_18_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_18_port);
   DATAPATH_I_LATCH_RF2_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_19_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_19_port);
   DATAPATH_I_LATCH_RF2_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_20_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_20_port);
   DATAPATH_I_LATCH_RF2_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_21_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_21_port);
   DATAPATH_I_LATCH_RF2_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_22_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_22_port);
   DATAPATH_I_LATCH_RF2_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_23_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_23_port);
   DATAPATH_I_LATCH_RF2_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_24_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_24_port);
   DATAPATH_I_LATCH_RF2_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_25_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_25_port);
   DATAPATH_I_LATCH_RF2_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_26_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_26_port);
   DATAPATH_I_LATCH_RF2_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_27_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_27_port);
   DATAPATH_I_LATCH_RF2_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_28_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_28_port);
   DATAPATH_I_LATCH_RF2_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_29_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_29_port);
   DATAPATH_I_LATCH_RF2_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_30_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_30_port);
   DATAPATH_I_LATCH_RF2_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_31_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_31_port);
   DATAPATH_I_LATCH_RF1_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_0_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_0_port);
   DATAPATH_I_LATCH_RF1_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_1_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_1_port);
   DATAPATH_I_LATCH_RF1_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_2_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_2_port);
   DATAPATH_I_LATCH_RF1_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_3_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_3_port);
   DATAPATH_I_LATCH_RF1_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_4_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_4_port);
   DATAPATH_I_LATCH_RF1_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_5_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_5_port);
   DATAPATH_I_LATCH_RF1_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_6_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_6_port);
   DATAPATH_I_LATCH_RF1_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_7_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_7_port);
   DATAPATH_I_LATCH_RF1_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_8_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_8_port);
   DATAPATH_I_LATCH_RF1_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_9_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_9_port);
   DATAPATH_I_LATCH_RF1_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_10_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_10_port);
   DATAPATH_I_LATCH_RF1_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_11_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_11_port);
   DATAPATH_I_LATCH_RF1_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_12_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_12_port);
   DATAPATH_I_LATCH_RF1_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_13_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_13_port);
   DATAPATH_I_LATCH_RF1_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_14_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_14_port);
   DATAPATH_I_LATCH_RF1_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_15_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_15_port);
   DATAPATH_I_LATCH_RF1_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_16_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_16_port);
   DATAPATH_I_LATCH_RF1_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_17_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_17_port);
   DATAPATH_I_LATCH_RF1_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_18_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_18_port);
   DATAPATH_I_LATCH_RF1_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_19_N3, GN => n317, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_19_port);
   DATAPATH_I_LATCH_RF1_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_20_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_20_port);
   DATAPATH_I_LATCH_RF1_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_21_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_21_port);
   DATAPATH_I_LATCH_RF1_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_22_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_22_port);
   DATAPATH_I_LATCH_RF1_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_23_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_23_port);
   DATAPATH_I_LATCH_RF1_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_24_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_24_port);
   DATAPATH_I_LATCH_RF1_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_25_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_25_port);
   DATAPATH_I_LATCH_RF1_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_26_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_26_port);
   DATAPATH_I_LATCH_RF1_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_27_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_27_port);
   DATAPATH_I_LATCH_RF1_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_28_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_28_port);
   DATAPATH_I_LATCH_RF1_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_29_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_29_port);
   DATAPATH_I_LATCH_RF1_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_30_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_30_port);
   DATAPATH_I_LATCH_RF1_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_31_N3, GN => n318, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_31_port);
   CU_I_aluOpcode2_reg_0_inst : DFFR_X1 port map( D => CU_I_aluOpcode1_0_port, 
                           CK => CLK, RN => n317, Q => CU_I_aluOpcode2_0_port, 
                           QN => n_1352);
   CU_I_aluOpcode3_reg_0_inst : DFFR_X1 port map( D => CU_I_aluOpcode2_0_port, 
                           CK => CLK, RN => n317, Q => ALU_OPCODE_i_6_port, QN 
                           => n_1353);
   CU_I_aluOpcode2_reg_3_inst : DFFR_X1 port map( D => CU_I_aluOpcode1_3_port, 
                           CK => CLK, RN => n317, Q => CU_I_aluOpcode2_3_port, 
                           QN => n_1354);
   CU_I_aluOpcode3_reg_3_inst : DFFR_X1 port map( D => CU_I_aluOpcode2_3_port, 
                           CK => CLK, RN => n317, Q => ALU_OPCODE_i_3_port, QN 
                           => n_1355);
   CU_I_aluOpcode2_reg_4_inst : DFFR_X1 port map( D => CU_I_aluOpcode1_4_port, 
                           CK => CLK, RN => n317, Q => CU_I_aluOpcode2_4_port, 
                           QN => n_1356);
   CU_I_aluOpcode3_reg_4_inst : DFFR_X1 port map( D => CU_I_aluOpcode2_4_port, 
                           CK => CLK, RN => n317, Q => ALU_OPCODE_i_2_port, QN 
                           => n_1357);
   CU_I_aluOpcode2_reg_2_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_2_port, 
                           CK => CLK, SN => n317, Q => CU_I_aluOpcode2_2_port, 
                           QN => n_1358);
   CU_I_aluOpcode3_reg_2_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_2_port, 
                           CK => CLK, SN => n317, Q => ALU_OPCODE_i_4_port, QN 
                           => n_1359);
   CU_I_aluOpcode2_reg_1_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_1_port, 
                           CK => CLK, SN => n317, Q => CU_I_aluOpcode2_1_port, 
                           QN => n_1360);
   CU_I_aluOpcode3_reg_1_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_1_port, 
                           CK => CLK, SN => n317, Q => ALU_OPCODE_i_5_port, QN 
                           => n_1361);
   CU_I_aluOpcode2_reg_5_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_5_port, 
                           CK => CLK, SN => n317, Q => CU_I_aluOpcode2_5_port, 
                           QN => n_1362);
   CU_I_aluOpcode3_reg_5_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_5_port, 
                           CK => CLK, SN => n317, Q => ALU_OPCODE_i_1_port, QN 
                           => n_1363);
   CU_I_aluOpcode2_reg_6_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_6_port, 
                           CK => CLK, SN => n317, Q => CU_I_aluOpcode2_6_port, 
                           QN => n_1364);
   CU_I_aluOpcode3_reg_6_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_6_port, 
                           CK => CLK, SN => n317, Q => ALU_OPCODE_i_0_port, QN 
                           => n_1365);
   DATAPATH_I_ID_EX_RD_reg_3_inst : DFF_X2 port map( D => DATAPATH_I_N112, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_3_port, QN => 
                           n_1366);
   DATAPATH_I_ID_EX_RD_reg_1_inst : DFF_X2 port map( D => DATAPATH_I_N110, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_1_port, QN => 
                           n_1367);
   DATAPATH_I_ID_EX_RD_reg_4_inst : DFFS_X2 port map( D => DATAPATH_I_N113, CK 
                           => CLK, SN => n475, Q => DATAPATH_I_ID_EX_RD_4_port,
                           QN => n_1368);
   DATAPATH_I_ID_EX_RD_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N111, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_2_port, QN => 
                           n_1369);
   DATAPATH_I_ID_EX_RD_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N109, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_0_port, QN => 
                           n_1370);
   U751 : INV_X2 port map( A => RST, ZN => n322);
   U752 : INV_X1 port map( A => RST, ZN => n321);
   U753 : INV_X8 port map( A => n321, ZN => n318);
   U754 : INV_X8 port map( A => n321, ZN => n319);
   U755 : INV_X8 port map( A => n322, ZN => n317);
   U756 : INV_X1 port map( A => n321, ZN => n320);
   U757 : AND2_X1 port map( A1 => n374, A2 => n375, ZN => n323);
   U758 : AND2_X1 port map( A1 => n375, A2 => n374, ZN => n385);
   U759 : AND2_X1 port map( A1 => n485, A2 => n486, ZN => n324);
   U760 : AND2_X2 port map( A1 => n326, A2 => n367, ZN => n325);
   U761 : AND2_X1 port map( A1 => n326, A2 => n367, ZN => n386);
   U762 : AND2_X1 port map( A1 => n324, A2 => n336, ZN => n326);
   U763 : NAND2_X1 port map( A1 => n328, A2 => n369, ZN => n327);
   U764 : BUF_X1 port map( A => n370, Z => n328);
   U765 : BUF_X1 port map( A => n374, Z => n329);
   U766 : AND2_X1 port map( A1 => n388, A2 => n327, ZN => n389);
   U767 : AND2_X1 port map( A1 => n382, A2 => n387, ZN => n383);
   U768 : AND2_X1 port map( A1 => n379, A2 => n327, ZN => n380);
   U769 : AND2_X1 port map( A1 => n376, A2 => n387, ZN => n377);
   U770 : OAI21_X1 port map( B1 => n337, B2 => n326, A => n366, ZN => n330);
   U771 : OAI21_X1 port map( B1 => n337, B2 => n368, A => n366, ZN => n375);
   U772 : NOR2_X1 port map( A1 => n479, A2 => n338, ZN => n331);
   U773 : NOR2_X1 port map( A1 => n477, A2 => n338, ZN => n332);
   U774 : NOR2_X1 port map( A1 => n476, A2 => n338, ZN => n333);
   U775 : NOR2_X1 port map( A1 => n478, A2 => n338, ZN => n334);
   U776 : NOR2_X1 port map( A1 => n480, A2 => n338, ZN => n335);
   n475 <= '1';
   U778 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_0_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_N3);
   U779 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_1_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_N3);
   U780 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_2_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_N3);
   U781 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_3_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_N3);
   U782 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_4_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_N3);
   U783 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_5_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_N3);
   U784 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_6_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_N3);
   U785 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_7_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_N3);
   U786 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_8_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_N3);
   U787 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_9_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_N3);
   U788 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_10_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_N3);
   U789 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_11_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_N3);
   U790 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_12_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_N3);
   U791 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_13_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_N3);
   U792 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_14_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_N3);
   U793 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_15_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_N3);
   U794 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_16_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_N3);
   U795 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_17_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_N3);
   U796 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_18_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_N3);
   U797 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_19_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_N3);
   U798 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_20_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_N3);
   U799 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_21_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_N3);
   U800 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_22_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_N3);
   U801 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_23_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_N3);
   U802 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_24_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_N3);
   U803 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_25_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_N3);
   U804 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_26_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_N3);
   U805 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_27_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_N3);
   U806 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_28_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_N3);
   U807 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_29_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_N3);
   U808 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_30_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_N3);
   U809 : AND2_X1 port map( A1 => n319, A2 => IR_BUS_31_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_N3);
   U810 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_0_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_0_N3);
   U811 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_1_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_1_N3);
   U812 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_2_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_2_N3);
   U813 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_3_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_3_N3);
   U814 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_4_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_4_N3);
   U815 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_5_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_5_N3);
   U816 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_6_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_6_N3);
   U817 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_7_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_7_N3);
   U818 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_8_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_8_N3);
   U819 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_9_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_9_N3);
   U820 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_10_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_10_N3);
   U821 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_11_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_11_N3);
   U822 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_12_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_12_N3);
   U823 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_13_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_13_N3);
   U824 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_14_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_14_N3);
   U825 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_15_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_15_N3);
   U826 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_16_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_16_N3);
   U827 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_17_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_17_N3);
   U828 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_18_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_18_N3);
   U829 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_19_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_19_N3);
   U830 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_20_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_20_N3);
   U831 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_21_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_21_N3);
   U832 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_22_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_22_N3);
   U833 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_23_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_23_N3);
   U834 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_24_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_24_N3);
   U835 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_25_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_25_N3);
   U836 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_26_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_26_N3);
   U837 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_27_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_27_N3);
   U838 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_28_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_28_N3);
   U839 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_29_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_29_N3);
   U840 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ALU_OUTPUT_31_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_31_N3);
   U841 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_0_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_0_N3);
   U842 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_1_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_1_N3);
   U843 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_2_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_2_N3);
   U844 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_3_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_3_N3);
   U845 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_4_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_4_N3);
   U846 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_5_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_5_N3);
   U847 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_6_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_6_N3);
   U848 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_7_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_7_N3);
   U849 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_8_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_8_N3);
   U850 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_9_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_9_N3);
   U851 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_10_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_10_N3);
   U852 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_11_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_11_N3);
   U853 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_12_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_12_N3);
   U854 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_13_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_13_N3);
   U855 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_14_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_14_N3);
   U856 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_15_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_15_N3);
   U857 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_16_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_16_N3);
   U858 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_17_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_17_N3);
   U859 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_18_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_18_N3);
   U860 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_19_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_19_N3);
   U861 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_20_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_20_N3);
   U862 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_21_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_21_N3);
   U863 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_22_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_22_N3);
   U864 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_23_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_23_N3);
   U865 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_24_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_24_N3);
   U866 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_25_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_25_N3);
   U867 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_26_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_26_N3);
   U868 : AND2_X1 port map( A1 => n320, A2 => DATA_OUT_27_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_27_N3);
   U869 : AND2_X1 port map( A1 => n319, A2 => DATA_OUT_28_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_28_N3);
   U870 : AND2_X1 port map( A1 => n320, A2 => DATA_OUT_29_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_29_N3);
   U871 : AND2_X1 port map( A1 => n320, A2 => DATA_OUT_30_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_30_N3);
   U872 : AND2_X1 port map( A1 => n320, A2 => DATA_OUT_31_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_31_N3);
   U873 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_0_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_0_N3);
   U874 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_1_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_1_N3);
   U875 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_2_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_2_N3);
   U876 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_3_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_3_N3);
   U877 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_4_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_4_N3);
   U878 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_5_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_5_N3);
   U879 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_6_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_6_N3);
   U880 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_7_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_7_N3);
   U881 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_8_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_8_N3);
   U882 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_9_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_9_N3);
   U883 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_10_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_10_N3);
   U884 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_11_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_11_N3);
   U885 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_12_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_12_N3);
   U886 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_13_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_13_N3);
   U887 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_14_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_14_N3);
   U888 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_15_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_15_N3);
   U889 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_16_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_16_N3);
   U890 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_17_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_17_N3);
   U891 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_18_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_18_N3);
   U892 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_19_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_19_N3);
   U893 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_20_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_20_N3);
   U894 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_21_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_21_N3);
   U895 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_22_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_22_N3);
   U896 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_23_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_23_N3);
   U897 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_24_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_24_N3);
   U898 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_25_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_25_N3);
   U899 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_26_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_26_N3);
   U900 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_27_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_27_N3);
   U901 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_ALU_OUTPUT_30_port, ZN
                           => DATAPATH_I_LATCH_ALUOUT_LDI_30_N3);
   U902 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_29_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_29_N3);
   U903 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_30_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_30_N3);
   U904 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_31_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_31_N3);
   U905 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT1_0_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_0_N3);
   U906 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT1_1_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_1_N3);
   U907 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT2_28_port, ZN =>
                           DATAPATH_I_LATCH_RF2_LDI_28_N3);
   U908 : AND2_X1 port map( A1 => n482, A2 => n481, ZN => n336);
   U909 : AND2_X1 port map( A1 => n486, A2 => n485, ZN => n339);
   U910 : AND2_X1 port map( A1 => n324, A2 => n336, ZN => n368);
   U911 : AND4_X2 port map( A1 => DATAPATH_I_IF_ID_IR_29_port, A2 => 
                           DATAPATH_I_IF_ID_IR_31_port, A3 => 
                           DATAPATH_I_IF_ID_IR_27_port, A4 => 
                           DATAPATH_I_IF_ID_IR_26_port, ZN => n337);
   U912 : AND2_X1 port map( A1 => n483, A2 => n484, ZN => n366);
   U913 : CLKBUF_X1 port map( A => n330, Z => n338);
   U914 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT1_2_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_2_N3);
   U915 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT1_3_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_3_N3);
   U916 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT1_4_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_4_N3);
   U917 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_RF_OUT1_5_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_5_N3);
   U918 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_6_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_6_N3);
   U919 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_7_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_7_N3);
   U920 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_8_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_8_N3);
   U921 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_9_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_9_N3);
   U922 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_10_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_10_N3);
   U923 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_11_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_11_N3);
   U924 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_12_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_12_N3);
   U925 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_13_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_13_N3);
   U926 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_14_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_14_N3);
   U927 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_15_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_15_N3);
   U928 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_16_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_16_N3);
   U929 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_17_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_17_N3);
   U930 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_18_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_18_N3);
   U931 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_19_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_19_N3);
   U932 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_28_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_28_N3);
   U933 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_20_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_20_N3);
   U934 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_27_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_27_N3);
   U935 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_21_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_21_N3);
   U936 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_30_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_30_N3);
   U937 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_22_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_22_N3);
   U938 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_31_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_31_N3);
   U939 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_23_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_23_N3);
   U940 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_29_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_29_N3);
   U941 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_24_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_24_N3);
   U942 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_25_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_25_N3);
   U943 : INV_X1 port map( A => IR_28_port, ZN => n442);
   U944 : NOR2_X1 port map( A1 => n322, A2 => n442, ZN => DATAPATH_I_N62);
   U945 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_RF_OUT1_26_port, ZN =>
                           DATAPATH_I_LATCH_RF1_LDI_26_N3);
   U946 : NOR2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_28_port, A2 => n482, ZN 
                           => n340);
   U947 : AND2_X1 port map( A1 => n340, A2 => n339, ZN => n370);
   U948 : CLKBUF_X1 port map( A => n328, Z => n342);
   U949 : INV_X1 port map( A => DATAPATH_I_IF_ID_IR_30_port, ZN => n341);
   U950 : NAND2_X1 port map( A1 => n342, A2 => n341, ZN => n343);
   U951 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_25_port, A2 => n343, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_4_port);
   U952 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_23_port, A2 => n343, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_2_port);
   U953 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_22_port, A2 => n343, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_1_port);
   U954 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_21_port, A2 => n343, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_0_port);
   U955 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_EX_MEM_RD_3_port, ZN 
                           => DATAPATH_I_N413);
   U956 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RD_0_port, ZN =>
                           DATAPATH_I_N308);
   U957 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RD_1_port, ZN =>
                           DATAPATH_I_N309);
   U958 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_EX_MEM_RD_1_port, ZN 
                           => DATAPATH_I_N411);
   U959 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RD_2_port, ZN =>
                           DATAPATH_I_N310);
   U960 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_EX_MEM_RD_0_port, ZN 
                           => DATAPATH_I_N410);
   U961 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RD_4_port, ZN =>
                           DATAPATH_I_N312);
   U962 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RD_3_port, ZN =>
                           DATAPATH_I_N311);
   U963 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_EX_MEM_RD_2_port, ZN 
                           => DATAPATH_I_N412);
   U964 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_EX_MEM_RD_4_port, ZN 
                           => DATAPATH_I_N414);
   U965 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_31_port, ZN => 
                           DATAPATH_I_N177);
   U966 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_8_port, ZN => 
                           DATAPATH_I_N122);
   U967 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_3_port, ZN => 
                           DATAPATH_I_N117);
   U968 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_27_port, ZN => 
                           DATAPATH_I_N173);
   U969 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_12_port, ZN => 
                           DATAPATH_I_N126);
   U970 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_6_port, ZN => 
                           DATAPATH_I_N120);
   U971 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_28_port, ZN => 
                           DATAPATH_I_N174);
   U972 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_2_port, ZN => 
                           DATAPATH_I_N116);
   U973 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_29_port, ZN => 
                           DATAPATH_I_N175);
   U974 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_14_port, ZN => 
                           DATAPATH_I_N128);
   U975 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_30_port, ZN => 
                           DATAPATH_I_N176);
   U976 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_13_port, ZN => 
                           DATAPATH_I_N127);
   U977 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_7_port, ZN => 
                           DATAPATH_I_N121);
   U978 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_24_port, ZN => 
                           DATAPATH_I_N170);
   U979 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_26_port, ZN => 
                           DATAPATH_I_N172);
   U980 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_4_port, ZN => 
                           DATAPATH_I_N118);
   U981 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_15_port, ZN => 
                           DATAPATH_I_N129);
   U982 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_9_port, ZN => 
                           DATAPATH_I_N123);
   U983 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_23_port, ZN => 
                           DATAPATH_I_N169);
   U984 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_5_port, ZN => 
                           DATAPATH_I_N119);
   U985 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_16_port, ZN => 
                           DATAPATH_I_N130);
   U986 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_10_port, ZN => 
                           DATAPATH_I_N124);
   U987 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_0_port, ZN => 
                           DATAPATH_I_N114);
   U988 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_22_port, ZN => 
                           DATAPATH_I_N168);
   U989 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_17_port, ZN => 
                           DATAPATH_I_N131);
   U990 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_11_port, ZN => 
                           DATAPATH_I_N125);
   U991 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_1_port, ZN => 
                           DATAPATH_I_N115);
   U992 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_25_port, ZN => 
                           DATAPATH_I_N171);
   U993 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_18_port, ZN => 
                           DATAPATH_I_N132);
   U994 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_21_port, ZN => 
                           DATAPATH_I_N167);
   U995 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_19_port, ZN => 
                           DATAPATH_I_N133);
   U996 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_20_port, ZN => 
                           DATAPATH_I_N134);
   U997 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_21_port, ZN => 
                           DATAPATH_I_N135);
   U998 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_22_port, ZN => 
                           DATAPATH_I_N136);
   U999 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_23_port, ZN => 
                           DATAPATH_I_N137);
   U1000 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_24_port, ZN => 
                           DATAPATH_I_N138);
   U1001 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_25_port, ZN => 
                           DATAPATH_I_N139);
   U1002 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_26_port, ZN => 
                           DATAPATH_I_N140);
   U1003 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_27_port, ZN => 
                           DATAPATH_I_N141);
   U1004 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_28_port, ZN => 
                           DATAPATH_I_N142);
   U1005 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_29_port, ZN => 
                           DATAPATH_I_N143);
   U1006 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_30_port, ZN => 
                           DATAPATH_I_N144);
   U1007 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_31_port, ZN => 
                           DATAPATH_I_N145);
   U1008 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_20_port, ZN => 
                           DATAPATH_I_N166);
   U1009 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n27, ZN => 
                           DATAPATH_I_N47);
   U1010 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n26, ZN => 
                           DATAPATH_I_N48);
   U1011 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n25, ZN => 
                           DATAPATH_I_N49);
   U1012 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n24, ZN => 
                           DATAPATH_I_N50);
   U1013 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n23, ZN => 
                           DATAPATH_I_N51);
   U1014 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n22, ZN => 
                           DATAPATH_I_N52);
   U1015 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n21, ZN => 
                           DATAPATH_I_N53);
   U1016 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n20, ZN => 
                           DATAPATH_I_N54);
   U1017 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n19, ZN => 
                           DATAPATH_I_N55);
   U1018 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n18, ZN => 
                           DATAPATH_I_N56);
   U1019 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n17, ZN => 
                           DATAPATH_I_N57);
   U1020 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n16, ZN => 
                           DATAPATH_I_N58);
   U1021 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n15, ZN => 
                           DATAPATH_I_N59);
   U1022 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_0_port, ZN => 
                           DATAPATH_I_N275);
   U1023 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_1_port, ZN => 
                           DATAPATH_I_N276);
   U1024 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_2_port, ZN => 
                           DATAPATH_I_N277);
   U1025 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_3_port, ZN => 
                           DATAPATH_I_N278);
   U1026 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_4_port, ZN => 
                           DATAPATH_I_N279);
   U1027 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_5_port, ZN => 
                           DATAPATH_I_N280);
   U1028 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_6_port, ZN => 
                           DATAPATH_I_N281);
   U1029 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_7_port, ZN => 
                           DATAPATH_I_N282);
   U1030 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_8_port, ZN => 
                           DATAPATH_I_N283);
   U1031 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_9_port, ZN => 
                           DATAPATH_I_N284);
   U1032 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_10_port, ZN => 
                           DATAPATH_I_N285);
   U1033 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_11_port, ZN => 
                           DATAPATH_I_N286);
   U1034 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_12_port, ZN => 
                           DATAPATH_I_N287);
   U1035 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_13_port, ZN => 
                           DATAPATH_I_N288);
   U1036 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_14_port, ZN => 
                           DATAPATH_I_N289);
   U1037 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_15_port, ZN => 
                           DATAPATH_I_N290);
   U1038 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_16_port, ZN => 
                           DATAPATH_I_N291);
   U1039 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_17_port, ZN => 
                           DATAPATH_I_N292);
   U1040 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_18_port, ZN => 
                           DATAPATH_I_N293);
   U1041 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_19_port, ZN => 
                           DATAPATH_I_N294);
   U1042 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_20_port, ZN => 
                           DATAPATH_I_N295);
   U1043 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_21_port, ZN => 
                           DATAPATH_I_N296);
   U1044 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_22_port, ZN => 
                           DATAPATH_I_N297);
   U1045 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_23_port, ZN => 
                           DATAPATH_I_N298);
   U1046 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_24_port, ZN => 
                           DATAPATH_I_N299);
   U1047 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_25_port, ZN => 
                           DATAPATH_I_N300);
   U1048 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_26_port, ZN => 
                           DATAPATH_I_N301);
   U1049 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_27_port, ZN => 
                           DATAPATH_I_N302);
   U1050 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_28_port, ZN => 
                           DATAPATH_I_N303);
   U1051 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_29_port, ZN => 
                           DATAPATH_I_N304);
   U1052 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_30_port, ZN => 
                           DATAPATH_I_N305);
   U1053 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_31_port, ZN => 
                           DATAPATH_I_N306);
   U1054 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_0_port, ZN => 
                           DATAPATH_I_N378);
   U1055 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n28, ZN => 
                           DATAPATH_I_N46);
   U1056 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_1_port, ZN => 
                           DATAPATH_I_N379);
   U1057 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_2_port, ZN => 
                           DATAPATH_I_N380);
   U1058 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_3_port, ZN => 
                           DATAPATH_I_N381);
   U1059 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_4_port, ZN => 
                           DATAPATH_I_N382);
   U1060 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_5_port, ZN => 
                           DATAPATH_I_N383);
   U1061 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_6_port, ZN => 
                           DATAPATH_I_N384);
   U1062 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_7_port, ZN => 
                           DATAPATH_I_N385);
   U1063 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_8_port, ZN => 
                           DATAPATH_I_N386);
   U1064 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_9_port, ZN => 
                           DATAPATH_I_N387);
   U1065 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_10_port, ZN => 
                           DATAPATH_I_N388);
   U1066 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_11_port, ZN => 
                           DATAPATH_I_N389);
   U1067 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_n29, ZN => 
                           DATAPATH_I_N45);
   U1068 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_13_port, ZN => 
                           DATAPATH_I_N391);
   U1069 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_14_port, ZN => 
                           DATAPATH_I_N392);
   U1070 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_15_port, ZN => 
                           DATAPATH_I_N393);
   U1071 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_16_port, ZN => 
                           DATAPATH_I_N394);
   U1072 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_17_port, ZN => 
                           DATAPATH_I_N395);
   U1073 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_18_port, ZN => 
                           DATAPATH_I_N396);
   U1074 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_19_port, ZN => 
                           DATAPATH_I_N397);
   U1075 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_20_port, ZN => 
                           DATAPATH_I_N398);
   U1076 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_21_port, ZN => 
                           DATAPATH_I_N399);
   U1077 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_22_port, ZN => 
                           DATAPATH_I_N400);
   U1078 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_23_port, ZN => 
                           DATAPATH_I_N401);
   U1079 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_24_port, ZN => 
                           DATAPATH_I_N402);
   U1080 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_25_port, ZN => 
                           DATAPATH_I_N403);
   U1081 : AND2_X1 port map( A1 => n318, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_26_port, ZN => 
                           DATAPATH_I_N404);
   U1082 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_27_port, ZN => 
                           DATAPATH_I_N405);
   U1083 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_28_port, ZN => 
                           DATAPATH_I_N406);
   U1084 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_29_port, ZN => 
                           DATAPATH_I_N407);
   U1085 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_30_port, ZN => 
                           DATAPATH_I_N408);
   U1086 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_31_port, ZN => 
                           DATAPATH_I_N409);
   U1087 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_0_port, ZN => 
                           DATAPATH_I_N146);
   U1088 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_1_port, ZN => 
                           DATAPATH_I_N147);
   U1089 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_2_port, ZN => 
                           DATAPATH_I_N148);
   U1090 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_3_port, ZN => 
                           DATAPATH_I_N149);
   U1091 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_4_port, ZN => 
                           DATAPATH_I_N150);
   U1092 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_5_port, ZN => 
                           DATAPATH_I_N151);
   U1093 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_6_port, ZN => 
                           DATAPATH_I_N152);
   U1094 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_7_port, ZN => 
                           DATAPATH_I_N153);
   U1095 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_8_port, ZN => 
                           DATAPATH_I_N154);
   U1096 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_9_port, ZN => 
                           DATAPATH_I_N155);
   U1097 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_10_port, ZN => 
                           DATAPATH_I_N156);
   U1098 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_11_port, ZN => 
                           DATAPATH_I_N157);
   U1099 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_12_port, ZN => 
                           DATAPATH_I_N158);
   U1100 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_13_port, ZN => 
                           DATAPATH_I_N159);
   U1101 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_14_port, ZN => 
                           DATAPATH_I_N160);
   U1102 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_15_port, ZN => 
                           DATAPATH_I_N161);
   U1103 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_16_port, ZN => 
                           DATAPATH_I_N162);
   U1104 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_17_port, ZN => 
                           DATAPATH_I_N163);
   U1105 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_18_port, ZN => 
                           DATAPATH_I_N164);
   U1106 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_19_port, ZN => 
                           DATAPATH_I_N165);
   U1107 : AND2_X1 port map( A1 => n319, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_12_port, ZN => 
                           DATAPATH_I_N390);
   U1108 : AND2_X1 port map( A1 => n319, A2 => IR_30_port, ZN => DATAPATH_I_N64
                           );
   U1109 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_24_port
                           , ZN => DATAPATH_I_N267);
   U1110 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_9_port,
                           ZN => DATAPATH_I_N252);
   U1111 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_12_port
                           , ZN => DATAPATH_I_N255);
   U1112 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_7_port,
                           ZN => DATAPATH_I_N250);
   U1113 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_13_port
                           , ZN => DATAPATH_I_N256);
   U1114 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_5_port,
                           ZN => DATAPATH_I_N248);
   U1115 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_15_port
                           , ZN => DATAPATH_I_N258);
   U1116 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_0_port,
                           ZN => DATAPATH_I_N243);
   U1117 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_1_port,
                           ZN => DATAPATH_I_N244);
   U1118 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_11_port
                           , ZN => DATAPATH_I_N254);
   U1119 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_4_port,
                           ZN => DATAPATH_I_N247);
   U1120 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_31_port
                           , ZN => DATAPATH_I_N274);
   U1121 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_3_port,
                           ZN => DATAPATH_I_N246);
   U1122 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_14_port
                           , ZN => DATAPATH_I_N257);
   U1123 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_30_port
                           , ZN => DATAPATH_I_N273);
   U1124 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_2_port,
                           ZN => DATAPATH_I_N245);
   U1125 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_28_port
                           , ZN => DATAPATH_I_N271);
   U1126 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_27_port
                           , ZN => DATAPATH_I_N270);
   U1127 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_17_port
                           , ZN => DATAPATH_I_N260);
   U1128 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_8_port,
                           ZN => DATAPATH_I_N251);
   U1129 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_18_port
                           , ZN => DATAPATH_I_N261);
   U1130 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_6_port,
                           ZN => DATAPATH_I_N249);
   U1131 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_19_port
                           , ZN => DATAPATH_I_N262);
   U1132 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_26_port
                           , ZN => DATAPATH_I_N269);
   U1133 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_20_port
                           , ZN => DATAPATH_I_N263);
   U1134 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_16_port
                           , ZN => DATAPATH_I_N259);
   U1135 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_21_port
                           , ZN => DATAPATH_I_N264);
   U1136 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_25_port
                           , ZN => DATAPATH_I_N268);
   U1137 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_22_port
                           , ZN => DATAPATH_I_N265);
   U1138 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_10_port
                           , ZN => DATAPATH_I_N253);
   U1139 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_23_port
                           , ZN => DATAPATH_I_N266);
   U1140 : AND2_X1 port map( A1 => n319, A2 => DATAPATH_I_ID_EX_RF_OUT2_29_port
                           , ZN => DATAPATH_I_N272);
   U1141 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_24_port, A2 => n343, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_3_port);
   U1142 : INV_X1 port map( A => IR_26_port, ZN => n422);
   U1143 : NOR2_X1 port map( A1 => n322, A2 => n422, ZN => DATAPATH_I_N60);
   U1144 : INV_X1 port map( A => IR_5_port, ZN => n419);
   U1145 : OR4_X1 port map( A1 => IR_6_port, A2 => IR_9_port, A3 => IR_7_port, 
                           A4 => IR_8_port, ZN => n344);
   U1146 : NOR2_X1 port map( A1 => IR_10_port, A2 => n344, ZN => n345);
   U1147 : INV_X1 port map( A => IR_4_port, ZN => n347);
   U1148 : NAND2_X1 port map( A1 => n345, A2 => n347, ZN => n349);
   U1149 : NOR2_X1 port map( A1 => n419, A2 => n349, ZN => n352);
   U1150 : INV_X1 port map( A => n352, ZN => n348);
   U1151 : NOR2_X1 port map( A1 => IR_1_port, A2 => n348, ZN => n402);
   U1152 : INV_X1 port map( A => IR_1_port, ZN => n405);
   U1153 : INV_X1 port map( A => IR_2_port, ZN => n350);
   U1154 : NAND2_X1 port map( A1 => n345, A2 => IR_3_port, ZN => n346);
   U1155 : NOR2_X1 port map( A1 => n347, A2 => n346, ZN => n420);
   U1156 : NAND2_X1 port map( A1 => IR_5_port, A2 => n420, ZN => n410);
   U1157 : AOI221_X1 port map( B1 => IR_1_port, B2 => IR_2_port, C1 => n405, C2
                           => n350, A => n410, ZN => n418);
   U1158 : AOI21_X1 port map( B1 => IR_3_port, B2 => n402, A => n418, ZN => 
                           n440);
   U1159 : NOR2_X1 port map( A1 => IR_31_port, A2 => IR_30_port, ZN => n397);
   U1160 : INV_X1 port map( A => IR_29_port, ZN => n392);
   U1161 : NAND2_X1 port map( A1 => n397, A2 => n392, ZN => n443);
   U1162 : NOR4_X1 port map( A1 => IR_28_port, A2 => IR_27_port, A3 => 
                           IR_26_port, A4 => n443, ZN => n474);
   U1163 : INV_X1 port map( A => IR_3_port, ZN => n401);
   U1164 : NAND2_X1 port map( A1 => n350, A2 => IR_1_port, ZN => n411);
   U1165 : NOR2_X1 port map( A1 => n411, A2 => n348, ZN => n406);
   U1166 : OR4_X1 port map( A1 => IR_5_port, A2 => IR_3_port, A3 => n350, A4 =>
                           n349, ZN => n407);
   U1167 : NOR2_X1 port map( A1 => n405, A2 => n407, ZN => n415);
   U1168 : AOI21_X1 port map( B1 => n401, B2 => n406, A => n415, ZN => n351);
   U1169 : INV_X1 port map( A => n351, ZN => n439);
   U1170 : INV_X1 port map( A => n402, ZN => n453);
   U1171 : NOR2_X1 port map( A1 => IR_2_port, A2 => n453, ZN => n417);
   U1172 : INV_X1 port map( A => IR_0_port, ZN => n456);
   U1173 : OAI211_X1 port map( C1 => n439, C2 => n417, A => n401, B => n456, ZN
                           => n354);
   U1174 : NAND3_X1 port map( A1 => IR_3_port, A2 => n406, A3 => IR_0_port, ZN 
                           => n353);
   U1175 : NAND4_X1 port map( A1 => IR_2_port, A2 => n352, A3 => n401, A4 => 
                           n456, ZN => n404);
   U1176 : AND4_X1 port map( A1 => n474, A2 => n354, A3 => n353, A4 => n404, ZN
                           => n364);
   U1177 : NAND2_X1 port map( A1 => IR_29_port, A2 => n397, ZN => n441);
   U1178 : INV_X1 port map( A => n441, ZN => n465);
   U1179 : INV_X1 port map( A => DATAPATH_I_N62, ZN => n433);
   U1180 : NOR4_X1 port map( A1 => IR_27_port, A2 => n443, A3 => n422, A4 => 
                           n433, ZN => n362);
   U1181 : INV_X1 port map( A => IR_27_port, ZN => n391);
   U1182 : NAND2_X1 port map( A1 => IR_28_port, A2 => n391, ZN => n462);
   U1183 : NAND3_X1 port map( A1 => IR_29_port, A2 => IR_31_port, A3 => 
                           IR_30_port, ZN => n424);
   U1184 : NOR2_X1 port map( A1 => n462, A2 => n424, ZN => n356);
   U1185 : INV_X1 port map( A => IR_31_port, ZN => n393);
   U1186 : NAND3_X1 port map( A1 => IR_29_port, A2 => IR_30_port, A3 => n393, 
                           ZN => n435);
   U1187 : NAND2_X1 port map( A1 => IR_27_port, A2 => n442, ZN => n446);
   U1188 : NOR2_X1 port map( A1 => n435, A2 => n446, ZN => n394);
   U1189 : NAND2_X1 port map( A1 => n391, A2 => n422, ZN => n434);
   U1190 : INV_X1 port map( A => n474, ZN => n355);
   U1191 : OAI21_X1 port map( B1 => n434, B2 => n435, A => n355, ZN => n414);
   U1192 : AOI221_X1 port map( B1 => n356, B2 => IR_26_port, C1 => n394, C2 => 
                           n422, A => n414, ZN => n360);
   U1193 : INV_X1 port map( A => n446, ZN => n395);
   U1194 : NAND2_X1 port map( A1 => IR_26_port, A2 => n395, ZN => n425);
   U1195 : NOR3_X1 port map( A1 => IR_30_port, A2 => n393, A3 => n425, ZN => 
                           n452);
   U1196 : AOI21_X1 port map( B1 => n443, B2 => n424, A => n425, ZN => n358);
   U1197 : NAND3_X1 port map( A1 => IR_30_port, A2 => n392, A3 => n393, ZN => 
                           n447);
   U1198 : NOR3_X1 port map( A1 => n442, A2 => n391, A3 => n447, ZN => n437);
   U1199 : INV_X1 port map( A => n437, ZN => n357);
   U1200 : OAI22_X1 port map( A1 => IR_26_port, A2 => n357, B1 => n447, B2 => 
                           n425, ZN => n426);
   U1201 : AOI211_X1 port map( C1 => n452, C2 => n392, A => n358, B => n426, ZN
                           => n359);
   U1202 : AOI21_X1 port map( B1 => n360, B2 => n359, A => n322, ZN => n361);
   U1203 : AOI211_X1 port map( C1 => n465, C2 => DATAPATH_I_N60, A => n362, B 
                           => n361, ZN => n363);
   U1204 : AOI221_X1 port map( B1 => n440, B2 => n364, C1 => n456, C2 => n364, 
                           A => n363, ZN => CU_I_aluOpcode1_0_port);
   U1205 : NOR2_X1 port map( A1 => n370, A2 => n322, ZN => n374);
   U1206 : AND2_X1 port map( A1 => n330, A2 => DATAPATH_I_IF_ID_IR_20_port, ZN 
                           => n365);
   U1207 : NAND2_X1 port map( A1 => n365, A2 => n329, ZN => n373);
   U1208 : AND2_X1 port map( A1 => n366, A2 => n318, ZN => n367);
   U1209 : NAND2_X1 port map( A1 => n325, A2 => DATAPATH_I_IF_ID_IR_15_port, ZN
                           => n371);
   U1210 : AND2_X1 port map( A1 => n318, A2 => DATAPATH_I_IF_ID_IR_26_port, ZN 
                           => n369);
   U1211 : NAND2_X1 port map( A1 => n328, A2 => n369, ZN => n387);
   U1212 : AND2_X1 port map( A1 => n371, A2 => n387, ZN => n372);
   U1213 : NAND2_X1 port map( A1 => n372, A2 => n373, ZN => DATAPATH_I_N113);
   U1214 : NAND2_X1 port map( A1 => n385, A2 => DATAPATH_I_IF_ID_IR_16_port, ZN
                           => n378);
   U1215 : NAND2_X1 port map( A1 => n386, A2 => DATAPATH_I_IF_ID_IR_11_port, ZN
                           => n376);
   U1216 : NAND2_X1 port map( A1 => n378, A2 => n377, ZN => DATAPATH_I_N109);
   U1217 : NAND2_X1 port map( A1 => n385, A2 => DATAPATH_I_IF_ID_IR_17_port, ZN
                           => n381);
   U1218 : NAND2_X1 port map( A1 => n325, A2 => DATAPATH_I_IF_ID_IR_12_port, ZN
                           => n379);
   U1219 : NAND2_X1 port map( A1 => n380, A2 => n381, ZN => DATAPATH_I_N110);
   U1220 : NAND2_X1 port map( A1 => n323, A2 => DATAPATH_I_IF_ID_IR_18_port, ZN
                           => n384);
   U1221 : NAND2_X1 port map( A1 => n386, A2 => DATAPATH_I_IF_ID_IR_13_port, ZN
                           => n382);
   U1222 : NAND2_X1 port map( A1 => n384, A2 => n383, ZN => DATAPATH_I_N111);
   U1223 : NAND2_X1 port map( A1 => n323, A2 => DATAPATH_I_IF_ID_IR_19_port, ZN
                           => n390);
   U1224 : NAND2_X1 port map( A1 => n325, A2 => DATAPATH_I_IF_ID_IR_14_port, ZN
                           => n388);
   U1225 : NAND2_X1 port map( A1 => n389, A2 => n390, ZN => DATAPATH_I_N112);
   DATAPATH_I_MEM_WB_RF_WE <= '0';
   U1227 : NOR2_X1 port map( A1 => n322, A2 => n391, ZN => DATAPATH_I_N61);
   U1228 : NOR2_X1 port map( A1 => n322, A2 => n392, ZN => DATAPATH_I_N63);
   U1229 : NOR2_X1 port map( A1 => n322, A2 => n393, ZN => DATAPATH_I_N65);
   U1230 : INV_X1 port map( A => n452, ZN => n400);
   U1231 : INV_X1 port map( A => n447, ZN => n423);
   U1232 : OAI221_X1 port map( B1 => IR_28_port, B2 => n423, C1 => n442, C2 => 
                           n465, A => IR_27_port, ZN => n459);
   U1233 : OAI21_X1 port map( B1 => n437, B2 => n394, A => IR_26_port, ZN => 
                           n399);
   U1234 : INV_X1 port map( A => n424, ZN => n396);
   U1235 : OAI21_X1 port map( B1 => n397, B2 => n396, A => n395, ZN => n398);
   U1236 : NAND4_X1 port map( A1 => n400, A2 => n459, A3 => n399, A4 => n398, 
                           ZN => n413);
   U1237 : NAND2_X1 port map( A1 => IR_0_port, A2 => n401, ZN => n416);
   U1238 : INV_X1 port map( A => n416, ZN => n408);
   U1239 : NAND3_X1 port map( A1 => IR_2_port, A2 => n408, A3 => n402, ZN => 
                           n403);
   U1240 : OAI21_X1 port map( B1 => n405, B2 => n404, A => n403, ZN => n432);
   U1241 : AOI21_X1 port map( B1 => n406, B2 => n416, A => n432, ZN => n454);
   U1242 : OAI21_X1 port map( B1 => IR_0_port, B2 => n407, A => n474, ZN => 
                           n438);
   U1243 : AOI21_X1 port map( B1 => n408, B2 => n417, A => n438, ZN => n409);
   U1244 : OAI211_X1 port map( C1 => n411, C2 => n410, A => n454, B => n409, ZN
                           => n412);
   U1245 : OAI211_X1 port map( C1 => n414, C2 => n413, A => n317, B => n412, ZN
                           => CU_I_aluOpcode1_1_port);
   U1246 : AOI211_X1 port map( C1 => n417, C2 => n416, A => n415, B => n438, ZN
                           => n421);
   U1247 : INV_X1 port map( A => n418, ZN => n470);
   U1248 : NAND4_X1 port map( A1 => IR_1_port, A2 => IR_2_port, A3 => n420, A4 
                           => n419, ZN => n469);
   U1249 : NAND3_X1 port map( A1 => n421, A2 => n470, A3 => n469, ZN => n431);
   U1250 : OR2_X1 port map( A1 => n443, A2 => IR_27_port, ZN => n429);
   U1251 : NAND2_X1 port map( A1 => n462, A2 => n446, ZN => n464);
   U1252 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n461);
   U1253 : NAND3_X1 port map( A1 => n441, A2 => n461, A3 => n424, ZN => n427);
   U1254 : AOI21_X1 port map( B1 => n462, B2 => n425, A => n435, ZN => n451);
   U1255 : AOI211_X1 port map( C1 => n464, C2 => n427, A => n451, B => n426, ZN
                           => n428);
   U1256 : OAI221_X1 port map( B1 => n429, B2 => IR_26_port, C1 => n429, C2 => 
                           n442, A => n428, ZN => n430);
   U1257 : OAI211_X1 port map( C1 => n432, C2 => n431, A => n317, B => n430, ZN
                           => CU_I_aluOpcode1_2_port);
   U1258 : OR3_X1 port map( A1 => n434, A2 => n433, A3 => n447, ZN => n450);
   U1259 : AOI211_X1 port map( C1 => IR_27_port, C2 => IR_26_port, A => 
                           IR_28_port, B => n435, ZN => n436);
   U1260 : NOR2_X1 port map( A1 => n437, A2 => n436, ZN => n460);
   U1261 : NOR2_X1 port map( A1 => n439, A2 => n438, ZN => n455);
   U1262 : OAI211_X1 port map( C1 => IR_0_port, C2 => n469, A => n454, B => 
                           n440, ZN => n444);
   U1263 : AOI221_X1 port map( B1 => IR_28_port, B2 => n443, C1 => n442, C2 => 
                           n441, A => IR_27_port, ZN => n473);
   U1264 : AOI21_X1 port map( B1 => n455, B2 => n444, A => n473, ZN => n445);
   U1265 : OAI211_X1 port map( C1 => n447, C2 => n446, A => n460, B => n445, ZN
                           => n448);
   U1266 : AOI22_X1 port map( A1 => n317, A2 => n448, B1 => n452, B2 => 
                           DATAPATH_I_N63, ZN => n449);
   U1267 : NAND2_X1 port map( A1 => n450, A2 => n449, ZN => 
                           CU_I_aluOpcode1_3_port);
   U1268 : NOR2_X1 port map( A1 => n452, A2 => n451, ZN => n466);
   U1269 : AND3_X1 port map( A1 => n455, A2 => n454, A3 => n453, ZN => n471);
   U1270 : OAI21_X1 port map( B1 => n456, B2 => n469, A => n470, ZN => n457);
   U1271 : AOI21_X1 port map( B1 => n471, B2 => n457, A => n473, ZN => n458);
   U1272 : AOI21_X1 port map( B1 => n466, B2 => n458, A => n322, ZN => 
                           CU_I_aluOpcode1_4_port);
   U1273 : OAI211_X1 port map( C1 => n462, C2 => n461, A => n460, B => n459, ZN
                           => n463);
   U1274 : AOI211_X1 port map( C1 => n465, C2 => n464, A => n474, B => n463, ZN
                           => n467);
   U1275 : AOI22_X1 port map( A1 => n467, A2 => n466, B1 => n471, B2 => n470, 
                           ZN => n468);
   U1276 : NAND2_X1 port map( A1 => n317, A2 => n468, ZN => 
                           CU_I_aluOpcode1_5_port);
   U1277 : NAND3_X1 port map( A1 => n471, A2 => n470, A3 => n469, ZN => n472);
   U1278 : OAI211_X1 port map( C1 => n474, C2 => n473, A => n317, B => n472, ZN
                           => CU_I_aluOpcode1_6_port);
   n285 <= '1';

end SYN_DLX_RTL;


library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (OP_SLL, OP_SRL, OP_SRA, OP_ADD, OP_ADDU, OP_SUB, OP_SUBU, 
   OP_AND, OP_OR, OP_XOR, OP_SEQ, OP_SNE, OP_SLT, OP_SGT, OP_SLE, OP_SGE, 
   OP_MOVI2S, OP_MOVS2I, OP_MOVF, OP_MOVD, OP_MOVFP2I, OP_MOVI2FP, OP_MOVI2T, 
   OP_MOVT2I, OP_SLTU, OP_SGTU, OP_SLEU, OP_SGEU, OP_ADDF, OP_SUBF, OP_MULTF, 
   OP_DIVF, OP_ADDD, OP_SUBD, OP_MULTD, OP_DIVD, OP_CVTF2D, OP_CVTF2I, 
   OP_CVTD2F, OP_CVTD2I, OP_CVTI2F, OP_CVTI2D, OP_MULT, OP_DIV, OP_EQF, OP_NEF,
   OP_LTF, OP_GTF, OP_LEF, OP_GEF, OP_MULTU, OP_DIVU, OP_EQD, OP_NED, OP_LTD, 
   OP_GTD, OP_LED, OP_GED, OP_BEQZ, OP_BNEZ, OP_BFPT, OP_BFPF, OP_ADDI, 
   OP_ADDUI, OP_SUBI, OP_SUBUI, OP_ANDI, OP_ORI, OP_XORI, OP_LHI, OP_RFE, 
   OP_TRAP, OP_JR, OP_JALR, OP_SLLI, OP_SRLI, OP_SRAI, OP_SEQI, OP_SNEI, 
   OP_SLTI, OP_SGTI, OP_SLEI, OP_SGEI, OP_LB, OP_LH, OP_LW, OP_LBU, OP_LHU, 
   OP_LF, OP_LD, OP_SB, OP_SH, OP_SW, OP_SF, OP_SD, OP_ITLB, OP_SLTUI, 
   OP_SGTUI, OP_SLEUI, OP_SGEUI, OP_J, OP_JAL, OP_NOP);
attribute ENUM_ENCODING of aluOp : type is 
   "0000000 0000001 0000010 0000011 0000100 0000101 0000110 0000111 0001000 0001001 0001010 0001011 0001100 0001101 0001110 0001111 0010000 0010001 0010010 0010011 0010100 0010101 0010110 0010111 0011000 0011001 0011010 0011011 0011100 0011101 0011110 0011111 0100000 0100001 0100010 0100011 0100100 0100101 0100110 0100111 0101000 0101001 0101010 0101011 0101100 0101101 0101110 0101111 0110000 0110001 0110010 0110011 0110100 0110101 0110110 0110111 0111000 0111001 0111010 0111011 0111100 0111101 0111110 0111111 1000000 1000001 1000010 1000011 1000100 1000101 1000110 1000111 1001000 1001001 1001010 1001011 1001100 1001101 1001110 1001111 1010000 1010001 1010010 1010011 1010100 1010101 1010110 1010111 1011000 1011001 1011010 1011011 1011100 1011101 1011110 1011111 1100000 1100001 1100010 1100011 1100100 1100101 1100110";
   
   -- Declarations for conversion functions.
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when OP_SLL => return "0000000";
         when OP_SRL => return "0000001";
         when OP_SRA => return "0000010";
         when OP_ADD => return "0000011";
         when OP_ADDU => return "0000100";
         when OP_SUB => return "0000101";
         when OP_SUBU => return "0000110";
         when OP_AND => return "0000111";
         when OP_OR => return "0001000";
         when OP_XOR => return "0001001";
         when OP_SEQ => return "0001010";
         when OP_SNE => return "0001011";
         when OP_SLT => return "0001100";
         when OP_SGT => return "0001101";
         when OP_SLE => return "0001110";
         when OP_SGE => return "0001111";
         when OP_MOVI2S => return "0010000";
         when OP_MOVS2I => return "0010001";
         when OP_MOVF => return "0010010";
         when OP_MOVD => return "0010011";
         when OP_MOVFP2I => return "0010100";
         when OP_MOVI2FP => return "0010101";
         when OP_MOVI2T => return "0010110";
         when OP_MOVT2I => return "0010111";
         when OP_SLTU => return "0011000";
         when OP_SGTU => return "0011001";
         when OP_SLEU => return "0011010";
         when OP_SGEU => return "0011011";
         when OP_ADDF => return "0011100";
         when OP_SUBF => return "0011101";
         when OP_MULTF => return "0011110";
         when OP_DIVF => return "0011111";
         when OP_ADDD => return "0100000";
         when OP_SUBD => return "0100001";
         when OP_MULTD => return "0100010";
         when OP_DIVD => return "0100011";
         when OP_CVTF2D => return "0100100";
         when OP_CVTF2I => return "0100101";
         when OP_CVTD2F => return "0100110";
         when OP_CVTD2I => return "0100111";
         when OP_CVTI2F => return "0101000";
         when OP_CVTI2D => return "0101001";
         when OP_MULT => return "0101010";
         when OP_DIV => return "0101011";
         when OP_EQF => return "0101100";
         when OP_NEF => return "0101101";
         when OP_LTF => return "0101110";
         when OP_GTF => return "0101111";
         when OP_LEF => return "0110000";
         when OP_GEF => return "0110001";
         when OP_MULTU => return "0110010";
         when OP_DIVU => return "0110011";
         when OP_EQD => return "0110100";
         when OP_NED => return "0110101";
         when OP_LTD => return "0110110";
         when OP_GTD => return "0110111";
         when OP_LED => return "0111000";
         when OP_GED => return "0111001";
         when OP_BEQZ => return "0111010";
         when OP_BNEZ => return "0111011";
         when OP_BFPT => return "0111100";
         when OP_BFPF => return "0111101";
         when OP_ADDI => return "0111110";
         when OP_ADDUI => return "0111111";
         when OP_SUBI => return "1000000";
         when OP_SUBUI => return "1000001";
         when OP_ANDI => return "1000010";
         when OP_ORI => return "1000011";
         when OP_XORI => return "1000100";
         when OP_LHI => return "1000101";
         when OP_RFE => return "1000110";
         when OP_TRAP => return "1000111";
         when OP_JR => return "1001000";
         when OP_JALR => return "1001001";
         when OP_SLLI => return "1001010";
         when OP_SRLI => return "1001011";
         when OP_SRAI => return "1001100";
         when OP_SEQI => return "1001101";
         when OP_SNEI => return "1001110";
         when OP_SLTI => return "1001111";
         when OP_SGTI => return "1010000";
         when OP_SLEI => return "1010001";
         when OP_SGEI => return "1010010";
         when OP_LB => return "1010011";
         when OP_LH => return "1010100";
         when OP_LW => return "1010101";
         when OP_LBU => return "1010110";
         when OP_LHU => return "1010111";
         when OP_LF => return "1011000";
         when OP_LD => return "1011001";
         when OP_SB => return "1011010";
         when OP_SH => return "1011011";
         when OP_SW => return "1011100";
         when OP_SF => return "1011101";
         when OP_SD => return "1011110";
         when OP_ITLB => return "1011111";
         when OP_SLTUI => return "1100000";
         when OP_SGTUI => return "1100001";
         when OP_SLEUI => return "1100010";
         when OP_SGEUI => return "1100011";
         when OP_J => return "1100100";
         when OP_JAL => return "1100101";
         when OP_NOP => return "1100110";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

   port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  DOUT :
         out std_logic_vector (31 downto 0));

end DLX_IRAM_RAM_DEPTH256_I_SIZE32;

architecture SYN_BEHAVIORAL of DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_DRAM_N256_NW32 is

   port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector (31 
         downto 0);  DOUT : out std_logic_vector (31 downto 0));

end DLX_DRAM_N256_NW32;

architecture SYN_BEHAVIORAL of DLX_DRAM_N256_NW32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RF_N32_NA5 is

   port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
         ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_N32_NA5;

architecture SYN_BEHAVIORAL of RF_N32_NA5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REG_0_31_port, REG_0_30_port, REG_0_29_port, REG_0_28_port, 
      REG_0_27_port, REG_0_26_port, REG_0_25_port, REG_0_24_port, REG_0_23_port
      , REG_0_22_port, REG_0_21_port, REG_0_20_port, REG_0_19_port, 
      REG_0_18_port, REG_0_17_port, REG_0_16_port, REG_0_15_port, REG_0_14_port
      , REG_0_13_port, REG_0_12_port, REG_0_11_port, REG_0_10_port, 
      REG_0_9_port, REG_0_8_port, REG_0_7_port, REG_0_6_port, REG_0_5_port, 
      REG_0_4_port, REG_0_3_port, REG_0_2_port, REG_0_1_port, REG_0_0_port, 
      REG_31_31_port, REG_31_30_port, REG_31_29_port, REG_31_28_port, 
      REG_31_27_port, REG_31_26_port, REG_31_25_port, REG_31_24_port, 
      REG_31_23_port, REG_31_22_port, REG_31_21_port, REG_31_20_port, 
      REG_31_19_port, REG_31_18_port, REG_31_17_port, REG_31_16_port, 
      REG_31_15_port, REG_31_14_port, REG_31_13_port, REG_31_12_port, 
      REG_31_11_port, REG_31_10_port, REG_31_9_port, REG_31_8_port, 
      REG_31_7_port, REG_31_6_port, REG_31_5_port, REG_31_4_port, REG_31_3_port
      , REG_31_2_port, REG_31_1_port, REG_31_0_port, N156, N157, N158, N159, 
      N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, 
      N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, 
      N184, N185, N186, N187, N219, N220, N221, N222, N223, N224, N225, N226, 
      N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, 
      N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, 
      n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50 : 
      std_logic;

begin
   
   REG_reg_0_31_inst : DLH_X1 port map( G => n10, D => N250, Q => REG_0_31_port
                           );
   REG_reg_0_30_inst : DLH_X1 port map( G => n11, D => N249, Q => REG_0_30_port
                           );
   REG_reg_0_29_inst : DLH_X1 port map( G => n10, D => N248, Q => REG_0_29_port
                           );
   REG_reg_0_28_inst : DLH_X1 port map( G => n11, D => N247, Q => REG_0_28_port
                           );
   REG_reg_0_27_inst : DLH_X1 port map( G => n11, D => N246, Q => REG_0_27_port
                           );
   REG_reg_0_26_inst : DLH_X1 port map( G => n11, D => N245, Q => REG_0_26_port
                           );
   REG_reg_0_25_inst : DLH_X1 port map( G => n11, D => N244, Q => REG_0_25_port
                           );
   REG_reg_0_24_inst : DLH_X1 port map( G => n11, D => N243, Q => REG_0_24_port
                           );
   REG_reg_0_23_inst : DLH_X1 port map( G => n10, D => N242, Q => REG_0_23_port
                           );
   REG_reg_0_22_inst : DLH_X1 port map( G => n10, D => N241, Q => REG_0_22_port
                           );
   REG_reg_0_21_inst : DLH_X1 port map( G => n11, D => N240, Q => REG_0_21_port
                           );
   REG_reg_0_20_inst : DLH_X1 port map( G => n11, D => N239, Q => REG_0_20_port
                           );
   REG_reg_0_19_inst : DLH_X1 port map( G => n11, D => N238, Q => REG_0_19_port
                           );
   REG_reg_0_18_inst : DLH_X1 port map( G => n11, D => N237, Q => REG_0_18_port
                           );
   REG_reg_0_17_inst : DLH_X1 port map( G => n10, D => N236, Q => REG_0_17_port
                           );
   REG_reg_0_16_inst : DLH_X1 port map( G => n10, D => N235, Q => REG_0_16_port
                           );
   REG_reg_0_15_inst : DLH_X1 port map( G => n10, D => N234, Q => REG_0_15_port
                           );
   REG_reg_0_14_inst : DLH_X1 port map( G => n10, D => N233, Q => REG_0_14_port
                           );
   REG_reg_0_13_inst : DLH_X1 port map( G => n10, D => N232, Q => REG_0_13_port
                           );
   REG_reg_0_12_inst : DLH_X1 port map( G => n10, D => N231, Q => REG_0_12_port
                           );
   REG_reg_0_11_inst : DLH_X1 port map( G => n11, D => N230, Q => REG_0_11_port
                           );
   REG_reg_0_10_inst : DLH_X1 port map( G => n10, D => N229, Q => REG_0_10_port
                           );
   REG_reg_0_9_inst : DLH_X1 port map( G => n11, D => N228, Q => REG_0_9_port);
   REG_reg_0_8_inst : DLH_X1 port map( G => n11, D => N227, Q => REG_0_8_port);
   REG_reg_0_7_inst : DLH_X1 port map( G => n10, D => N226, Q => REG_0_7_port);
   REG_reg_0_6_inst : DLH_X1 port map( G => n10, D => N225, Q => REG_0_6_port);
   REG_reg_0_5_inst : DLH_X1 port map( G => n10, D => N224, Q => REG_0_5_port);
   REG_reg_0_4_inst : DLH_X1 port map( G => n10, D => N223, Q => REG_0_4_port);
   REG_reg_0_3_inst : DLH_X1 port map( G => n10, D => N222, Q => REG_0_3_port);
   REG_reg_0_2_inst : DLH_X1 port map( G => n10, D => N221, Q => REG_0_2_port);
   REG_reg_0_1_inst : DLH_X1 port map( G => n10, D => N220, Q => REG_0_1_port);
   REG_reg_0_0_inst : DLH_X1 port map( G => n10, D => N219, Q => REG_0_0_port);
   REG_reg_31_31_inst : DLH_X1 port map( G => n10, D => N187, Q => 
                           REG_31_31_port);
   REG_reg_31_30_inst : DLH_X1 port map( G => n10, D => N186, Q => 
                           REG_31_30_port);
   REG_reg_31_29_inst : DLH_X1 port map( G => n10, D => N185, Q => 
                           REG_31_29_port);
   REG_reg_31_28_inst : DLH_X1 port map( G => n10, D => N184, Q => 
                           REG_31_28_port);
   REG_reg_31_27_inst : DLH_X1 port map( G => n11, D => N183, Q => 
                           REG_31_27_port);
   REG_reg_31_26_inst : DLH_X1 port map( G => n11, D => N182, Q => 
                           REG_31_26_port);
   REG_reg_31_25_inst : DLH_X1 port map( G => n11, D => N181, Q => 
                           REG_31_25_port);
   REG_reg_31_24_inst : DLH_X1 port map( G => n11, D => N180, Q => 
                           REG_31_24_port);
   REG_reg_31_23_inst : DLH_X1 port map( G => n11, D => N179, Q => 
                           REG_31_23_port);
   REG_reg_31_22_inst : DLH_X1 port map( G => n11, D => N178, Q => 
                           REG_31_22_port);
   REG_reg_31_21_inst : DLH_X1 port map( G => n11, D => N177, Q => 
                           REG_31_21_port);
   REG_reg_31_20_inst : DLH_X1 port map( G => n11, D => N176, Q => 
                           REG_31_20_port);
   REG_reg_31_19_inst : DLH_X1 port map( G => n11, D => N175, Q => 
                           REG_31_19_port);
   REG_reg_31_18_inst : DLH_X1 port map( G => n11, D => N174, Q => 
                           REG_31_18_port);
   REG_reg_31_17_inst : DLH_X1 port map( G => n10, D => N173, Q => 
                           REG_31_17_port);
   REG_reg_31_16_inst : DLH_X1 port map( G => n10, D => N172, Q => 
                           REG_31_16_port);
   REG_reg_31_15_inst : DLH_X1 port map( G => n10, D => N171, Q => 
                           REG_31_15_port);
   REG_reg_31_14_inst : DLH_X1 port map( G => n10, D => N170, Q => 
                           REG_31_14_port);
   REG_reg_31_13_inst : DLH_X1 port map( G => n11, D => N169, Q => 
                           REG_31_13_port);
   REG_reg_31_12_inst : DLH_X1 port map( G => n10, D => N168, Q => 
                           REG_31_12_port);
   REG_reg_31_11_inst : DLH_X1 port map( G => n11, D => N167, Q => 
                           REG_31_11_port);
   REG_reg_31_10_inst : DLH_X1 port map( G => n10, D => N166, Q => 
                           REG_31_10_port);
   REG_reg_31_9_inst : DLH_X1 port map( G => n11, D => N165, Q => REG_31_9_port
                           );
   REG_reg_31_8_inst : DLH_X1 port map( G => n11, D => N164, Q => REG_31_8_port
                           );
   REG_reg_31_7_inst : DLH_X1 port map( G => n11, D => N163, Q => REG_31_7_port
                           );
   REG_reg_31_6_inst : DLH_X1 port map( G => n10, D => N162, Q => REG_31_6_port
                           );
   REG_reg_31_5_inst : DLH_X1 port map( G => n11, D => N161, Q => REG_31_5_port
                           );
   REG_reg_31_4_inst : DLH_X1 port map( G => n11, D => N160, Q => REG_31_4_port
                           );
   REG_reg_31_3_inst : DLH_X1 port map( G => n11, D => N159, Q => REG_31_3_port
                           );
   REG_reg_31_2_inst : DLH_X1 port map( G => n11, D => N158, Q => REG_31_2_port
                           );
   REG_reg_31_1_inst : DLH_X1 port map( G => n10, D => N157, Q => REG_31_1_port
                           );
   REG_reg_31_0_inst : DLH_X1 port map( G => n10, D => N156, Q => REG_31_0_port
                           );
   U3 : CLKBUF_X2 port map( A => n48, Z => n7);
   U4 : CLKBUF_X2 port map( A => n50, Z => n8);
   U5 : INV_X1 port map( A => RST, ZN => n10);
   U6 : INV_X1 port map( A => RST, ZN => n11);
   U7 : OR4_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), A3 => ADD_WR(0), A4 
                           => ADD_WR(2), ZN => n12);
   U8 : NOR2_X1 port map( A1 => ADD_WR(1), A2 => n12, ZN => n35);
   U9 : CLKBUF_X1 port map( A => n35, Z => n46);
   U10 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(0), ZN => n13);
   U11 : INV_X1 port map( A => n13, ZN => N156);
   U12 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(31), ZN => n45);
   U13 : INV_X1 port map( A => n45, ZN => N187);
   U14 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(30), ZN => n44);
   U15 : INV_X1 port map( A => n44, ZN => N186);
   U16 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(29), ZN => n43);
   U17 : INV_X1 port map( A => n43, ZN => N185);
   U18 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(28), ZN => n42);
   U19 : INV_X1 port map( A => n42, ZN => N184);
   U20 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(27), ZN => n41);
   U21 : INV_X1 port map( A => n41, ZN => N183);
   U22 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(26), ZN => n40);
   U23 : INV_X1 port map( A => n40, ZN => N182);
   U24 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(25), ZN => n39);
   U25 : INV_X1 port map( A => n39, ZN => N181);
   U26 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(24), ZN => n38);
   U27 : INV_X1 port map( A => n38, ZN => N180);
   U28 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(23), ZN => n37);
   U29 : INV_X1 port map( A => n37, ZN => N179);
   U30 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(22), ZN => n36);
   U31 : INV_X1 port map( A => n36, ZN => N178);
   U32 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(21), ZN => n34);
   U33 : INV_X1 port map( A => n34, ZN => N177);
   U34 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(20), ZN => n33);
   U35 : INV_X1 port map( A => n33, ZN => N176);
   U36 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(19), ZN => n32);
   U37 : INV_X1 port map( A => n32, ZN => N175);
   U38 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(18), ZN => n31);
   U39 : INV_X1 port map( A => n31, ZN => N174);
   U40 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(17), ZN => n30);
   U41 : INV_X1 port map( A => n30, ZN => N173);
   U42 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(16), ZN => n29);
   U43 : INV_X1 port map( A => n29, ZN => N172);
   U44 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(15), ZN => n28);
   U45 : INV_X1 port map( A => n28, ZN => N171);
   U46 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(14), ZN => n27);
   U47 : INV_X1 port map( A => n27, ZN => N170);
   U48 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(13), ZN => n26);
   U49 : INV_X1 port map( A => n26, ZN => N169);
   U50 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(12), ZN => n25);
   U51 : INV_X1 port map( A => n25, ZN => N168);
   U52 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(11), ZN => n24);
   U53 : INV_X1 port map( A => n24, ZN => N167);
   U54 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(10), ZN => n23);
   U55 : INV_X1 port map( A => n23, ZN => N166);
   U56 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(9), ZN => n22);
   U57 : INV_X1 port map( A => n22, ZN => N165);
   U58 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(8), ZN => n21);
   U59 : INV_X1 port map( A => n21, ZN => N164);
   U60 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(7), ZN => n20);
   U61 : INV_X1 port map( A => n20, ZN => N163);
   U62 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(6), ZN => n19);
   U63 : INV_X1 port map( A => n19, ZN => N162);
   U64 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(5), ZN => n18);
   U65 : INV_X1 port map( A => n18, ZN => N161);
   U66 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(4), ZN => n17);
   U67 : INV_X1 port map( A => n17, ZN => N160);
   U68 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(3), ZN => n16);
   U69 : INV_X1 port map( A => n16, ZN => N159);
   U70 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(2), ZN => n15);
   U71 : INV_X1 port map( A => n15, ZN => N158);
   U72 : NAND2_X1 port map( A1 => RST, A2 => DATAIN(1), ZN => n14);
   U73 : INV_X1 port map( A => n14, ZN => N157);
   U74 : NOR2_X1 port map( A1 => n46, A2 => n13, ZN => N219);
   U75 : NOR2_X1 port map( A1 => n46, A2 => n14, ZN => N220);
   U76 : NOR2_X1 port map( A1 => n46, A2 => n15, ZN => N221);
   U77 : NOR2_X1 port map( A1 => n46, A2 => n16, ZN => N222);
   U78 : NOR2_X1 port map( A1 => n46, A2 => n17, ZN => N223);
   U79 : NOR2_X1 port map( A1 => n46, A2 => n18, ZN => N224);
   U80 : NOR2_X1 port map( A1 => n46, A2 => n19, ZN => N225);
   U81 : NOR2_X1 port map( A1 => n46, A2 => n20, ZN => N226);
   U82 : NOR2_X1 port map( A1 => n46, A2 => n21, ZN => N227);
   U83 : NOR2_X1 port map( A1 => n46, A2 => n22, ZN => N228);
   U84 : NOR2_X1 port map( A1 => n35, A2 => n23, ZN => N229);
   U85 : NOR2_X1 port map( A1 => n46, A2 => n24, ZN => N230);
   U86 : NOR2_X1 port map( A1 => n46, A2 => n25, ZN => N231);
   U87 : NOR2_X1 port map( A1 => n35, A2 => n26, ZN => N232);
   U88 : NOR2_X1 port map( A1 => n35, A2 => n27, ZN => N233);
   U89 : NOR2_X1 port map( A1 => n35, A2 => n28, ZN => N234);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n29, ZN => N235);
   U91 : NOR2_X1 port map( A1 => n35, A2 => n30, ZN => N236);
   U92 : NOR2_X1 port map( A1 => n35, A2 => n31, ZN => N237);
   U93 : NOR2_X1 port map( A1 => n35, A2 => n32, ZN => N238);
   U94 : NOR2_X1 port map( A1 => n35, A2 => n33, ZN => N239);
   U95 : NOR2_X1 port map( A1 => n35, A2 => n34, ZN => N240);
   U96 : NOR2_X1 port map( A1 => n46, A2 => n36, ZN => N241);
   U97 : NOR2_X1 port map( A1 => n46, A2 => n37, ZN => N242);
   U98 : NOR2_X1 port map( A1 => n46, A2 => n38, ZN => N243);
   U99 : NOR2_X1 port map( A1 => n46, A2 => n39, ZN => N244);
   U100 : NOR2_X1 port map( A1 => n46, A2 => n40, ZN => N245);
   U101 : NOR2_X1 port map( A1 => n46, A2 => n41, ZN => N246);
   U102 : NOR2_X1 port map( A1 => n46, A2 => n42, ZN => N247);
   U103 : NOR2_X1 port map( A1 => n46, A2 => n43, ZN => N248);
   U104 : NOR2_X1 port map( A1 => n46, A2 => n44, ZN => N249);
   U105 : NOR2_X1 port map( A1 => n46, A2 => n45, ZN => N250);
   U106 : OR4_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => ADD_RD2(2)
                           , A4 => ADD_RD2(4), ZN => n47);
   U107 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => n47, ZN => n48);
   U108 : MUX2_X1 port map( A => REG_31_31_port, B => REG_0_31_port, S => n7, Z
                           => OUT2(31));
   U109 : MUX2_X1 port map( A => REG_31_30_port, B => REG_0_30_port, S => n7, Z
                           => OUT2(30));
   U110 : MUX2_X1 port map( A => REG_31_29_port, B => REG_0_29_port, S => n7, Z
                           => OUT2(29));
   U111 : MUX2_X1 port map( A => REG_31_28_port, B => REG_0_28_port, S => n7, Z
                           => OUT2(28));
   U112 : MUX2_X1 port map( A => REG_31_27_port, B => REG_0_27_port, S => n7, Z
                           => OUT2(27));
   U113 : MUX2_X1 port map( A => REG_31_26_port, B => REG_0_26_port, S => n7, Z
                           => OUT2(26));
   U114 : MUX2_X1 port map( A => REG_31_25_port, B => REG_0_25_port, S => n7, Z
                           => OUT2(25));
   U115 : MUX2_X1 port map( A => REG_31_24_port, B => REG_0_24_port, S => n7, Z
                           => OUT2(24));
   U116 : MUX2_X1 port map( A => REG_31_23_port, B => REG_0_23_port, S => n7, Z
                           => OUT2(23));
   U117 : MUX2_X1 port map( A => REG_31_22_port, B => REG_0_22_port, S => n7, Z
                           => OUT2(22));
   U118 : MUX2_X1 port map( A => REG_31_21_port, B => REG_0_21_port, S => n7, Z
                           => OUT2(21));
   U119 : MUX2_X1 port map( A => REG_31_20_port, B => REG_0_20_port, S => n7, Z
                           => OUT2(20));
   U120 : MUX2_X1 port map( A => REG_31_19_port, B => REG_0_19_port, S => n7, Z
                           => OUT2(19));
   U121 : MUX2_X1 port map( A => REG_31_18_port, B => REG_0_18_port, S => n48, 
                           Z => OUT2(18));
   U122 : MUX2_X1 port map( A => REG_31_17_port, B => REG_0_17_port, S => n48, 
                           Z => OUT2(17));
   U123 : MUX2_X1 port map( A => REG_31_16_port, B => REG_0_16_port, S => n48, 
                           Z => OUT2(16));
   U124 : MUX2_X1 port map( A => REG_31_15_port, B => REG_0_15_port, S => n48, 
                           Z => OUT2(15));
   U125 : MUX2_X1 port map( A => REG_31_14_port, B => REG_0_14_port, S => n48, 
                           Z => OUT2(14));
   U126 : MUX2_X1 port map( A => REG_31_13_port, B => REG_0_13_port, S => n48, 
                           Z => OUT2(13));
   U127 : MUX2_X1 port map( A => REG_31_12_port, B => REG_0_12_port, S => n48, 
                           Z => OUT2(12));
   U128 : MUX2_X1 port map( A => REG_31_11_port, B => REG_0_11_port, S => n48, 
                           Z => OUT2(11));
   U129 : MUX2_X1 port map( A => REG_31_10_port, B => REG_0_10_port, S => n48, 
                           Z => OUT2(10));
   U130 : MUX2_X1 port map( A => REG_31_9_port, B => REG_0_9_port, S => n7, Z 
                           => OUT2(9));
   U131 : MUX2_X1 port map( A => REG_31_8_port, B => REG_0_8_port, S => n7, Z 
                           => OUT2(8));
   U132 : MUX2_X1 port map( A => REG_31_7_port, B => REG_0_7_port, S => n7, Z 
                           => OUT2(7));
   U133 : MUX2_X1 port map( A => REG_31_6_port, B => REG_0_6_port, S => n7, Z 
                           => OUT2(6));
   U134 : MUX2_X1 port map( A => REG_31_5_port, B => REG_0_5_port, S => n7, Z 
                           => OUT2(5));
   U135 : MUX2_X1 port map( A => REG_31_4_port, B => REG_0_4_port, S => n7, Z 
                           => OUT2(4));
   U136 : MUX2_X1 port map( A => REG_31_3_port, B => REG_0_3_port, S => n7, Z 
                           => OUT2(3));
   U137 : MUX2_X1 port map( A => REG_31_2_port, B => REG_0_2_port, S => n7, Z 
                           => OUT2(2));
   U138 : MUX2_X1 port map( A => REG_31_1_port, B => REG_0_1_port, S => n7, Z 
                           => OUT2(1));
   U139 : MUX2_X1 port map( A => REG_31_0_port, B => REG_0_0_port, S => n7, Z 
                           => OUT2(0));
   U140 : OR4_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => ADD_RD1(2)
                           , A4 => ADD_RD1(4), ZN => n49);
   U141 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => n49, ZN => n50);
   U142 : MUX2_X1 port map( A => REG_31_31_port, B => REG_0_31_port, S => n8, Z
                           => OUT1(31));
   U143 : MUX2_X1 port map( A => REG_31_30_port, B => REG_0_30_port, S => n8, Z
                           => OUT1(30));
   U144 : MUX2_X1 port map( A => REG_31_29_port, B => REG_0_29_port, S => n8, Z
                           => OUT1(29));
   U145 : MUX2_X1 port map( A => REG_31_28_port, B => REG_0_28_port, S => n8, Z
                           => OUT1(28));
   U146 : MUX2_X1 port map( A => REG_31_27_port, B => REG_0_27_port, S => n8, Z
                           => OUT1(27));
   U147 : MUX2_X1 port map( A => REG_31_26_port, B => REG_0_26_port, S => n8, Z
                           => OUT1(26));
   U148 : MUX2_X1 port map( A => REG_31_25_port, B => REG_0_25_port, S => n8, Z
                           => OUT1(25));
   U149 : MUX2_X1 port map( A => REG_31_24_port, B => REG_0_24_port, S => n8, Z
                           => OUT1(24));
   U150 : MUX2_X1 port map( A => REG_31_23_port, B => REG_0_23_port, S => n8, Z
                           => OUT1(23));
   U151 : MUX2_X1 port map( A => REG_31_22_port, B => REG_0_22_port, S => n8, Z
                           => OUT1(22));
   U152 : MUX2_X1 port map( A => REG_31_21_port, B => REG_0_21_port, S => n8, Z
                           => OUT1(21));
   U153 : MUX2_X1 port map( A => REG_31_20_port, B => REG_0_20_port, S => n8, Z
                           => OUT1(20));
   U154 : MUX2_X1 port map( A => REG_31_19_port, B => REG_0_19_port, S => n8, Z
                           => OUT1(19));
   U155 : MUX2_X1 port map( A => REG_31_18_port, B => REG_0_18_port, S => n50, 
                           Z => OUT1(18));
   U156 : MUX2_X1 port map( A => REG_31_17_port, B => REG_0_17_port, S => n50, 
                           Z => OUT1(17));
   U157 : MUX2_X1 port map( A => REG_31_16_port, B => REG_0_16_port, S => n50, 
                           Z => OUT1(16));
   U158 : MUX2_X1 port map( A => REG_31_15_port, B => REG_0_15_port, S => n50, 
                           Z => OUT1(15));
   U159 : MUX2_X1 port map( A => REG_31_14_port, B => REG_0_14_port, S => n50, 
                           Z => OUT1(14));
   U160 : MUX2_X1 port map( A => REG_31_13_port, B => REG_0_13_port, S => n50, 
                           Z => OUT1(13));
   U161 : MUX2_X1 port map( A => REG_31_12_port, B => REG_0_12_port, S => n50, 
                           Z => OUT1(12));
   U162 : MUX2_X1 port map( A => REG_31_11_port, B => REG_0_11_port, S => n50, 
                           Z => OUT1(11));
   U163 : MUX2_X1 port map( A => REG_31_10_port, B => REG_0_10_port, S => n50, 
                           Z => OUT1(10));
   U164 : MUX2_X1 port map( A => REG_31_9_port, B => REG_0_9_port, S => n8, Z 
                           => OUT1(9));
   U165 : MUX2_X1 port map( A => REG_31_8_port, B => REG_0_8_port, S => n8, Z 
                           => OUT1(8));
   U166 : MUX2_X1 port map( A => REG_31_7_port, B => REG_0_7_port, S => n8, Z 
                           => OUT1(7));
   U167 : MUX2_X1 port map( A => REG_31_6_port, B => REG_0_6_port, S => n8, Z 
                           => OUT1(6));
   U168 : MUX2_X1 port map( A => REG_31_5_port, B => REG_0_5_port, S => n8, Z 
                           => OUT1(5));
   U169 : MUX2_X1 port map( A => REG_31_4_port, B => REG_0_4_port, S => n8, Z 
                           => OUT1(4));
   U170 : MUX2_X1 port map( A => REG_31_3_port, B => REG_0_3_port, S => n8, Z 
                           => OUT1(3));
   U171 : MUX2_X1 port map( A => REG_31_2_port, B => REG_0_2_port, S => n8, Z 
                           => OUT1(2));
   U172 : MUX2_X1 port map( A => REG_31_1_port, B => REG_0_1_port, S => n8, Z 
                           => OUT1(1));
   U173 : MUX2_X1 port map( A => REG_31_0_port, B => REG_0_0_port, S => n8, Z 
                           => OUT1(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_NB8 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
         std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);  Z
         : out std_logic);

end ALU_N32_NB8;

architecture SYN_BEHAVIORAL of ALU_N32_NB8 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X2
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal N96, OP_A_31_port, OP_A_30_port, OP_A_29_port, OP_A_28_port, 
      OP_A_27_port, OP_A_26_port, OP_A_25_port, OP_A_24_port, OP_A_23_port, 
      OP_A_22_port, OP_A_21_port, OP_A_20_port, OP_A_19_port, OP_A_18_port, 
      OP_A_17_port, OP_A_16_port, OP_A_15_port, OP_A_14_port, OP_A_13_port, 
      OP_A_12_port, OP_A_11_port, OP_A_10_port, OP_A_9_port, OP_A_8_port, 
      OP_A_7_port, OP_A_6_port, OP_A_5_port, OP_A_4_port, OP_A_3_port, 
      OP_A_2_port, OP_A_1_port, OP_A_0_port, OP_B_31_port, OP_B_30_port, 
      OP_B_29_port, OP_B_28_port, OP_B_27_port, OP_B_26_port, OP_B_25_port, 
      OP_B_24_port, OP_B_23_port, OP_B_22_port, OP_B_21_port, OP_B_20_port, 
      OP_B_19_port, OP_B_18_port, OP_B_17_port, OP_B_16_port, OP_B_15_port, 
      OP_B_14_port, OP_B_13_port, OP_B_12_port, OP_B_11_port, OP_B_10_port, 
      OP_B_9_port, OP_B_8_port, OP_B_7_port, OP_B_6_port, OP_B_5_port, 
      OP_B_4_port, OP_B_3_port, OP_B_2_port, OP_B_1_port, OP_B_0_port, OP_Ci, 
      OP_LOGIC_1_port, OP_LOGIC_0_port, OP_SHIFT, OP_COMPARE_3_port, 
      OP_COMPARE_2_port, OP_COMPARE_1_port, OP_COMPARE_0_port, N246, N247, N248
      , N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
      N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, 
      N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, 
      N285, N286, N287, N288, N289, C431_DATA4_3, C431_DATA4_4, C431_DATA4_5, 
      C431_DATA4_6, C431_DATA4_7, C431_DATA4_8, C431_DATA4_9, C431_DATA4_10, 
      C431_DATA4_11, C431_DATA4_12, C431_DATA4_13, C431_DATA4_14, C431_DATA4_15
      , C431_DATA4_16, C431_DATA4_17, C430_DATA4_5, C430_DATA4_6, C430_DATA4_7,
      C430_DATA4_8, C430_DATA4_9, C430_DATA4_10, C430_DATA4_11, C430_DATA4_12, 
      C430_DATA4_13, C430_DATA4_14, C430_DATA4_15, C430_DATA4_16, C430_DATA4_17
      , C430_DATA4_18, C430_DATA4_19, C429_DATA4_7, C429_DATA4_8, C429_DATA4_9,
      C429_DATA4_10, C429_DATA4_11, C429_DATA4_12, C429_DATA4_13, C429_DATA4_14
      , C429_DATA4_15, C429_DATA4_16, C429_DATA4_17, C429_DATA4_18, 
      C429_DATA4_19, C429_DATA4_20, C429_DATA4_21, C428_DATA4_1, C428_DATA4_2, 
      C428_DATA4_3, C428_DATA4_4, C428_DATA4_5, C428_DATA4_6, C428_DATA4_7, 
      C428_DATA4_8, C428_DATA4_9, C428_DATA4_10, C428_DATA4_11, C428_DATA4_12, 
      C428_DATA4_13, C428_DATA4_14, C428_DATA4_15, C2_DATA1_2, C2_DATA1_4, 
      C2_DATA1_6, DP_OP_440J3_122_9847_n80, DP_OP_440J3_122_9847_n79, 
      DP_OP_440J3_122_9847_n78, DP_OP_440J3_122_9847_n77, 
      DP_OP_440J3_122_9847_n76, DP_OP_440J3_122_9847_n75, 
      DP_OP_440J3_122_9847_n74, DP_OP_440J3_122_9847_n73, 
      DP_OP_440J3_122_9847_n72, DP_OP_440J3_122_9847_n71, 
      DP_OP_440J3_122_9847_n70, DP_OP_440J3_122_9847_n69, 
      DP_OP_440J3_122_9847_n68, DP_OP_440J3_122_9847_n67, 
      DP_OP_440J3_122_9847_n66, DP_OP_440J3_122_9847_n35, 
      DP_OP_440J3_122_9847_n34, DP_OP_440J3_122_9847_n33, 
      DP_OP_440J3_122_9847_n32, DP_OP_440J3_122_9847_n31, 
      DP_OP_440J3_122_9847_n30, DP_OP_440J3_122_9847_n29, 
      DP_OP_440J3_122_9847_n28, DP_OP_440J3_122_9847_n27, 
      DP_OP_440J3_122_9847_n26, DP_OP_440J3_122_9847_n25, 
      DP_OP_440J3_122_9847_n24, DP_OP_440J3_122_9847_n23, 
      DP_OP_440J3_122_9847_n22, DP_OP_440J3_122_9847_n21, 
      DP_OP_440J3_122_9847_n20, DP_OP_446J3_125_4819_n87, 
      DP_OP_446J3_125_4819_n86, DP_OP_446J3_125_4819_n85, 
      DP_OP_446J3_125_4819_n84, DP_OP_446J3_125_4819_n83, 
      DP_OP_446J3_125_4819_n82, DP_OP_446J3_125_4819_n81, 
      DP_OP_446J3_125_4819_n80, DP_OP_446J3_125_4819_n79, 
      DP_OP_446J3_125_4819_n78, DP_OP_446J3_125_4819_n77, 
      DP_OP_446J3_125_4819_n76, DP_OP_446J3_125_4819_n75, 
      DP_OP_446J3_125_4819_n74, DP_OP_446J3_125_4819_n73, 
      DP_OP_446J3_125_4819_n72, DP_OP_446J3_125_4819_n27, 
      DP_OP_446J3_125_4819_n26, DP_OP_446J3_125_4819_n25, 
      DP_OP_446J3_125_4819_n24, DP_OP_446J3_125_4819_n23, 
      DP_OP_446J3_125_4819_n22, DP_OP_446J3_125_4819_n21, 
      DP_OP_446J3_125_4819_n20, DP_OP_446J3_125_4819_n19, 
      DP_OP_446J3_125_4819_n18, DP_OP_446J3_125_4819_n17, 
      DP_OP_446J3_125_4819_n16, DP_OP_446J3_125_4819_n15, 
      DP_OP_446J3_125_4819_n14, DP_OP_446J3_125_4819_n13, 
      DP_OP_446J3_125_4819_n12, DP_OP_451J3_128_3502_n85, 
      DP_OP_451J3_128_3502_n84, DP_OP_451J3_128_3502_n83, 
      DP_OP_451J3_128_3502_n82, DP_OP_451J3_128_3502_n81, 
      DP_OP_451J3_128_3502_n80, DP_OP_451J3_128_3502_n79, 
      DP_OP_451J3_128_3502_n78, DP_OP_451J3_128_3502_n77, 
      DP_OP_451J3_128_3502_n76, DP_OP_451J3_128_3502_n75, 
      DP_OP_451J3_128_3502_n74, DP_OP_451J3_128_3502_n73, 
      DP_OP_451J3_128_3502_n72, DP_OP_451J3_128_3502_n71, 
      DP_OP_451J3_128_3502_n70, DP_OP_451J3_128_3502_n30, 
      DP_OP_451J3_128_3502_n29, DP_OP_451J3_128_3502_n28, 
      DP_OP_451J3_128_3502_n27, DP_OP_451J3_128_3502_n26, 
      DP_OP_451J3_128_3502_n25, DP_OP_451J3_128_3502_n24, 
      DP_OP_451J3_128_3502_n23, DP_OP_451J3_128_3502_n22, 
      DP_OP_451J3_128_3502_n21, DP_OP_451J3_128_3502_n20, 
      DP_OP_451J3_128_3502_n19, DP_OP_451J3_128_3502_n18, 
      DP_OP_451J3_128_3502_n17, DP_OP_451J3_128_3502_n16, 
      DP_OP_451J3_128_3502_n15, DP_OP_456J3_131_2158_n82, 
      DP_OP_456J3_131_2158_n81, DP_OP_456J3_131_2158_n80, 
      DP_OP_456J3_131_2158_n79, DP_OP_456J3_131_2158_n78, 
      DP_OP_456J3_131_2158_n77, DP_OP_456J3_131_2158_n76, 
      DP_OP_456J3_131_2158_n75, DP_OP_456J3_131_2158_n74, 
      DP_OP_456J3_131_2158_n73, DP_OP_456J3_131_2158_n72, 
      DP_OP_456J3_131_2158_n71, DP_OP_456J3_131_2158_n70, 
      DP_OP_456J3_131_2158_n69, DP_OP_456J3_131_2158_n68, 
      DP_OP_456J3_131_2158_n67, DP_OP_456J3_131_2158_n32, 
      DP_OP_456J3_131_2158_n31, DP_OP_456J3_131_2158_n30, 
      DP_OP_456J3_131_2158_n29, DP_OP_456J3_131_2158_n28, 
      DP_OP_456J3_131_2158_n27, DP_OP_456J3_131_2158_n26, 
      DP_OP_456J3_131_2158_n25, DP_OP_456J3_131_2158_n24, 
      DP_OP_456J3_131_2158_n23, DP_OP_456J3_131_2158_n22, 
      DP_OP_456J3_131_2158_n21, DP_OP_456J3_131_2158_n20, 
      DP_OP_456J3_131_2158_n19, DP_OP_456J3_131_2158_n18, 
      DP_OP_456J3_131_2158_n17, intadd_0_A_16_port, intadd_0_A_12_port, 
      intadd_0_A_11_port, intadd_0_A_10_port, intadd_0_A_9_port, 
      intadd_0_A_8_port, intadd_0_A_7_port, intadd_0_A_6_port, 
      intadd_0_A_5_port, intadd_0_A_4_port, intadd_0_A_3_port, 
      intadd_0_A_2_port, intadd_0_A_1_port, intadd_0_A_0_port, 
      intadd_0_B_14_port, intadd_0_B_13_port, intadd_0_B_12_port, 
      intadd_0_B_11_port, intadd_0_B_10_port, intadd_0_B_9_port, 
      intadd_0_B_8_port, intadd_0_B_7_port, intadd_0_B_6_port, 
      intadd_0_B_5_port, intadd_0_B_4_port, intadd_0_B_3_port, 
      intadd_0_B_2_port, intadd_0_B_1_port, intadd_0_B_0_port, intadd_0_CI, 
      intadd_0_SUM_26_port, intadd_0_SUM_25_port, intadd_0_SUM_24_port, 
      intadd_0_SUM_23_port, intadd_0_SUM_22_port, intadd_0_SUM_21_port, 
      intadd_0_SUM_20_port, intadd_0_SUM_19_port, intadd_0_SUM_18_port, 
      intadd_0_SUM_17_port, intadd_0_SUM_16_port, intadd_0_SUM_15_port, 
      intadd_0_SUM_14_port, intadd_0_SUM_13_port, intadd_0_SUM_12_port, 
      intadd_0_SUM_11_port, intadd_0_SUM_10_port, intadd_0_SUM_9_port, 
      intadd_0_SUM_8_port, intadd_0_SUM_7_port, intadd_0_SUM_6_port, 
      intadd_0_SUM_5_port, intadd_0_SUM_4_port, intadd_0_SUM_3_port, 
      intadd_0_SUM_2_port, intadd_0_SUM_1_port, intadd_0_SUM_0_port, 
      intadd_0_n27, intadd_0_n26, intadd_0_n25, intadd_0_n24, intadd_0_n23, 
      intadd_0_n22, intadd_0_n21, intadd_0_n20, intadd_0_n19, intadd_0_n18, 
      intadd_0_n17, intadd_0_n16, intadd_0_n15, intadd_0_n14, intadd_0_n13, 
      intadd_0_n12, intadd_0_n11, intadd_0_n10, intadd_0_n9, intadd_0_n8, 
      intadd_0_n7, intadd_0_n6, intadd_0_n5, intadd_0_n4, intadd_0_n3, 
      intadd_0_n2, intadd_0_n1, intadd_1_A_0_port, intadd_1_B_18_port, 
      intadd_1_B_14_port, intadd_1_B_13_port, intadd_1_B_12_port, 
      intadd_1_B_11_port, intadd_1_B_10_port, intadd_1_B_9_port, 
      intadd_1_B_8_port, intadd_1_B_7_port, intadd_1_B_6_port, 
      intadd_1_B_5_port, intadd_1_B_4_port, intadd_1_B_3_port, 
      intadd_1_B_2_port, intadd_1_B_1_port, intadd_1_B_0_port, 
      intadd_1_SUM_24_port, intadd_1_SUM_23_port, intadd_1_SUM_22_port, 
      intadd_1_SUM_21_port, intadd_1_SUM_20_port, intadd_1_SUM_19_port, 
      intadd_1_SUM_18_port, intadd_1_SUM_17_port, intadd_1_SUM_16_port, 
      intadd_1_SUM_15_port, intadd_1_SUM_14_port, intadd_1_SUM_13_port, 
      intadd_1_SUM_12_port, intadd_1_SUM_11_port, intadd_1_SUM_10_port, 
      intadd_1_SUM_9_port, intadd_1_SUM_8_port, intadd_1_SUM_7_port, 
      intadd_1_SUM_6_port, intadd_1_SUM_5_port, intadd_1_SUM_4_port, 
      intadd_1_SUM_3_port, intadd_1_SUM_2_port, intadd_1_SUM_1_port, 
      intadd_1_SUM_0_port, intadd_1_n25, intadd_1_n24, intadd_1_n23, 
      intadd_1_n22, intadd_1_n21, intadd_1_n20, intadd_1_n19, intadd_1_n18, 
      intadd_1_n17, intadd_1_n16, intadd_1_n15, intadd_1_n14, intadd_1_n13, 
      intadd_1_n12, intadd_1_n11, intadd_1_n10, intadd_1_n9, intadd_1_n8, 
      intadd_1_n7, intadd_1_n6, intadd_1_n5, intadd_1_n4, intadd_1_n3, 
      intadd_1_n2, intadd_1_n1, intadd_2_A_9_port, intadd_2_A_8_port, 
      intadd_2_A_7_port, intadd_2_A_6_port, intadd_2_A_5_port, 
      intadd_2_A_4_port, intadd_2_A_3_port, intadd_2_A_2_port, 
      intadd_2_A_1_port, intadd_2_A_0_port, intadd_2_B_0_port, 
      intadd_2_SUM_9_port, intadd_2_SUM_8_port, intadd_2_SUM_7_port, 
      intadd_2_SUM_6_port, intadd_2_SUM_5_port, intadd_2_SUM_4_port, 
      intadd_2_SUM_3_port, intadd_2_SUM_2_port, intadd_2_SUM_1_port, 
      intadd_2_SUM_0_port, intadd_2_n10, intadd_2_n9, intadd_2_n8, intadd_2_n7,
      intadd_2_n6, intadd_2_n5, intadd_2_n4, intadd_2_n3, intadd_2_n2, 
      intadd_2_n1, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
      n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96_port, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246_port, n247_port, n248_port, 
      n249_port, n250_port, n251_port, n252_port, n253_port, n254_port, 
      n255_port, n256_port, n257_port, n258_port, n259_port, n260_port, 
      n261_port, n262_port, n263_port, n264_port, n265_port, n266_port, 
      n267_port, n268_port, n269_port, n270_port, n271_port, n272_port, 
      n273_port, n274_port, n275_port, n276_port, n277_port, n278_port, 
      n279_port, n280_port, n281_port, n282_port, n283_port, n284_port, 
      n285_port, n286_port, n287_port, n288_port, n289_port, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
      n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, 
      n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
      n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
      n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
      n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, 
      n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
      n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
      n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n1415, n_1170 : std_logic;

begin
   
   OP_COMPARE_reg_3_inst : DLH_X1 port map( G => N285, D => N289, Q => 
                           OP_COMPARE_3_port);
   OP_COMPARE_reg_2_inst : DLH_X1 port map( G => N285, D => N288, Q => 
                           OP_COMPARE_2_port);
   OP_COMPARE_reg_1_inst : DLH_X1 port map( G => N285, D => N287, Q => 
                           OP_COMPARE_1_port);
   OP_COMPARE_reg_0_inst : DLH_X1 port map( G => N285, D => N286, Q => 
                           OP_COMPARE_0_port);
   OP_A_reg_31_inst : DLH_X1 port map( G => n1412, D => OP1(31), Q => 
                           OP_A_31_port);
   OP_A_reg_30_inst : DLH_X1 port map( G => n1412, D => OP1(30), Q => 
                           OP_A_30_port);
   OP_A_reg_29_inst : DLH_X1 port map( G => n1412, D => OP1(29), Q => 
                           OP_A_29_port);
   OP_A_reg_28_inst : DLH_X1 port map( G => n1412, D => OP1(28), Q => 
                           OP_A_28_port);
   OP_A_reg_27_inst : DLH_X1 port map( G => N246, D => OP1(27), Q => 
                           OP_A_27_port);
   OP_A_reg_26_inst : DLH_X1 port map( G => N246, D => OP1(26), Q => 
                           OP_A_26_port);
   OP_A_reg_25_inst : DLH_X1 port map( G => N246, D => OP1(25), Q => 
                           OP_A_25_port);
   OP_A_reg_24_inst : DLH_X1 port map( G => n1412, D => OP1(24), Q => 
                           OP_A_24_port);
   OP_A_reg_23_inst : DLH_X1 port map( G => N246, D => OP1(23), Q => 
                           OP_A_23_port);
   OP_A_reg_22_inst : DLH_X1 port map( G => n1412, D => OP1(22), Q => 
                           OP_A_22_port);
   OP_A_reg_21_inst : DLH_X1 port map( G => n1412, D => OP1(21), Q => 
                           OP_A_21_port);
   OP_A_reg_20_inst : DLH_X1 port map( G => N246, D => OP1(20), Q => 
                           OP_A_20_port);
   OP_A_reg_19_inst : DLH_X1 port map( G => N246, D => OP1(19), Q => 
                           OP_A_19_port);
   OP_A_reg_18_inst : DLH_X1 port map( G => n1412, D => OP1(18), Q => 
                           OP_A_18_port);
   OP_A_reg_17_inst : DLH_X1 port map( G => n1412, D => OP1(17), Q => 
                           OP_A_17_port);
   OP_A_reg_16_inst : DLH_X1 port map( G => n1412, D => OP1(16), Q => 
                           OP_A_16_port);
   OP_B_reg_31_inst : DLH_X1 port map( G => N246, D => N278, Q => OP_B_31_port)
                           ;
   OP_B_reg_30_inst : DLH_X1 port map( G => n1412, D => N277, Q => OP_B_30_port
                           );
   OP_B_reg_29_inst : DLH_X1 port map( G => N246, D => N276, Q => OP_B_29_port)
                           ;
   OP_B_reg_28_inst : DLH_X1 port map( G => N246, D => N275, Q => OP_B_28_port)
                           ;
   OP_B_reg_27_inst : DLH_X1 port map( G => N246, D => N274, Q => OP_B_27_port)
                           ;
   OP_B_reg_26_inst : DLH_X1 port map( G => N246, D => N273, Q => OP_B_26_port)
                           ;
   OP_B_reg_25_inst : DLH_X1 port map( G => N246, D => N272, Q => OP_B_25_port)
                           ;
   OP_B_reg_24_inst : DLH_X1 port map( G => N246, D => N271, Q => OP_B_24_port)
                           ;
   OP_B_reg_23_inst : DLH_X1 port map( G => N246, D => N270, Q => OP_B_23_port)
                           ;
   OP_B_reg_22_inst : DLH_X1 port map( G => N246, D => N269, Q => OP_B_22_port)
                           ;
   OP_B_reg_21_inst : DLH_X1 port map( G => N246, D => N268, Q => OP_B_21_port)
                           ;
   OP_B_reg_20_inst : DLH_X1 port map( G => N246, D => N267, Q => OP_B_20_port)
                           ;
   OP_B_reg_19_inst : DLH_X1 port map( G => n1412, D => N266, Q => OP_B_19_port
                           );
   OP_B_reg_18_inst : DLH_X1 port map( G => n1412, D => N265, Q => OP_B_18_port
                           );
   OP_B_reg_17_inst : DLH_X1 port map( G => n1412, D => N264, Q => OP_B_17_port
                           );
   OP_B_reg_16_inst : DLH_X1 port map( G => n1412, D => N263, Q => OP_B_16_port
                           );
   OP_B_reg_15_inst : DLH_X1 port map( G => n1412, D => N262, Q => OP_B_15_port
                           );
   OP_B_reg_14_inst : DLH_X1 port map( G => n1412, D => N261, Q => OP_B_14_port
                           );
   OP_B_reg_13_inst : DLH_X1 port map( G => n1412, D => N260, Q => OP_B_13_port
                           );
   OP_B_reg_12_inst : DLH_X1 port map( G => n1412, D => N259, Q => OP_B_12_port
                           );
   OP_B_reg_11_inst : DLH_X1 port map( G => n1412, D => N258, Q => OP_B_11_port
                           );
   OP_B_reg_10_inst : DLH_X1 port map( G => n1412, D => N257, Q => OP_B_10_port
                           );
   OP_B_reg_9_inst : DLH_X1 port map( G => N246, D => N256, Q => OP_B_9_port);
   OP_B_reg_8_inst : DLH_X1 port map( G => N246, D => N255, Q => OP_B_8_port);
   OP_B_reg_7_inst : DLH_X1 port map( G => n1412, D => N254, Q => OP_B_7_port);
   OP_B_reg_6_inst : DLH_X1 port map( G => N246, D => N253, Q => OP_B_6_port);
   OP_B_reg_0_inst : DLH_X1 port map( G => n1412, D => N247, Q => OP_B_0_port);
   OP_Ci_reg : DLH_X1 port map( G => N279, D => N280, Q => OP_Ci);
   OP_LOGIC_reg_1_inst : DLH_X1 port map( G => N281, D => N283, Q => 
                           OP_LOGIC_1_port);
   OP_LOGIC_reg_0_inst : DLH_X1 port map( G => N281, D => N282, Q => 
                           OP_LOGIC_0_port);
   OP_SHIFT_reg : DLH_X1 port map( G => N284, D => N96, Q => OP_SHIFT);
   DP_OP_440J3_122_9847_U43 : HA_X1 port map( A => DP_OP_440J3_122_9847_n35, B 
                           => DP_OP_440J3_122_9847_n66, CO => 
                           DP_OP_440J3_122_9847_n34, S => C428_DATA4_1);
   DP_OP_440J3_122_9847_U42 : HA_X1 port map( A => DP_OP_440J3_122_9847_n34, B 
                           => DP_OP_440J3_122_9847_n67, CO => 
                           DP_OP_440J3_122_9847_n33, S => C428_DATA4_2);
   DP_OP_440J3_122_9847_U41 : HA_X1 port map( A => DP_OP_440J3_122_9847_n33, B 
                           => DP_OP_440J3_122_9847_n68, CO => 
                           DP_OP_440J3_122_9847_n32, S => C428_DATA4_3);
   DP_OP_440J3_122_9847_U40 : HA_X1 port map( A => DP_OP_440J3_122_9847_n32, B 
                           => DP_OP_440J3_122_9847_n69, CO => 
                           DP_OP_440J3_122_9847_n31, S => C428_DATA4_4);
   DP_OP_440J3_122_9847_U39 : HA_X1 port map( A => DP_OP_440J3_122_9847_n31, B 
                           => DP_OP_440J3_122_9847_n70, CO => 
                           DP_OP_440J3_122_9847_n30, S => C428_DATA4_5);
   DP_OP_440J3_122_9847_U38 : HA_X1 port map( A => DP_OP_440J3_122_9847_n30, B 
                           => DP_OP_440J3_122_9847_n71, CO => 
                           DP_OP_440J3_122_9847_n29, S => C428_DATA4_6);
   DP_OP_440J3_122_9847_U37 : HA_X1 port map( A => DP_OP_440J3_122_9847_n29, B 
                           => DP_OP_440J3_122_9847_n72, CO => 
                           DP_OP_440J3_122_9847_n28, S => C428_DATA4_7);
   DP_OP_440J3_122_9847_U36 : HA_X1 port map( A => DP_OP_440J3_122_9847_n28, B 
                           => DP_OP_440J3_122_9847_n73, CO => 
                           DP_OP_440J3_122_9847_n27, S => C428_DATA4_8);
   DP_OP_440J3_122_9847_U35 : HA_X1 port map( A => DP_OP_440J3_122_9847_n27, B 
                           => DP_OP_440J3_122_9847_n74, CO => 
                           DP_OP_440J3_122_9847_n26, S => C428_DATA4_9);
   DP_OP_440J3_122_9847_U34 : HA_X1 port map( A => DP_OP_440J3_122_9847_n26, B 
                           => DP_OP_440J3_122_9847_n75, CO => 
                           DP_OP_440J3_122_9847_n25, S => C428_DATA4_10);
   DP_OP_440J3_122_9847_U33 : HA_X1 port map( A => DP_OP_440J3_122_9847_n25, B 
                           => DP_OP_440J3_122_9847_n76, CO => 
                           DP_OP_440J3_122_9847_n24, S => C428_DATA4_11);
   DP_OP_440J3_122_9847_U32 : HA_X1 port map( A => DP_OP_440J3_122_9847_n24, B 
                           => DP_OP_440J3_122_9847_n77, CO => 
                           DP_OP_440J3_122_9847_n23, S => C428_DATA4_12);
   DP_OP_440J3_122_9847_U31 : HA_X1 port map( A => DP_OP_440J3_122_9847_n23, B 
                           => DP_OP_440J3_122_9847_n78, CO => 
                           DP_OP_440J3_122_9847_n22, S => C428_DATA4_13);
   DP_OP_440J3_122_9847_U30 : HA_X1 port map( A => DP_OP_440J3_122_9847_n22, B 
                           => DP_OP_440J3_122_9847_n79, CO => 
                           DP_OP_440J3_122_9847_n21, S => C428_DATA4_14);
   DP_OP_440J3_122_9847_U29 : HA_X1 port map( A => DP_OP_440J3_122_9847_n21, B 
                           => DP_OP_440J3_122_9847_n80, CO => 
                           DP_OP_440J3_122_9847_n20, S => C428_DATA4_15);
   DP_OP_446J3_125_4819_U33 : HA_X1 port map( A => n1414, B => 
                           DP_OP_446J3_125_4819_n72, CO => 
                           DP_OP_446J3_125_4819_n27, S => C2_DATA1_6);
   DP_OP_446J3_125_4819_U32 : HA_X1 port map( A => DP_OP_446J3_125_4819_n27, B 
                           => DP_OP_446J3_125_4819_n73, CO => 
                           DP_OP_446J3_125_4819_n26, S => C429_DATA4_7);
   DP_OP_446J3_125_4819_U31 : HA_X1 port map( A => DP_OP_446J3_125_4819_n26, B 
                           => DP_OP_446J3_125_4819_n74, CO => 
                           DP_OP_446J3_125_4819_n25, S => C429_DATA4_8);
   DP_OP_446J3_125_4819_U30 : HA_X1 port map( A => DP_OP_446J3_125_4819_n25, B 
                           => DP_OP_446J3_125_4819_n75, CO => 
                           DP_OP_446J3_125_4819_n24, S => C429_DATA4_9);
   DP_OP_446J3_125_4819_U29 : HA_X1 port map( A => DP_OP_446J3_125_4819_n24, B 
                           => DP_OP_446J3_125_4819_n76, CO => 
                           DP_OP_446J3_125_4819_n23, S => C429_DATA4_10);
   DP_OP_446J3_125_4819_U28 : HA_X1 port map( A => DP_OP_446J3_125_4819_n23, B 
                           => DP_OP_446J3_125_4819_n77, CO => 
                           DP_OP_446J3_125_4819_n22, S => C429_DATA4_11);
   DP_OP_446J3_125_4819_U27 : HA_X1 port map( A => DP_OP_446J3_125_4819_n22, B 
                           => DP_OP_446J3_125_4819_n78, CO => 
                           DP_OP_446J3_125_4819_n21, S => C429_DATA4_12);
   DP_OP_446J3_125_4819_U26 : HA_X1 port map( A => DP_OP_446J3_125_4819_n21, B 
                           => DP_OP_446J3_125_4819_n79, CO => 
                           DP_OP_446J3_125_4819_n20, S => C429_DATA4_13);
   DP_OP_446J3_125_4819_U25 : HA_X1 port map( A => DP_OP_446J3_125_4819_n20, B 
                           => DP_OP_446J3_125_4819_n80, CO => 
                           DP_OP_446J3_125_4819_n19, S => C429_DATA4_14);
   DP_OP_446J3_125_4819_U24 : HA_X1 port map( A => DP_OP_446J3_125_4819_n19, B 
                           => DP_OP_446J3_125_4819_n81, CO => 
                           DP_OP_446J3_125_4819_n18, S => C429_DATA4_15);
   DP_OP_446J3_125_4819_U23 : HA_X1 port map( A => DP_OP_446J3_125_4819_n18, B 
                           => DP_OP_446J3_125_4819_n82, CO => 
                           DP_OP_446J3_125_4819_n17, S => C429_DATA4_16);
   DP_OP_446J3_125_4819_U22 : HA_X1 port map( A => DP_OP_446J3_125_4819_n17, B 
                           => DP_OP_446J3_125_4819_n83, CO => 
                           DP_OP_446J3_125_4819_n16, S => C429_DATA4_17);
   DP_OP_446J3_125_4819_U21 : HA_X1 port map( A => DP_OP_446J3_125_4819_n16, B 
                           => DP_OP_446J3_125_4819_n84, CO => 
                           DP_OP_446J3_125_4819_n15, S => C429_DATA4_18);
   DP_OP_446J3_125_4819_U20 : HA_X1 port map( A => DP_OP_446J3_125_4819_n15, B 
                           => DP_OP_446J3_125_4819_n85, CO => 
                           DP_OP_446J3_125_4819_n14, S => C429_DATA4_19);
   DP_OP_446J3_125_4819_U19 : HA_X1 port map( A => DP_OP_446J3_125_4819_n14, B 
                           => DP_OP_446J3_125_4819_n86, CO => 
                           DP_OP_446J3_125_4819_n13, S => C429_DATA4_20);
   DP_OP_446J3_125_4819_U18 : HA_X1 port map( A => DP_OP_446J3_125_4819_n13, B 
                           => DP_OP_446J3_125_4819_n87, CO => 
                           DP_OP_446J3_125_4819_n12, S => C429_DATA4_21);
   DP_OP_451J3_128_3502_U37 : HA_X1 port map( A => n1413, B => 
                           DP_OP_451J3_128_3502_n70, CO => 
                           DP_OP_451J3_128_3502_n30, S => C2_DATA1_4);
   DP_OP_451J3_128_3502_U36 : HA_X1 port map( A => DP_OP_451J3_128_3502_n30, B 
                           => DP_OP_451J3_128_3502_n71, CO => 
                           DP_OP_451J3_128_3502_n29, S => C430_DATA4_5);
   DP_OP_451J3_128_3502_U35 : HA_X1 port map( A => DP_OP_451J3_128_3502_n29, B 
                           => DP_OP_451J3_128_3502_n72, CO => 
                           DP_OP_451J3_128_3502_n28, S => C430_DATA4_6);
   DP_OP_451J3_128_3502_U34 : HA_X1 port map( A => DP_OP_451J3_128_3502_n28, B 
                           => DP_OP_451J3_128_3502_n73, CO => 
                           DP_OP_451J3_128_3502_n27, S => C430_DATA4_7);
   DP_OP_451J3_128_3502_U33 : HA_X1 port map( A => DP_OP_451J3_128_3502_n27, B 
                           => DP_OP_451J3_128_3502_n74, CO => 
                           DP_OP_451J3_128_3502_n26, S => C430_DATA4_8);
   DP_OP_451J3_128_3502_U32 : HA_X1 port map( A => DP_OP_451J3_128_3502_n26, B 
                           => DP_OP_451J3_128_3502_n75, CO => 
                           DP_OP_451J3_128_3502_n25, S => C430_DATA4_9);
   DP_OP_451J3_128_3502_U31 : HA_X1 port map( A => DP_OP_451J3_128_3502_n25, B 
                           => DP_OP_451J3_128_3502_n76, CO => 
                           DP_OP_451J3_128_3502_n24, S => C430_DATA4_10);
   DP_OP_451J3_128_3502_U30 : HA_X1 port map( A => DP_OP_451J3_128_3502_n24, B 
                           => DP_OP_451J3_128_3502_n77, CO => 
                           DP_OP_451J3_128_3502_n23, S => C430_DATA4_11);
   DP_OP_451J3_128_3502_U29 : HA_X1 port map( A => DP_OP_451J3_128_3502_n23, B 
                           => DP_OP_451J3_128_3502_n78, CO => 
                           DP_OP_451J3_128_3502_n22, S => C430_DATA4_12);
   DP_OP_451J3_128_3502_U28 : HA_X1 port map( A => DP_OP_451J3_128_3502_n22, B 
                           => DP_OP_451J3_128_3502_n79, CO => 
                           DP_OP_451J3_128_3502_n21, S => C430_DATA4_13);
   DP_OP_451J3_128_3502_U27 : HA_X1 port map( A => DP_OP_451J3_128_3502_n21, B 
                           => DP_OP_451J3_128_3502_n80, CO => 
                           DP_OP_451J3_128_3502_n20, S => C430_DATA4_14);
   DP_OP_451J3_128_3502_U26 : HA_X1 port map( A => DP_OP_451J3_128_3502_n20, B 
                           => DP_OP_451J3_128_3502_n81, CO => 
                           DP_OP_451J3_128_3502_n19, S => C430_DATA4_15);
   DP_OP_451J3_128_3502_U25 : HA_X1 port map( A => DP_OP_451J3_128_3502_n19, B 
                           => DP_OP_451J3_128_3502_n82, CO => 
                           DP_OP_451J3_128_3502_n18, S => C430_DATA4_16);
   DP_OP_451J3_128_3502_U24 : HA_X1 port map( A => DP_OP_451J3_128_3502_n18, B 
                           => DP_OP_451J3_128_3502_n83, CO => 
                           DP_OP_451J3_128_3502_n17, S => C430_DATA4_17);
   DP_OP_451J3_128_3502_U23 : HA_X1 port map( A => DP_OP_451J3_128_3502_n17, B 
                           => DP_OP_451J3_128_3502_n84, CO => 
                           DP_OP_451J3_128_3502_n16, S => C430_DATA4_18);
   DP_OP_451J3_128_3502_U22 : HA_X1 port map( A => DP_OP_451J3_128_3502_n16, B 
                           => DP_OP_451J3_128_3502_n85, CO => 
                           DP_OP_451J3_128_3502_n15, S => C430_DATA4_19);
   DP_OP_456J3_131_2158_U40 : HA_X1 port map( A => n1415, B => 
                           DP_OP_456J3_131_2158_n67, CO => 
                           DP_OP_456J3_131_2158_n32, S => C2_DATA1_2);
   DP_OP_456J3_131_2158_U39 : HA_X1 port map( A => DP_OP_456J3_131_2158_n32, B 
                           => DP_OP_456J3_131_2158_n68, CO => 
                           DP_OP_456J3_131_2158_n31, S => C431_DATA4_3);
   DP_OP_456J3_131_2158_U38 : HA_X1 port map( A => DP_OP_456J3_131_2158_n31, B 
                           => DP_OP_456J3_131_2158_n69, CO => 
                           DP_OP_456J3_131_2158_n30, S => C431_DATA4_4);
   DP_OP_456J3_131_2158_U37 : HA_X1 port map( A => DP_OP_456J3_131_2158_n30, B 
                           => DP_OP_456J3_131_2158_n70, CO => 
                           DP_OP_456J3_131_2158_n29, S => C431_DATA4_5);
   DP_OP_456J3_131_2158_U36 : HA_X1 port map( A => DP_OP_456J3_131_2158_n29, B 
                           => DP_OP_456J3_131_2158_n71, CO => 
                           DP_OP_456J3_131_2158_n28, S => C431_DATA4_6);
   DP_OP_456J3_131_2158_U35 : HA_X1 port map( A => DP_OP_456J3_131_2158_n28, B 
                           => DP_OP_456J3_131_2158_n72, CO => 
                           DP_OP_456J3_131_2158_n27, S => C431_DATA4_7);
   DP_OP_456J3_131_2158_U34 : HA_X1 port map( A => DP_OP_456J3_131_2158_n27, B 
                           => DP_OP_456J3_131_2158_n73, CO => 
                           DP_OP_456J3_131_2158_n26, S => C431_DATA4_8);
   DP_OP_456J3_131_2158_U33 : HA_X1 port map( A => DP_OP_456J3_131_2158_n26, B 
                           => DP_OP_456J3_131_2158_n74, CO => 
                           DP_OP_456J3_131_2158_n25, S => C431_DATA4_9);
   DP_OP_456J3_131_2158_U32 : HA_X1 port map( A => DP_OP_456J3_131_2158_n25, B 
                           => DP_OP_456J3_131_2158_n75, CO => 
                           DP_OP_456J3_131_2158_n24, S => C431_DATA4_10);
   DP_OP_456J3_131_2158_U31 : HA_X1 port map( A => DP_OP_456J3_131_2158_n24, B 
                           => DP_OP_456J3_131_2158_n76, CO => 
                           DP_OP_456J3_131_2158_n23, S => C431_DATA4_11);
   DP_OP_456J3_131_2158_U30 : HA_X1 port map( A => DP_OP_456J3_131_2158_n23, B 
                           => DP_OP_456J3_131_2158_n77, CO => 
                           DP_OP_456J3_131_2158_n22, S => C431_DATA4_12);
   DP_OP_456J3_131_2158_U29 : HA_X1 port map( A => DP_OP_456J3_131_2158_n22, B 
                           => DP_OP_456J3_131_2158_n78, CO => 
                           DP_OP_456J3_131_2158_n21, S => C431_DATA4_13);
   DP_OP_456J3_131_2158_U28 : HA_X1 port map( A => DP_OP_456J3_131_2158_n21, B 
                           => DP_OP_456J3_131_2158_n79, CO => 
                           DP_OP_456J3_131_2158_n20, S => C431_DATA4_14);
   DP_OP_456J3_131_2158_U27 : HA_X1 port map( A => DP_OP_456J3_131_2158_n20, B 
                           => DP_OP_456J3_131_2158_n80, CO => 
                           DP_OP_456J3_131_2158_n19, S => C431_DATA4_15);
   DP_OP_456J3_131_2158_U26 : HA_X1 port map( A => DP_OP_456J3_131_2158_n19, B 
                           => DP_OP_456J3_131_2158_n81, CO => 
                           DP_OP_456J3_131_2158_n18, S => C431_DATA4_16);
   DP_OP_456J3_131_2158_U25 : HA_X1 port map( A => DP_OP_456J3_131_2158_n18, B 
                           => DP_OP_456J3_131_2158_n82, CO => 
                           DP_OP_456J3_131_2158_n17, S => C431_DATA4_17);
   intadd_0_U28 : FA_X1 port map( A => intadd_0_A_0_port, B => 
                           intadd_0_B_0_port, CI => intadd_0_CI, CO => 
                           intadd_0_n27, S => intadd_0_SUM_0_port);
   intadd_0_U27 : FA_X1 port map( A => intadd_0_A_1_port, B => 
                           intadd_0_B_1_port, CI => intadd_0_n27, CO => 
                           intadd_0_n26, S => intadd_0_SUM_1_port);
   intadd_0_U26 : FA_X1 port map( A => intadd_0_A_2_port, B => 
                           intadd_0_B_2_port, CI => intadd_0_n26, CO => 
                           intadd_0_n25, S => intadd_0_SUM_2_port);
   intadd_0_U25 : FA_X1 port map( A => intadd_0_A_3_port, B => 
                           intadd_0_B_3_port, CI => intadd_0_n25, CO => 
                           intadd_0_n24, S => intadd_0_SUM_3_port);
   intadd_0_U24 : FA_X1 port map( A => intadd_0_A_4_port, B => 
                           intadd_0_B_4_port, CI => intadd_0_n24, CO => 
                           intadd_0_n23, S => intadd_0_SUM_4_port);
   intadd_0_U23 : FA_X1 port map( A => intadd_0_A_5_port, B => 
                           intadd_0_B_5_port, CI => intadd_0_n23, CO => 
                           intadd_0_n22, S => intadd_0_SUM_5_port);
   intadd_0_U22 : FA_X1 port map( A => intadd_0_A_6_port, B => 
                           intadd_0_B_6_port, CI => intadd_0_n22, CO => 
                           intadd_0_n21, S => intadd_0_SUM_6_port);
   intadd_0_U21 : FA_X1 port map( A => intadd_0_A_7_port, B => 
                           intadd_0_B_7_port, CI => intadd_0_n21, CO => 
                           intadd_0_n20, S => intadd_0_SUM_7_port);
   intadd_0_U20 : FA_X1 port map( A => intadd_0_A_8_port, B => 
                           intadd_0_B_8_port, CI => intadd_0_n20, CO => 
                           intadd_0_n19, S => intadd_0_SUM_8_port);
   intadd_0_U19 : FA_X1 port map( A => intadd_0_A_9_port, B => 
                           intadd_0_B_9_port, CI => intadd_0_n19, CO => 
                           intadd_0_n18, S => intadd_0_SUM_9_port);
   intadd_0_U18 : FA_X1 port map( A => intadd_0_A_10_port, B => 
                           intadd_0_B_10_port, CI => intadd_0_n18, CO => 
                           intadd_0_n17, S => intadd_0_SUM_10_port);
   intadd_0_U17 : FA_X1 port map( A => intadd_0_A_11_port, B => 
                           intadd_0_B_11_port, CI => intadd_0_n17, CO => 
                           intadd_0_n16, S => intadd_0_SUM_11_port);
   intadd_0_U16 : FA_X1 port map( A => intadd_0_A_12_port, B => 
                           intadd_0_B_12_port, CI => intadd_0_n16, CO => 
                           intadd_0_n15, S => intadd_0_SUM_12_port);
   intadd_0_U15 : FA_X1 port map( A => intadd_0_A_16_port, B => 
                           intadd_0_B_13_port, CI => intadd_0_n15, CO => 
                           intadd_0_n14, S => intadd_0_SUM_13_port);
   intadd_0_U14 : FA_X1 port map( A => intadd_0_A_16_port, B => 
                           intadd_0_B_14_port, CI => intadd_0_n14, CO => 
                           intadd_0_n13, S => intadd_0_SUM_14_port);
   intadd_0_U13 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n13, CO => intadd_0_n12, S => 
                           intadd_0_SUM_15_port);
   intadd_0_U12 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n12, CO => intadd_0_n11, S => 
                           intadd_0_SUM_16_port);
   intadd_0_U11 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n11, CO => intadd_0_n10, S => 
                           intadd_0_SUM_17_port);
   intadd_0_U10 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n10, CO => intadd_0_n9, S => 
                           intadd_0_SUM_18_port);
   intadd_0_U9 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n9, CO => intadd_0_n8, S => 
                           intadd_0_SUM_19_port);
   intadd_0_U8 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n8, CO => intadd_0_n7, S => 
                           intadd_0_SUM_20_port);
   intadd_0_U7 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n7, CO => intadd_0_n6, S => 
                           intadd_0_SUM_21_port);
   intadd_0_U6 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n6, CO => intadd_0_n5, S => 
                           intadd_0_SUM_22_port);
   intadd_0_U5 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n5, CO => intadd_0_n4, S => 
                           intadd_0_SUM_23_port);
   intadd_0_U4 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n4, CO => intadd_0_n3, S => 
                           intadd_0_SUM_24_port);
   intadd_0_U3 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n3, CO => intadd_0_n2, S => 
                           intadd_0_SUM_25_port);
   intadd_0_U2 : FA_X1 port map( A => intadd_0_A_16_port, B => n61, CI => 
                           intadd_0_n2, CO => intadd_0_n1, S => 
                           intadd_0_SUM_26_port);
   intadd_1_U26 : FA_X1 port map( A => intadd_1_A_0_port, B => 
                           intadd_1_B_0_port, CI => intadd_0_SUM_2_port, CO => 
                           intadd_1_n25, S => intadd_1_SUM_0_port);
   intadd_1_U25 : FA_X1 port map( A => intadd_0_SUM_3_port, B => 
                           intadd_1_B_1_port, CI => intadd_1_n25, CO => 
                           intadd_1_n24, S => intadd_1_SUM_1_port);
   intadd_1_U24 : FA_X1 port map( A => intadd_0_SUM_4_port, B => 
                           intadd_1_B_2_port, CI => intadd_1_n24, CO => 
                           intadd_1_n23, S => intadd_1_SUM_2_port);
   intadd_1_U23 : FA_X1 port map( A => intadd_0_SUM_5_port, B => 
                           intadd_1_B_3_port, CI => intadd_1_n23, CO => 
                           intadd_1_n22, S => intadd_1_SUM_3_port);
   intadd_1_U22 : FA_X1 port map( A => intadd_0_SUM_6_port, B => 
                           intadd_1_B_4_port, CI => intadd_1_n22, CO => 
                           intadd_1_n21, S => intadd_1_SUM_4_port);
   intadd_1_U21 : FA_X1 port map( A => intadd_0_SUM_7_port, B => 
                           intadd_1_B_5_port, CI => intadd_1_n21, CO => 
                           intadd_1_n20, S => intadd_1_SUM_5_port);
   intadd_1_U20 : FA_X1 port map( A => intadd_0_SUM_8_port, B => 
                           intadd_1_B_6_port, CI => intadd_1_n20, CO => 
                           intadd_1_n19, S => intadd_1_SUM_6_port);
   intadd_1_U19 : FA_X1 port map( A => intadd_0_SUM_9_port, B => 
                           intadd_1_B_7_port, CI => intadd_1_n19, CO => 
                           intadd_1_n18, S => intadd_1_SUM_7_port);
   intadd_1_U18 : FA_X1 port map( A => intadd_0_SUM_10_port, B => 
                           intadd_1_B_8_port, CI => intadd_1_n18, CO => 
                           intadd_1_n17, S => intadd_1_SUM_8_port);
   intadd_1_U17 : FA_X1 port map( A => intadd_0_SUM_11_port, B => 
                           intadd_1_B_9_port, CI => intadd_1_n17, CO => 
                           intadd_1_n16, S => intadd_1_SUM_9_port);
   intadd_1_U16 : FA_X1 port map( A => intadd_0_SUM_12_port, B => 
                           intadd_1_B_10_port, CI => intadd_1_n16, CO => 
                           intadd_1_n15, S => intadd_1_SUM_10_port);
   intadd_1_U15 : FA_X1 port map( A => intadd_0_SUM_13_port, B => 
                           intadd_1_B_11_port, CI => intadd_1_n15, CO => 
                           intadd_1_n14, S => intadd_1_SUM_11_port);
   intadd_1_U14 : FA_X1 port map( A => intadd_0_SUM_14_port, B => 
                           intadd_1_B_12_port, CI => intadd_1_n14, CO => 
                           intadd_1_n13, S => intadd_1_SUM_12_port);
   intadd_1_U13 : FA_X1 port map( A => intadd_0_SUM_15_port, B => 
                           intadd_1_B_13_port, CI => intadd_1_n13, CO => 
                           intadd_1_n12, S => intadd_1_SUM_13_port);
   intadd_1_U12 : FA_X1 port map( A => intadd_0_SUM_16_port, B => 
                           intadd_1_B_14_port, CI => intadd_1_n12, CO => 
                           intadd_1_n11, S => intadd_1_SUM_14_port);
   intadd_1_U11 : FA_X1 port map( A => intadd_0_SUM_17_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n11, CO => 
                           intadd_1_n10, S => intadd_1_SUM_15_port);
   intadd_1_U10 : FA_X1 port map( A => intadd_0_SUM_18_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n10, CO => 
                           intadd_1_n9, S => intadd_1_SUM_16_port);
   intadd_1_U9 : FA_X1 port map( A => intadd_0_SUM_19_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n9, CO => 
                           intadd_1_n8, S => intadd_1_SUM_17_port);
   intadd_1_U8 : FA_X1 port map( A => intadd_0_SUM_20_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n8, CO => 
                           intadd_1_n7, S => intadd_1_SUM_18_port);
   intadd_1_U7 : FA_X1 port map( A => intadd_0_SUM_21_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n7, CO => 
                           intadd_1_n6, S => intadd_1_SUM_19_port);
   intadd_1_U6 : FA_X1 port map( A => intadd_0_SUM_22_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n6, CO => 
                           intadd_1_n5, S => intadd_1_SUM_20_port);
   intadd_1_U5 : FA_X1 port map( A => intadd_0_SUM_23_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n5, CO => 
                           intadd_1_n4, S => intadd_1_SUM_21_port);
   intadd_1_U4 : FA_X1 port map( A => intadd_0_SUM_24_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n4, CO => 
                           intadd_1_n3, S => intadd_1_SUM_22_port);
   intadd_1_U3 : FA_X1 port map( A => intadd_0_SUM_25_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n3, CO => 
                           intadd_1_n2, S => intadd_1_SUM_23_port);
   intadd_1_U2 : FA_X1 port map( A => intadd_0_SUM_26_port, B => 
                           intadd_1_B_18_port, CI => intadd_1_n2, CO => 
                           intadd_1_n1, S => intadd_1_SUM_24_port);
   intadd_2_U11 : FA_X1 port map( A => intadd_2_A_0_port, B => 
                           intadd_2_B_0_port, CI => intadd_1_SUM_2_port, CO => 
                           intadd_2_n10, S => intadd_2_SUM_0_port);
   intadd_2_U10 : FA_X1 port map( A => intadd_2_A_1_port, B => 
                           intadd_1_SUM_3_port, CI => intadd_2_n10, CO => 
                           intadd_2_n9, S => intadd_2_SUM_1_port);
   intadd_2_U9 : FA_X1 port map( A => intadd_2_A_2_port, B => 
                           intadd_1_SUM_4_port, CI => intadd_2_n9, CO => 
                           intadd_2_n8, S => intadd_2_SUM_2_port);
   intadd_2_U8 : FA_X1 port map( A => intadd_2_A_3_port, B => 
                           intadd_1_SUM_5_port, CI => intadd_2_n8, CO => 
                           intadd_2_n7, S => intadd_2_SUM_3_port);
   intadd_2_U7 : FA_X1 port map( A => intadd_2_A_4_port, B => 
                           intadd_1_SUM_6_port, CI => intadd_2_n7, CO => 
                           intadd_2_n6, S => intadd_2_SUM_4_port);
   intadd_2_U6 : FA_X1 port map( A => intadd_2_A_5_port, B => 
                           intadd_1_SUM_7_port, CI => intadd_2_n6, CO => 
                           intadd_2_n5, S => intadd_2_SUM_5_port);
   intadd_2_U5 : FA_X1 port map( A => intadd_2_A_6_port, B => 
                           intadd_1_SUM_8_port, CI => intadd_2_n5, CO => 
                           intadd_2_n4, S => intadd_2_SUM_6_port);
   intadd_2_U4 : FA_X1 port map( A => intadd_2_A_7_port, B => 
                           intadd_1_SUM_9_port, CI => intadd_2_n4, CO => 
                           intadd_2_n3, S => intadd_2_SUM_7_port);
   intadd_2_U3 : FA_X1 port map( A => intadd_2_A_8_port, B => 
                           intadd_1_SUM_10_port, CI => intadd_2_n3, CO => 
                           intadd_2_n2, S => intadd_2_SUM_8_port);
   intadd_2_U2 : FA_X1 port map( A => intadd_2_A_9_port, B => 
                           intadd_1_SUM_11_port, CI => intadd_2_n2, CO => 
                           intadd_2_n1, S => intadd_2_SUM_9_port);
   OP_A_reg_7_inst : DLH_X1 port map( G => N246, D => OP1(7), Q => OP_A_7_port)
                           ;
   OP_A_reg_12_inst : DLH_X1 port map( G => N246, D => OP1(12), Q => 
                           OP_A_12_port);
   OP_A_reg_13_inst : DLH_X1 port map( G => n1412, D => OP1(13), Q => 
                           OP_A_13_port);
   OP_A_reg_10_inst : DLH_X1 port map( G => n1412, D => OP1(10), Q => 
                           OP_A_10_port);
   OP_A_reg_0_inst : DLH_X1 port map( G => n1412, D => OP1(0), Q => OP_A_0_port
                           );
   OP_A_reg_4_inst : DLH_X1 port map( G => N246, D => OP1(4), Q => OP_A_4_port)
                           ;
   OP_A_reg_8_inst : DLH_X1 port map( G => n1412, D => OP1(8), Q => OP_A_8_port
                           );
   OP_A_reg_6_inst : DLH_X1 port map( G => N246, D => OP1(6), Q => OP_A_6_port)
                           ;
   OP_A_reg_11_inst : DLH_X1 port map( G => n1412, D => OP1(11), Q => 
                           OP_A_11_port);
   OP_A_reg_14_inst : DLH_X1 port map( G => n1412, D => OP1(14), Q => 
                           OP_A_14_port);
   OP_A_reg_1_inst : DLH_X1 port map( G => N246, D => OP1(1), Q => OP_A_1_port)
                           ;
   OP_A_reg_3_inst : DLH_X1 port map( G => N246, D => OP1(3), Q => OP_A_3_port)
                           ;
   OP_A_reg_9_inst : DLH_X1 port map( G => n1412, D => OP1(9), Q => OP_A_9_port
                           );
   OP_A_reg_5_inst : DLH_X1 port map( G => n1412, D => OP1(5), Q => OP_A_5_port
                           );
   OP_B_reg_2_inst : DLH_X1 port map( G => N246, D => N249, Q => OP_B_2_port);
   OP_B_reg_5_inst : DLH_X1 port map( G => n1412, D => N252, Q => OP_B_5_port);
   OP_B_reg_3_inst : DLH_X1 port map( G => N246, D => N250, Q => OP_B_3_port);
   OP_A_reg_15_inst : DLH_X1 port map( G => n1412, D => OP1(15), Q => 
                           OP_A_15_port);
   OP_B_reg_4_inst : DLH_X1 port map( G => N246, D => N251, Q => OP_B_4_port);
   OP_A_reg_2_inst : DLH_X1 port map( G => N246, D => OP1(2), Q => OP_A_2_port)
                           ;
   OP_B_reg_1_inst : DLH_X2 port map( G => N246, D => N248, Q => OP_B_1_port);
   U3 : CLKBUF_X1 port map( A => n148, Z => n59);
   U4 : INV_X2 port map( A => n577, ZN => n55);
   U5 : INV_X2 port map( A => n607, ZN => n56);
   U6 : INV_X1 port map( A => n1368, ZN => n1367);
   U7 : INV_X1 port map( A => n1245, ZN => n1369);
   U8 : INV_X1 port map( A => n1372, ZN => n1344);
   U9 : INV_X2 port map( A => N280, ZN => n195);
   U10 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_15, B1 => 
                           OP_A_11_port, B2 => n159, C1 => n160, C2 => 
                           OP_A_10_port, ZN => intadd_1_B_9_port);
   U11 : AOI211_X1 port map( C1 => n63, C2 => n863, A => n540, B => n539, ZN =>
                           n964);
   U12 : OR3_X1 port map( A1 => n1081, A2 => OP_B_7_port, A3 => n161, ZN => n57
                           );
   U13 : OR2_X1 port map( A1 => n145, A2 => n114, ZN => n58);
   U14 : NOR2_X2 port map( A1 => OP_B_2_port, A2 => n1160, ZN => n855);
   U15 : NOR2_X2 port map( A1 => OP_B_7_port, A2 => n162, ZN => n1027);
   U16 : NOR2_X2 port map( A1 => n223, A2 => n742, ZN => n147);
   U17 : NOR2_X2 port map( A1 => OP_B_5_port, A2 => n154, ZN => n160);
   U18 : AOI21_X2 port map( B1 => OP_B_3_port, B2 => OP_B_4_port, A => n296, ZN
                           => n1413);
   U19 : NOR2_X2 port map( A1 => OP_B_3_port, A2 => OP_B_2_port, ZN => n894);
   U20 : INV_X1 port map( A => n57, ZN => n60);
   U21 : INV_X1 port map( A => n58, ZN => n61);
   U22 : NOR2_X2 port map( A1 => n900, A2 => n1261, ZN => n1228);
   U23 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n581, ZN => n62);
   U24 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n581, ZN => n63);
   U25 : NOR2_X2 port map( A1 => n1381, A2 => n111, ZN => intadd_1_B_18_port);
   U26 : AOI21_X2 port map( B1 => OP_B_2_port, B2 => OP_B_1_port, A => n1160, 
                           ZN => n1415);
   U27 : NOR3_X4 port map( A1 => n150, A2 => OP_B_5_port, A3 => n153, ZN => 
                           n159);
   U28 : NOR2_X4 port map( A1 => n126, A2 => n109, ZN => intadd_0_A_16_port);
   U29 : NOR3_X4 port map( A1 => n1081, A2 => OP_B_7_port, A3 => n1080, ZN => 
                           n1380);
   U30 : OR2_X1 port map( A1 => n1413, A2 => n1381, ZN => n64);
   U31 : NOR2_X2 port map( A1 => DP_OP_446J3_125_4819_n12, A2 => n1092, ZN => 
                           n65);
   U32 : INV_X1 port map( A => OPC(4), ZN => n69);
   U33 : NOR2_X1 port map( A1 => OPC(2), A2 => OPC(1), ZN => n72);
   U34 : INV_X1 port map( A => OPC(6), ZN => n170);
   U35 : NOR3_X1 port map( A1 => OPC(5), A2 => n69, A3 => n170, ZN => n80);
   U36 : NAND2_X1 port map( A1 => OPC(4), A2 => OPC(5), ZN => n81);
   U37 : NOR2_X1 port map( A1 => OPC(6), A2 => n81, ZN => n77);
   U38 : NOR2_X1 port map( A1 => n80, A2 => n77, ZN => n175);
   U39 : INV_X1 port map( A => OPC(3), ZN => n66);
   U40 : INV_X1 port map( A => OPC(0), ZN => n67);
   U41 : NAND3_X1 port map( A1 => n72, A2 => n66, A3 => n67, ZN => n96_port);
   U42 : INV_X1 port map( A => OPC(5), ZN => n68);
   U43 : NAND2_X1 port map( A1 => n69, A2 => n68, ZN => n215);
   U44 : NOR2_X1 port map( A1 => OPC(3), A2 => n67, ZN => n83);
   U45 : NAND2_X1 port map( A1 => n72, A2 => n83, ZN => n1411);
   U46 : OAI22_X1 port map( A1 => n175, A2 => n96_port, B1 => n215, B2 => n1411
                           , ZN => N280);
   U47 : NOR2_X1 port map( A1 => OPC(4), A2 => n68, ZN => n88);
   U48 : NAND2_X1 port map( A1 => n88, A2 => n170, ZN => n171);
   U49 : NOR3_X1 port map( A1 => OPC(6), A2 => OPC(5), A3 => n69, ZN => n100);
   U50 : INV_X1 port map( A => n100, ZN => n1410);
   U51 : NAND3_X1 port map( A1 => OPC(3), A2 => OPC(0), A3 => n72, ZN => n214);
   U52 : OAI22_X1 port map( A1 => n171, A2 => n96_port, B1 => n1410, B2 => n214
                           , ZN => N96);
   U53 : NAND3_X1 port map( A1 => OPC(6), A2 => OPC(5), A3 => n69, ZN => n1406)
                           ;
   U54 : INV_X1 port map( A => n96_port, ZN => n102);
   U55 : INV_X1 port map( A => n215, ZN => n101);
   U56 : NAND2_X1 port map( A1 => OPC(6), A2 => n101, ZN => n1409);
   U57 : INV_X1 port map( A => n1409, ZN => n70);
   U58 : AOI21_X1 port map( B1 => n102, B2 => n70, A => N96, ZN => n71);
   U59 : OAI21_X1 port map( B1 => n1406, B2 => n214, A => n71, ZN => N284);
   U60 : NAND2_X1 port map( A1 => OPC(3), A2 => n72, ZN => n73);
   U61 : NOR2_X1 port map( A1 => OPC(0), A2 => n73, ZN => n86);
   U62 : INV_X1 port map( A => n86, ZN => n1408);
   U63 : INV_X1 port map( A => n214, ZN => n78);
   U64 : NAND2_X1 port map( A1 => OPC(2), A2 => OPC(3), ZN => n74);
   U65 : NOR2_X1 port map( A1 => OPC(0), A2 => n74, ZN => n94);
   U66 : INV_X1 port map( A => OPC(1), ZN => n104);
   U67 : INV_X1 port map( A => OPC(2), ZN => n75);
   U68 : NAND3_X1 port map( A1 => OPC(1), A2 => n83, A3 => n75, ZN => n93);
   U69 : INV_X1 port map( A => n93, ZN => n76);
   U70 : AOI21_X1 port map( B1 => n94, B2 => n104, A => n76, ZN => n178);
   U71 : NOR2_X1 port map( A1 => OPC(4), A2 => n178, ZN => n168);
   U72 : AOI21_X1 port map( B1 => n78, B2 => n77, A => n168, ZN => n79);
   U73 : OAI21_X1 port map( B1 => n1406, B2 => n1408, A => n79, ZN => N286);
   U74 : INV_X1 port map( A => n80, ZN => n216);
   U75 : AOI21_X1 port map( B1 => n171, B2 => n216, A => n1408, ZN => n84);
   U76 : NAND2_X1 port map( A1 => OPC(4), A2 => n170, ZN => n82);
   U77 : OR2_X1 port map( A1 => n170, A2 => n81, ZN => n90);
   U78 : OAI22_X1 port map( A1 => n82, A2 => n1408, B1 => n214, B2 => n90, ZN 
                           => n167);
   U79 : NAND3_X1 port map( A1 => OPC(2), A2 => n83, A3 => n104, ZN => n92);
   U80 : OAI22_X1 port map( A1 => n171, A2 => n92, B1 => n1408, B2 => n90, ZN 
                           => n176);
   U81 : NOR4_X1 port map( A1 => n84, A2 => n167, A3 => N286, A4 => n176, ZN =>
                           n85);
   U82 : OR2_X1 port map( A1 => n215, A2 => n92, ZN => n173);
   U83 : OAI211_X1 port map( C1 => n214, C2 => n216, A => n85, B => n173, ZN =>
                           N285);
   U84 : NAND2_X1 port map( A1 => n101, A2 => n86, ZN => n1407);
   U85 : INV_X1 port map( A => n1411, ZN => n87);
   U86 : OAI21_X1 port map( B1 => n88, B2 => n100, A => n87, ZN => n89);
   U87 : OAI211_X1 port map( C1 => n96_port, C2 => n90, A => n1407, B => n89, 
                           ZN => N281);
   U88 : NAND3_X1 port map( A1 => OPC(2), A2 => OPC(3), A3 => OPC(0), ZN => n91
                           );
   U89 : OAI211_X1 port map( C1 => OPC(1), C2 => n91, A => n93, B => n96_port, 
                           ZN => n99);
   U90 : AOI21_X1 port map( B1 => n93, B2 => n92, A => n216, ZN => n98);
   U91 : NAND3_X1 port map( A1 => OPC(5), A2 => OPC(1), A3 => n94, ZN => n95);
   U92 : OAI21_X1 port map( B1 => n96_port, B2 => n1406, A => n95, ZN => n97);
   U93 : AOI211_X1 port map( C1 => n100, C2 => n99, A => n98, B => n97, ZN => 
                           n115);
   U94 : INV_X1 port map( A => N281, ZN => n218);
   U95 : NAND3_X1 port map( A1 => n102, A2 => n101, A3 => n170, ZN => n103);
   U96 : OAI21_X1 port map( B1 => n214, B2 => n171, A => n103, ZN => n1366);
   U97 : INV_X1 port map( A => n1366, ZN => n900);
   U98 : INV_X1 port map( A => n171, ZN => n106);
   U99 : AOI211_X1 port map( C1 => OPC(3), C2 => OPC(2), A => OPC(0), B => n104
                           , ZN => n105);
   U100 : OAI211_X1 port map( C1 => OPC(2), C2 => OPC(3), A => n106, B => n105,
                           ZN => n1396);
   U101 : NAND4_X1 port map( A1 => n115, A2 => n218, A3 => n900, A4 => n1396, 
                           ZN => n107);
   U102 : NOR3_X2 port map( A1 => N284, A2 => N285, A3 => n107, ZN => n193);
   U103 : CLKBUF_X1 port map( A => n193, Z => n204);
   U104 : NAND2_X1 port map( A1 => n195, A2 => n204, ZN => N246);
   U105 : CLKBUF_X1 port map( A => N246, Z => n1412);
   U106 : INV_X1 port map( A => OP_A_15_port, ZN => n1080);
   U107 : INV_X1 port map( A => OP_B_1_port, ZN => n223);
   U108 : INV_X1 port map( A => OP_B_0_port, ZN => n222);
   U109 : OR2_X1 port map( A1 => OP_B_1_port, A2 => n222, ZN => n509);
   U110 : NOR2_X1 port map( A1 => n1080, A2 => n509, ZN => n126);
   U111 : NOR2_X1 port map( A1 => OP_B_0_port, A2 => n223, ZN => n603);
   U112 : INV_X1 port map( A => n603, ZN => n575);
   U113 : OR2_X1 port map( A1 => n223, A2 => n222, ZN => n577);
   U114 : NAND2_X1 port map( A1 => n55, A2 => n1080, ZN => n116);
   U115 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n575, A => n116, ZN => 
                           n108);
   U116 : INV_X1 port map( A => n108, ZN => n123);
   U117 : NOR2_X1 port map( A1 => DP_OP_440J3_122_9847_n20, A2 => n123, ZN => 
                           n109);
   U118 : INV_X1 port map( A => OP_B_7_port, ZN => n294);
   U119 : AOI21_X1 port map( B1 => OP_B_6_port, B2 => OP_B_5_port, A => n294, 
                           ZN => n1414);
   U120 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => OP_B_3_port, ZN => n150);
   U121 : NOR3_X1 port map( A1 => n150, A2 => OP_B_5_port, A3 => n1080, ZN => 
                           n1381);
   U122 : NAND2_X1 port map( A1 => n150, A2 => OP_B_5_port, ZN => n121);
   U123 : INV_X1 port map( A => OP_B_3_port, ZN => n1160);
   U124 : INV_X1 port map( A => OP_B_4_port, ZN => n1363);
   U125 : NOR2_X1 port map( A1 => n1160, A2 => n1363, ZN => n153);
   U126 : INV_X1 port map( A => OP_B_5_port, ZN => n296);
   U127 : NOR3_X1 port map( A1 => n150, A2 => n153, A3 => n296, ZN => n151);
   U128 : NAND2_X1 port map( A1 => n151, A2 => n1080, ZN => n120);
   U129 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n121, A => n120, ZN => 
                           n110);
   U130 : INV_X1 port map( A => n110, ZN => n157);
   U131 : OR2_X1 port map( A1 => DP_OP_451J3_128_3502_n15, A2 => n157, ZN => 
                           n1383);
   U132 : INV_X1 port map( A => n1383, ZN => n111);
   U133 : INV_X1 port map( A => OP_B_2_port, ZN => n581);
   U134 : AOI211_X1 port map( C1 => n581, C2 => n223, A => OP_B_3_port, B => 
                           n1080, ZN => n145);
   U135 : NAND2_X1 port map( A1 => n855, A2 => n223, ZN => n118);
   U136 : NAND2_X1 port map( A1 => OP_B_3_port, A2 => OP_B_2_port, ZN => n857);
   U137 : NAND2_X1 port map( A1 => OP_B_1_port, A2 => n855, ZN => n112);
   U138 : OAI21_X1 port map( B1 => OP_B_1_port, B2 => n857, A => n112, ZN => 
                           n137);
   U139 : NAND2_X1 port map( A1 => n1080, A2 => n137, ZN => n117);
   U140 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n118, A => n117, ZN => 
                           n113);
   U141 : INV_X1 port map( A => n113, ZN => n142);
   U142 : NOR2_X1 port map( A1 => DP_OP_456J3_131_2158_n17, A2 => n142, ZN => 
                           n114);
   U143 : NAND2_X1 port map( A1 => n195, A2 => n115, ZN => N279);
   U144 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n575, A => n116, ZN => 
                           DP_OP_440J3_122_9847_n80);
   U145 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n577, B1 => OP_A_13_port
                           , B2 => n575, ZN => DP_OP_440J3_122_9847_n79);
   U146 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n577, B1 => OP_A_12_port
                           , B2 => n575, ZN => DP_OP_440J3_122_9847_n78);
   U147 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n575, B1 => OP_A_12_port
                           , B2 => n577, ZN => DP_OP_440J3_122_9847_n77);
   U148 : OAI22_X1 port map( A1 => OP_A_10_port, A2 => n575, B1 => OP_A_11_port
                           , B2 => n577, ZN => DP_OP_440J3_122_9847_n76);
   U149 : OAI22_X1 port map( A1 => OP_A_9_port, A2 => n575, B1 => OP_A_10_port,
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n75);
   U150 : OAI22_X1 port map( A1 => OP_A_8_port, A2 => n575, B1 => OP_A_9_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n74);
   U151 : OAI22_X1 port map( A1 => OP_A_7_port, A2 => n575, B1 => OP_A_8_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n73);
   U152 : OAI22_X1 port map( A1 => OP_A_6_port, A2 => n575, B1 => OP_A_7_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n72);
   U153 : OAI22_X1 port map( A1 => OP_A_5_port, A2 => n575, B1 => OP_A_6_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n71);
   U154 : OAI22_X1 port map( A1 => OP_A_4_port, A2 => n575, B1 => OP_A_5_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n70);
   U155 : OAI22_X1 port map( A1 => OP_A_3_port, A2 => n575, B1 => OP_A_4_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n69);
   U156 : OAI22_X1 port map( A1 => OP_A_2_port, A2 => n575, B1 => OP_A_3_port, 
                           B2 => n577, ZN => DP_OP_440J3_122_9847_n68);
   U157 : OAI22_X1 port map( A1 => OP_A_2_port, A2 => n577, B1 => OP_A_1_port, 
                           B2 => n575, ZN => DP_OP_440J3_122_9847_n67);
   U158 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n577, B1 => OP_A_0_port, 
                           B2 => n575, ZN => DP_OP_440J3_122_9847_n66);
   U159 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n577, A => n575, ZN => 
                           DP_OP_440J3_122_9847_n35);
   U160 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n118, A => n117, ZN => 
                           DP_OP_456J3_131_2158_n82);
   U161 : INV_X1 port map( A => n137, ZN => n119);
   U162 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n119, B1 => OP_A_13_port
                           , B2 => n118, ZN => DP_OP_456J3_131_2158_n81);
   U163 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n119, B1 => OP_A_12_port
                           , B2 => n118, ZN => DP_OP_456J3_131_2158_n80);
   U164 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n118, B1 => OP_A_12_port
                           , B2 => n119, ZN => DP_OP_456J3_131_2158_n79);
   U165 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n119, B1 => OP_A_10_port
                           , B2 => n118, ZN => DP_OP_456J3_131_2158_n78);
   U166 : OAI22_X1 port map( A1 => n119, A2 => OP_A_10_port, B1 => OP_A_9_port,
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n77);
   U167 : OAI22_X1 port map( A1 => n119, A2 => OP_A_9_port, B1 => OP_A_8_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n76);
   U168 : OAI22_X1 port map( A1 => n119, A2 => OP_A_8_port, B1 => OP_A_7_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n75);
   U169 : OAI22_X1 port map( A1 => n119, A2 => OP_A_7_port, B1 => OP_A_6_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n74);
   U170 : OAI22_X1 port map( A1 => n119, A2 => OP_A_6_port, B1 => OP_A_5_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n73);
   U171 : OAI22_X1 port map( A1 => n119, A2 => OP_A_5_port, B1 => OP_A_4_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n72);
   U172 : OAI22_X1 port map( A1 => n119, A2 => OP_A_4_port, B1 => OP_A_3_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n71);
   U173 : OAI22_X1 port map( A1 => n119, A2 => OP_A_3_port, B1 => OP_A_2_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n70);
   U174 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n118, B1 => n119, B2 => 
                           OP_A_2_port, ZN => DP_OP_456J3_131_2158_n69);
   U175 : OAI22_X1 port map( A1 => n119, A2 => OP_A_1_port, B1 => OP_A_0_port, 
                           B2 => n118, ZN => DP_OP_456J3_131_2158_n68);
   U176 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n119, A => n118, ZN => 
                           DP_OP_456J3_131_2158_n67);
   U177 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n121, A => n120, ZN => 
                           DP_OP_451J3_128_3502_n85);
   U178 : INV_X1 port map( A => n151, ZN => n122);
   U179 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n122, B1 => OP_A_13_port
                           , B2 => n121, ZN => DP_OP_451J3_128_3502_n84);
   U180 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n122, B1 => OP_A_12_port
                           , B2 => n121, ZN => DP_OP_451J3_128_3502_n83);
   U181 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n121, B1 => OP_A_12_port
                           , B2 => n122, ZN => DP_OP_451J3_128_3502_n82);
   U182 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n122, B1 => OP_A_10_port
                           , B2 => n121, ZN => DP_OP_451J3_128_3502_n81);
   U183 : OAI22_X1 port map( A1 => OP_A_10_port, A2 => n122, B1 => OP_A_9_port,
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n80);
   U184 : OAI22_X1 port map( A1 => OP_A_9_port, A2 => n122, B1 => OP_A_8_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n79);
   U185 : OAI22_X1 port map( A1 => OP_A_8_port, A2 => n122, B1 => OP_A_7_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n78);
   U186 : OAI22_X1 port map( A1 => OP_A_7_port, A2 => n122, B1 => OP_A_6_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n77);
   U187 : OAI22_X1 port map( A1 => OP_A_6_port, A2 => n122, B1 => OP_A_5_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n76);
   U188 : OAI22_X1 port map( A1 => OP_A_5_port, A2 => n122, B1 => OP_A_4_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n75);
   U189 : OAI22_X1 port map( A1 => OP_A_4_port, A2 => n122, B1 => OP_A_3_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n74);
   U190 : OAI22_X1 port map( A1 => OP_A_3_port, A2 => n122, B1 => OP_A_2_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n73);
   U191 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n121, B1 => OP_A_2_port, 
                           B2 => n122, ZN => DP_OP_451J3_128_3502_n72);
   U192 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n122, B1 => OP_A_0_port, 
                           B2 => n121, ZN => DP_OP_451J3_128_3502_n71);
   U193 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n122, A => n121, ZN => 
                           DP_OP_451J3_128_3502_n70);
   U194 : XNOR2_X1 port map( A => DP_OP_440J3_122_9847_n20, B => n123, ZN => 
                           n124);
   U195 : INV_X1 port map( A => n126, ZN => n890);
   U196 : NAND2_X1 port map( A1 => n223, A2 => n890, ZN => n125);
   U197 : OAI21_X1 port map( B1 => n126, B2 => n124, A => n125, ZN => 
                           intadd_0_A_12_port);
   U198 : OAI21_X1 port map( B1 => n126, B2 => C428_DATA4_15, A => n125, ZN => 
                           intadd_0_A_11_port);
   U199 : INV_X1 port map( A => n509, ZN => n542);
   U200 : NAND2_X1 port map( A1 => n542, A2 => OP_A_14_port, ZN => n852);
   U201 : INV_X1 port map( A => n852, ZN => n127);
   U202 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_14, A => n127,
                           ZN => intadd_0_A_10_port);
   U203 : INV_X1 port map( A => n509, ZN => n491);
   U204 : NAND2_X1 port map( A1 => n491, A2 => OP_A_13_port, ZN => n819);
   U205 : INV_X1 port map( A => n819, ZN => n128);
   U206 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_13, A => n128,
                           ZN => intadd_0_A_9_port);
   U207 : NAND2_X1 port map( A1 => n542, A2 => OP_A_12_port, ZN => n804);
   U208 : INV_X1 port map( A => n804, ZN => n129);
   U209 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_12, A => n129,
                           ZN => intadd_0_A_8_port);
   U210 : NAND2_X1 port map( A1 => n542, A2 => OP_A_11_port, ZN => n769);
   U211 : INV_X1 port map( A => n769, ZN => n130);
   U212 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_11, A => n130,
                           ZN => intadd_0_A_7_port);
   U213 : NAND2_X1 port map( A1 => n542, A2 => OP_A_10_port, ZN => n740);
   U214 : INV_X1 port map( A => n740, ZN => n131);
   U215 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_10, A => n131,
                           ZN => intadd_0_A_6_port);
   U216 : NAND2_X1 port map( A1 => n491, A2 => OP_A_9_port, ZN => n726);
   U217 : INV_X1 port map( A => n726, ZN => n132);
   U218 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_9, A => n132, 
                           ZN => intadd_0_A_5_port);
   U219 : NAND2_X1 port map( A1 => n542, A2 => OP_A_8_port, ZN => n696);
   U220 : INV_X1 port map( A => n696, ZN => n133);
   U221 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_8, A => n133, 
                           ZN => intadd_0_A_4_port);
   U222 : NAND2_X1 port map( A1 => n542, A2 => OP_A_7_port, ZN => n675);
   U223 : INV_X1 port map( A => n675, ZN => n134);
   U224 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_7, A => n134, 
                           ZN => intadd_0_A_3_port);
   U225 : NAND2_X1 port map( A1 => n542, A2 => OP_A_6_port, ZN => n658);
   U226 : INV_X1 port map( A => n658, ZN => n135);
   U227 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_6, A => n135, 
                           ZN => intadd_0_A_2_port);
   U228 : NAND2_X1 port map( A1 => n491, A2 => OP_A_5_port, ZN => n628);
   U229 : INV_X1 port map( A => n628, ZN => n136);
   U230 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_5, A => n136, 
                           ZN => intadd_0_A_1_port);
   U231 : INV_X1 port map( A => n894, ZN => n765);
   U232 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n581, ZN => n853);
   U233 : INV_X1 port map( A => n853, ZN => n742);
   U234 : AOI22_X1 port map( A1 => OP_B_1_port, A2 => n765, B1 => n742, B2 => 
                           n223, ZN => n148);
   U235 : AND2_X1 port map( A1 => n137, A2 => C2_DATA1_2, ZN => n138);
   U236 : AOI21_X1 port map( B1 => n59, B2 => OP_A_0_port, A => n138, ZN => 
                           n525);
   U237 : INV_X1 port map( A => OP_A_2_port, ZN => n576);
   U238 : NOR2_X1 port map( A1 => n509, A2 => n576, ZN => n552);
   U239 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_2, A => n552, 
                           ZN => n526);
   U240 : NOR2_X1 port map( A1 => n525, A2 => n526, ZN => n537);
   U241 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_3, B1 => 
                           OP_A_0_port, B2 => n147, C1 => n59, C2 => 
                           OP_A_1_port, ZN => n140);
   U242 : INV_X1 port map( A => n140, ZN => n534);
   U243 : INV_X1 port map( A => n537, ZN => n139);
   U244 : INV_X1 port map( A => OP_A_3_port, ZN => n550);
   U245 : NOR2_X1 port map( A1 => n509, A2 => n550, ZN => n580);
   U246 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_3, A => n580, 
                           ZN => n535);
   U247 : OAI21_X1 port map( B1 => n140, B2 => n139, A => n535, ZN => n141);
   U248 : OAI21_X1 port map( B1 => n537, B2 => n534, A => n141, ZN => 
                           intadd_0_A_0_port);
   U249 : XNOR2_X1 port map( A => DP_OP_456J3_131_2158_n17, B => n142, ZN => 
                           n144);
   U250 : OR2_X1 port map( A1 => n145, A2 => n1415, ZN => n143);
   U251 : OAI21_X1 port map( B1 => n145, B2 => n144, A => n143, ZN => 
                           intadd_0_B_14_port);
   U252 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_17, B1 => 
                           OP_A_15_port, B2 => n59, C1 => OP_A_14_port, C2 => 
                           n147, ZN => intadd_0_B_13_port);
   U253 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_16, B1 => 
                           OP_A_13_port, B2 => n147, C1 => OP_A_14_port, C2 => 
                           n59, ZN => intadd_0_B_12_port);
   U254 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_15, B1 => 
                           OP_A_12_port, B2 => n147, C1 => OP_A_13_port, C2 => 
                           n59, ZN => intadd_0_B_11_port);
   U255 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_14, B1 => 
                           OP_A_12_port, B2 => n59, C1 => OP_A_11_port, C2 => 
                           n147, ZN => intadd_0_B_10_port);
   U256 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_13, B1 => 
                           OP_A_11_port, B2 => n59, C1 => n147, C2 => 
                           OP_A_10_port, ZN => intadd_0_B_9_port);
   U257 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_12, B1 => n59, B2 
                           => OP_A_10_port, C1 => n147, C2 => OP_A_9_port, ZN 
                           => intadd_0_B_8_port);
   U258 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_11, B1 => n59, B2 
                           => OP_A_9_port, C1 => n147, C2 => OP_A_8_port, ZN =>
                           intadd_0_B_7_port);
   U259 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_10, B1 => n59, B2 
                           => OP_A_8_port, C1 => n147, C2 => OP_A_7_port, ZN =>
                           intadd_0_B_6_port);
   U260 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_9, B1 => n59, B2 =>
                           OP_A_7_port, C1 => n147, C2 => OP_A_6_port, ZN => 
                           intadd_0_B_5_port);
   U261 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_8, B1 => n59, B2 =>
                           OP_A_6_port, C1 => n147, C2 => OP_A_5_port, ZN => 
                           intadd_0_B_4_port);
   U262 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_7, B1 => n59, B2 =>
                           OP_A_5_port, C1 => n147, C2 => OP_A_4_port, ZN => 
                           intadd_0_B_3_port);
   U263 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_6, B1 => n59, B2 =>
                           OP_A_4_port, C1 => n147, C2 => OP_A_3_port, ZN => 
                           intadd_0_B_2_port);
   U264 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_5, B1 => n59, B2 =>
                           OP_A_3_port, C1 => n147, C2 => OP_A_2_port, ZN => 
                           intadd_0_B_1_port);
   U265 : NAND2_X1 port map( A1 => n542, A2 => OP_A_4_port, ZN => n604);
   U266 : INV_X1 port map( A => n604, ZN => n146);
   U267 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_4, A => n146, 
                           ZN => intadd_0_B_0_port);
   U268 : AOI222_X1 port map( A1 => n1415, A2 => C431_DATA4_4, B1 => n59, B2 =>
                           OP_A_2_port, C1 => n147, C2 => OP_A_1_port, ZN => 
                           intadd_0_CI);
   U269 : NOR2_X1 port map( A1 => OP_B_5_port, A2 => OP_B_6_port, ZN => n1081);
   U270 : NAND2_X1 port map( A1 => n1081, A2 => OP_B_7_port, ZN => n1078);
   U271 : INV_X1 port map( A => OP_B_6_port, ZN => n377);
   U272 : NOR2_X1 port map( A1 => n296, A2 => n377, ZN => n161);
   U273 : NOR3_X1 port map( A1 => n1081, A2 => n161, A3 => n294, ZN => n163);
   U274 : NAND2_X1 port map( A1 => n163, A2 => n1080, ZN => n1077);
   U275 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => n1078, A => n1077, ZN =>
                           DP_OP_446J3_125_4819_n87);
   U276 : INV_X1 port map( A => n163, ZN => n149);
   U277 : OAI22_X1 port map( A1 => OP_A_14_port, A2 => n149, B1 => OP_A_13_port
                           , B2 => n1078, ZN => DP_OP_446J3_125_4819_n86);
   U278 : OAI22_X1 port map( A1 => OP_A_13_port, A2 => n149, B1 => OP_A_12_port
                           , B2 => n1078, ZN => DP_OP_446J3_125_4819_n85);
   U279 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n1078, B1 => 
                           OP_A_12_port, B2 => n149, ZN => 
                           DP_OP_446J3_125_4819_n84);
   U280 : OAI22_X1 port map( A1 => OP_A_11_port, A2 => n149, B1 => OP_A_10_port
                           , B2 => n1078, ZN => DP_OP_446J3_125_4819_n83);
   U281 : OAI22_X1 port map( A1 => OP_A_10_port, A2 => n149, B1 => OP_A_9_port,
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n82);
   U282 : OAI22_X1 port map( A1 => OP_A_9_port, A2 => n149, B1 => OP_A_8_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n81);
   U283 : OAI22_X1 port map( A1 => OP_A_8_port, A2 => n149, B1 => OP_A_7_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n80);
   U284 : OAI22_X1 port map( A1 => OP_A_7_port, A2 => n149, B1 => OP_A_6_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n79);
   U285 : OAI22_X1 port map( A1 => OP_A_6_port, A2 => n149, B1 => OP_A_5_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n78);
   U286 : OAI22_X1 port map( A1 => OP_A_5_port, A2 => n149, B1 => OP_A_4_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n77);
   U287 : OAI22_X1 port map( A1 => OP_A_4_port, A2 => n149, B1 => OP_A_3_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n76);
   U288 : OAI22_X1 port map( A1 => OP_A_3_port, A2 => n149, B1 => OP_A_2_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n75);
   U289 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n1078, B1 => OP_A_2_port,
                           B2 => n149, ZN => DP_OP_446J3_125_4819_n74);
   U290 : OAI22_X1 port map( A1 => OP_A_1_port, A2 => n149, B1 => OP_A_0_port, 
                           B2 => n1078, ZN => DP_OP_446J3_125_4819_n73);
   U291 : OAI21_X1 port map( B1 => OP_A_0_port, B2 => n149, A => n1078, ZN => 
                           DP_OP_446J3_125_4819_n72);
   U292 : AND2_X1 port map( A1 => C2_DATA1_4, A2 => n151, ZN => n152);
   U293 : AOI21_X1 port map( B1 => n159, B2 => OP_A_0_port, A => n152, ZN => 
                           n565);
   U294 : NOR2_X1 port map( A1 => intadd_0_SUM_0_port, A2 => n565, ZN => n564);
   U295 : INV_X1 port map( A => intadd_0_SUM_1_port, ZN => n156);
   U296 : INV_X1 port map( A => n564, ZN => n590);
   U297 : INV_X1 port map( A => n153, ZN => n154);
   U298 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_5, B1 => 
                           OP_A_0_port, B2 => n160, C1 => OP_A_1_port, C2 => 
                           n159, ZN => n591);
   U299 : OAI21_X1 port map( B1 => intadd_0_SUM_1_port, B2 => n590, A => n591, 
                           ZN => n155);
   U300 : OAI21_X1 port map( B1 => n564, B2 => n156, A => n155, ZN => 
                           intadd_1_A_0_port);
   U301 : XNOR2_X1 port map( A => DP_OP_451J3_128_3502_n15, B => n157, ZN => 
                           n158);
   U302 : OAI21_X1 port map( B1 => n1381, B2 => n158, A => n64, ZN => 
                           intadd_1_B_14_port);
   U303 : AOI222_X1 port map( A1 => OP_A_15_port, A2 => n159, B1 => n1413, B2 
                           => C430_DATA4_19, C1 => OP_A_14_port, C2 => n160, ZN
                           => intadd_1_B_13_port);
   U304 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_18, B1 => 
                           OP_A_13_port, B2 => n160, C1 => OP_A_14_port, C2 => 
                           n159, ZN => intadd_1_B_12_port);
   U305 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_17, B1 => 
                           OP_A_12_port, B2 => n160, C1 => OP_A_13_port, C2 => 
                           n159, ZN => intadd_1_B_11_port);
   U306 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_16, B1 => 
                           OP_A_12_port, B2 => n159, C1 => OP_A_11_port, C2 => 
                           n160, ZN => intadd_1_B_10_port);
   U307 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_14, B1 => n159, B2 
                           => OP_A_10_port, C1 => n160, C2 => OP_A_9_port, ZN 
                           => intadd_1_B_8_port);
   U308 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_13, B1 => n159, B2 
                           => OP_A_9_port, C1 => n160, C2 => OP_A_8_port, ZN =>
                           intadd_1_B_7_port);
   U309 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_12, B1 => n159, B2 
                           => OP_A_8_port, C1 => n160, C2 => OP_A_7_port, ZN =>
                           intadd_1_B_6_port);
   U310 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_11, B1 => n159, B2 
                           => OP_A_7_port, C1 => n160, C2 => OP_A_6_port, ZN =>
                           intadd_1_B_5_port);
   U311 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_10, B1 => n159, B2 
                           => OP_A_6_port, C1 => n160, C2 => OP_A_5_port, ZN =>
                           intadd_1_B_4_port);
   U312 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_9, B1 => n159, B2 
                           => OP_A_5_port, C1 => n160, C2 => OP_A_4_port, ZN =>
                           intadd_1_B_3_port);
   U313 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_8, B1 => n159, B2 
                           => OP_A_4_port, C1 => n160, C2 => OP_A_3_port, ZN =>
                           intadd_1_B_2_port);
   U314 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_7, B1 => n159, B2 
                           => OP_A_3_port, C1 => n160, C2 => OP_A_2_port, ZN =>
                           intadd_1_B_1_port);
   U315 : AOI222_X1 port map( A1 => n1413, A2 => C430_DATA4_6, B1 => 
                           OP_A_1_port, B2 => n160, C1 => n159, C2 => 
                           OP_A_2_port, ZN => intadd_1_B_0_port);
   U316 : INV_X1 port map( A => n161, ZN => n162);
   U317 : AOI222_X1 port map( A1 => n1083, A2 => C429_DATA4_17, B1 => n60, B2 
                           => OP_A_11_port, C1 => n1027, C2 => OP_A_10_port, ZN
                           => intadd_2_A_9_port);
   U318 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_16, B1 => n60, B2 
                           => OP_A_10_port, C1 => n1027, C2 => OP_A_9_port, ZN 
                           => intadd_2_A_8_port);
   U319 : AOI222_X1 port map( A1 => n1083, A2 => C429_DATA4_15, B1 => n60, B2 
                           => OP_A_9_port, C1 => n1027, C2 => OP_A_8_port, ZN 
                           => intadd_2_A_7_port);
   U320 : AOI222_X1 port map( A1 => n1083, A2 => C429_DATA4_14, B1 => n60, B2 
                           => OP_A_8_port, C1 => n1027, C2 => OP_A_7_port, ZN 
                           => intadd_2_A_6_port);
   U321 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_13, B1 => n60, B2 
                           => OP_A_7_port, C1 => n1027, C2 => OP_A_6_port, ZN 
                           => intadd_2_A_5_port);
   U322 : AOI222_X1 port map( A1 => n1083, A2 => C429_DATA4_12, B1 => n60, B2 
                           => OP_A_6_port, C1 => n1027, C2 => OP_A_5_port, ZN 
                           => intadd_2_A_4_port);
   U323 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_11, B1 => n60, B2 
                           => OP_A_5_port, C1 => n1027, C2 => OP_A_4_port, ZN 
                           => intadd_2_A_3_port);
   U324 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_10, B1 => n60, B2 
                           => OP_A_4_port, C1 => n1027, C2 => OP_A_3_port, ZN 
                           => intadd_2_A_2_port);
   U325 : AOI222_X1 port map( A1 => n1083, A2 => C429_DATA4_9, B1 => n60, B2 =>
                           OP_A_3_port, C1 => n1027, C2 => OP_A_2_port, ZN => 
                           intadd_2_A_1_port);
   U326 : AND2_X1 port map( A1 => C2_DATA1_6, A2 => n163, ZN => n164);
   U327 : AOI21_X1 port map( B1 => OP_A_0_port, B2 => n60, A => n164, ZN => 
                           n620);
   U328 : NOR2_X1 port map( A1 => intadd_1_SUM_0_port, A2 => n620, ZN => n619);
   U329 : INV_X1 port map( A => intadd_1_SUM_1_port, ZN => n166);
   U330 : INV_X1 port map( A => n619, ZN => n641);
   U331 : AOI222_X1 port map( A1 => n1083, A2 => C429_DATA4_7, B1 => n60, B2 =>
                           OP_A_1_port, C1 => n1027, C2 => OP_A_0_port, ZN => 
                           n642);
   U332 : OAI21_X1 port map( B1 => intadd_1_SUM_1_port, B2 => n641, A => n642, 
                           ZN => n165);
   U333 : OAI21_X1 port map( B1 => n619, B2 => n166, A => n165, ZN => 
                           intadd_2_A_0_port);
   U334 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_8, B1 => n60, B2 =>
                           OP_A_2_port, C1 => n1027, C2 => OP_A_1_port, ZN => 
                           intadd_2_B_0_port);
   U335 : AOI21_X1 port map( B1 => n168, B2 => n170, A => n167, ZN => n169);
   U336 : OAI21_X1 port map( B1 => n173, B2 => n170, A => n169, ZN => N287);
   U337 : AOI21_X1 port map( B1 => n171, B2 => n1409, A => n178, ZN => n172);
   U338 : INV_X1 port map( A => n172, ZN => n174);
   U339 : OAI211_X1 port map( C1 => n175, C2 => n1408, A => n174, B => n173, ZN
                           => N288);
   U340 : INV_X1 port map( A => n176, ZN => n177);
   U341 : OAI21_X1 port map( B1 => n178, B2 => n1406, A => n177, ZN => N289);
   U342 : INV_X1 port map( A => OP2(0), ZN => n217);
   U343 : AOI22_X1 port map( A1 => OP2(0), A2 => n193, B1 => n195, B2 => n217, 
                           ZN => N247);
   U344 : INV_X1 port map( A => OP2(1), ZN => n483);
   U345 : AOI22_X1 port map( A1 => OP2(1), A2 => n193, B1 => n195, B2 => n483, 
                           ZN => N248);
   U346 : INV_X1 port map( A => OP2(2), ZN => n179);
   U347 : AOI22_X1 port map( A1 => OP2(2), A2 => n193, B1 => n195, B2 => n179, 
                           ZN => N249);
   U348 : INV_X1 port map( A => OP2(3), ZN => n180);
   U349 : AOI22_X1 port map( A1 => OP2(3), A2 => n193, B1 => n195, B2 => n180, 
                           ZN => N250);
   U350 : INV_X1 port map( A => OP2(4), ZN => n181);
   U351 : AOI22_X1 port map( A1 => OP2(4), A2 => n193, B1 => n195, B2 => n181, 
                           ZN => N251);
   U352 : INV_X1 port map( A => OP2(5), ZN => n612);
   U353 : AOI22_X1 port map( A1 => OP2(5), A2 => n193, B1 => n195, B2 => n612, 
                           ZN => N252);
   U354 : INV_X1 port map( A => OP2(6), ZN => n182);
   U355 : AOI22_X1 port map( A1 => OP2(6), A2 => n193, B1 => n195, B2 => n182, 
                           ZN => N253);
   U356 : INV_X1 port map( A => OP2(7), ZN => n664);
   U357 : AOI22_X1 port map( A1 => OP2(7), A2 => n204, B1 => n195, B2 => n664, 
                           ZN => N254);
   U358 : INV_X1 port map( A => OP2(8), ZN => n183);
   U359 : AOI22_X1 port map( A1 => OP2(8), A2 => n204, B1 => n195, B2 => n183, 
                           ZN => N255);
   U360 : INV_X1 port map( A => OP2(9), ZN => n691);
   U361 : AOI22_X1 port map( A1 => OP2(9), A2 => n204, B1 => n195, B2 => n691, 
                           ZN => N256);
   U362 : INV_X1 port map( A => OP2(10), ZN => n184);
   U363 : AOI22_X1 port map( A1 => OP2(10), A2 => n204, B1 => n195, B2 => n184,
                           ZN => N257);
   U364 : INV_X1 port map( A => OP2(11), ZN => n185);
   U365 : AOI22_X1 port map( A1 => OP2(11), A2 => n204, B1 => n195, B2 => n185,
                           ZN => N258);
   U366 : INV_X1 port map( A => OP2(12), ZN => n776);
   U367 : AOI22_X1 port map( A1 => OP2(12), A2 => n204, B1 => n195, B2 => n776,
                           ZN => N259);
   U368 : INV_X1 port map( A => OP2(13), ZN => n800);
   U369 : AOI22_X1 port map( A1 => OP2(13), A2 => n204, B1 => n195, B2 => n800,
                           ZN => N260);
   U370 : INV_X1 port map( A => OP2(14), ZN => n186);
   U371 : AOI22_X1 port map( A1 => OP2(14), A2 => n204, B1 => n195, B2 => n186,
                           ZN => N261);
   U372 : INV_X1 port map( A => OP2(15), ZN => n859);
   U373 : AOI22_X1 port map( A1 => OP2(15), A2 => n204, B1 => n195, B2 => n859,
                           ZN => N262);
   U374 : INV_X1 port map( A => OP2(16), ZN => n187);
   U375 : AOI22_X1 port map( A1 => OP2(16), A2 => n204, B1 => n195, B2 => n187,
                           ZN => N263);
   U376 : INV_X1 port map( A => OP2(17), ZN => n188);
   U377 : AOI22_X1 port map( A1 => OP2(17), A2 => n193, B1 => n195, B2 => n188,
                           ZN => N264);
   U378 : INV_X1 port map( A => OP2(18), ZN => n189);
   U379 : AOI22_X1 port map( A1 => OP2(18), A2 => n193, B1 => n195, B2 => n189,
                           ZN => N265);
   U380 : INV_X1 port map( A => OP2(19), ZN => n190);
   U381 : AOI22_X1 port map( A1 => OP2(19), A2 => n193, B1 => n195, B2 => n190,
                           ZN => N266);
   U382 : INV_X1 port map( A => OP2(20), ZN => n191);
   U383 : AOI22_X1 port map( A1 => OP2(20), A2 => n193, B1 => n195, B2 => n191,
                           ZN => N267);
   U384 : INV_X1 port map( A => OP2(21), ZN => n192);
   U385 : AOI22_X1 port map( A1 => OP2(21), A2 => n193, B1 => n195, B2 => n192,
                           ZN => N268);
   U386 : INV_X1 port map( A => OP2(22), ZN => n194);
   U387 : AOI22_X1 port map( A1 => OP2(22), A2 => n204, B1 => n195, B2 => n194,
                           ZN => N269);
   U388 : INV_X1 port map( A => OP2(23), ZN => n196);
   U389 : AOI22_X1 port map( A1 => OP2(23), A2 => n204, B1 => n195, B2 => n196,
                           ZN => N270);
   U390 : INV_X1 port map( A => OP2(24), ZN => n1138);
   U391 : AOI22_X1 port map( A1 => OP2(24), A2 => n204, B1 => n195, B2 => n1138
                           , ZN => N271);
   U392 : INV_X1 port map( A => OP2(25), ZN => n197);
   U393 : AOI22_X1 port map( A1 => OP2(25), A2 => n204, B1 => n195, B2 => n197,
                           ZN => N272);
   U394 : INV_X1 port map( A => OP2(26), ZN => n198);
   U395 : AOI22_X1 port map( A1 => OP2(26), A2 => n204, B1 => n195, B2 => n198,
                           ZN => N273);
   U396 : INV_X1 port map( A => OP2(27), ZN => n199);
   U397 : AOI22_X1 port map( A1 => OP2(27), A2 => n204, B1 => n195, B2 => n199,
                           ZN => N274);
   U398 : INV_X1 port map( A => OP2(28), ZN => n200);
   U399 : AOI22_X1 port map( A1 => OP2(28), A2 => n204, B1 => n195, B2 => n200,
                           ZN => N275);
   U400 : INV_X1 port map( A => OP2(29), ZN => n201);
   U401 : AOI22_X1 port map( A1 => OP2(29), A2 => n204, B1 => n195, B2 => n201,
                           ZN => N276);
   U402 : INV_X1 port map( A => OP2(30), ZN => n202);
   U403 : AOI22_X1 port map( A1 => OP2(30), A2 => n204, B1 => n195, B2 => n202,
                           ZN => N277);
   U404 : INV_X1 port map( A => OP2(31), ZN => n203);
   U405 : AOI22_X1 port map( A1 => OP2(31), A2 => n204, B1 => n195, B2 => n203,
                           ZN => N278);
   U406 : INV_X1 port map( A => N284, ZN => n1159);
   U407 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => n55, ZN => n1204);
   U408 : NAND2_X1 port map( A1 => n542, A2 => OP_A_21_port, ZN => n1058);
   U409 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => n603, ZN => n1133);
   U410 : OR2_X1 port map( A1 => OP_B_1_port, A2 => OP_B_0_port, ZN => n607);
   U411 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => n56, ZN => n1002);
   U412 : AND4_X1 port map( A1 => n1204, A2 => n1058, A3 => n1133, A4 => n1002,
                           ZN => n784);
   U413 : NAND2_X1 port map( A1 => n491, A2 => OP_A_25_port, ZN => n1205);
   U414 : NAND2_X1 port map( A1 => OP_A_27_port, A2 => n55, ZN => n1318);
   U415 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => n56, ZN => n1130);
   U416 : CLKBUF_X1 port map( A => n603, Z => n553);
   U417 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => n553, ZN => n1272);
   U418 : NAND4_X1 port map( A1 => n1205, A2 => n1318, A3 => n1130, A4 => n1272
                           , ZN => n781);
   U419 : INV_X1 port map( A => n857, ZN => n510);
   U420 : INV_X1 port map( A => OP_A_31_port, ZN => n1370);
   U421 : AOI22_X1 port map( A1 => OP_A_30_port, A2 => n603, B1 => OP_A_28_port
                           , B2 => n56, ZN => n205);
   U422 : NAND2_X1 port map( A1 => n491, A2 => OP_A_29_port, ZN => n1319);
   U423 : OAI211_X1 port map( C1 => n577, C2 => n1370, A => n205, B => n1319, 
                           ZN => n1265);
   U424 : AOI22_X1 port map( A1 => n855, A2 => n781, B1 => n510, B2 => n1265, 
                           ZN => n207);
   U425 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => n55, ZN => n1057);
   U426 : NAND2_X1 port map( A1 => n491, A2 => OP_A_17_port, ZN => n937);
   U427 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => n553, ZN => n1005);
   U428 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n56, ZN => n887);
   U429 : NAND4_X1 port map( A1 => n1057, A2 => n937, A3 => n1005, A4 => n887, 
                           ZN => n777);
   U430 : NAND2_X1 port map( A1 => n894, A2 => n777, ZN => n206);
   U431 : OAI211_X1 port map( C1 => n784, C2 => n742, A => n207, B => n206, ZN 
                           => n898);
   U432 : NAND2_X1 port map( A1 => OP_A_15_port, A2 => n55, ZN => n936);
   U433 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => n56, ZN => n767);
   U434 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => n553, ZN => n889);
   U435 : AND4_X1 port map( A1 => n819, A2 => n936, A3 => n767, A4 => n889, ZN 
                           => n771);
   U436 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n857, ZN => n1352);
   U437 : INV_X1 port map( A => n1352, ZN => n891);
   U438 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => n55, ZN => n817);
   U439 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => n553, ZN => n768);
   U440 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => n56, ZN => n672);
   U441 : AND4_X1 port map( A1 => n817, A2 => n726, A3 => n768, A4 => n672, ZN 
                           => n681);
   U442 : INV_X1 port map( A => n855, ZN => n741);
   U443 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n741, ZN => n1350);
   U444 : INV_X1 port map( A => n1350, ZN => n566);
   U445 : OAI22_X1 port map( A1 => n771, A2 => n891, B1 => n681, B2 => n566, ZN
                           => n213);
   U446 : NAND2_X1 port map( A1 => OP_A_3_port, A2 => n55, ZN => n626);
   U447 : NAND2_X1 port map( A1 => n491, A2 => OP_A_1_port, ZN => n507);
   U448 : NAND2_X1 port map( A1 => OP_A_0_port, A2 => n56, ZN => n895);
   U449 : NAND2_X1 port map( A1 => OP_A_2_port, A2 => n553, ZN => n208);
   U450 : AND4_X1 port map( A1 => n626, A2 => n507, A3 => n895, A4 => n208, ZN 
                           => n211);
   U451 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n765, ZN => n1360);
   U452 : INV_X1 port map( A => n1360, ZN => n1261);
   U453 : NAND2_X1 port map( A1 => OP_A_7_port, A2 => n55, ZN => n725);
   U454 : NAND2_X1 port map( A1 => OP_A_4_port, A2 => n56, ZN => n209);
   U455 : NAND2_X1 port map( A1 => OP_A_6_port, A2 => n553, ZN => n674);
   U456 : NAND4_X1 port map( A1 => n725, A2 => n628, A3 => n209, A4 => n674, ZN
                           => n582);
   U457 : INV_X1 port map( A => n582, ZN => n210);
   U458 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n742, ZN => n1358);
   U459 : INV_X1 port map( A => n1358, ZN => n899);
   U460 : OAI22_X1 port map( A1 => n211, A2 => n1261, B1 => n210, B2 => n899, 
                           ZN => n212);
   U461 : AOI211_X1 port map( C1 => OP_B_4_port, C2 => n898, A => n213, B => 
                           n212, ZN => n481);
   U462 : NOR2_X1 port map( A1 => n215, A2 => n214, ZN => n1347);
   U463 : CLKBUF_X1 port map( A => n1347, Z => n1330);
   U464 : NAND2_X1 port map( A1 => OP_B_0_port, A2 => OP_A_0_port, ZN => n292);
   U465 : OR2_X1 port map( A1 => n216, A2 => n1411, ZN => n1139);
   U466 : OAI22_X1 port map( A1 => n1396, A2 => n292, B1 => n1139, B2 => n217, 
                           ZN => n220);
   U467 : NOR2_X1 port map( A1 => n218, A2 => OP_LOGIC_0_port, ZN => n474);
   U468 : INV_X1 port map( A => OP_LOGIC_1_port, ZN => n221);
   U469 : AND2_X1 port map( A1 => n474, A2 => n221, ZN => n1245);
   U470 : INV_X1 port map( A => n1228, ZN => n1061);
   U471 : OAI22_X1 port map( A1 => n292, A2 => n1369, B1 => n895, B2 => n1061, 
                           ZN => n219);
   U472 : AOI211_X1 port map( C1 => n1330, C2 => OP1(0), A => n220, B => n219, 
                           ZN => n480);
   U473 : NAND3_X1 port map( A1 => N281, A2 => n221, A3 => OP_LOGIC_0_port, ZN 
                           => n1368);
   U474 : INV_X1 port map( A => OP_A_0_port, ZN => n549);
   U475 : NAND2_X1 port map( A1 => n222, A2 => n549, ZN => n487);
   U476 : NOR2_X1 port map( A1 => OP_B_3_port, A2 => n550, ZN => n364);
   U477 : INV_X1 port map( A => n364, ZN => n315);
   U478 : INV_X1 port map( A => OP_A_5_port, ZN => n606);
   U479 : NAND2_X1 port map( A1 => n606, A2 => OP_B_5_port, ZN => n368);
   U480 : OAI21_X1 port map( B1 => n1363, B2 => OP_A_4_port, A => n368, ZN => 
                           n319);
   U481 : INV_X1 port map( A => OP_A_1_port, ZN => n578);
   U482 : OAI21_X1 port map( B1 => n223, B2 => OP_A_1_port, A => OP_A_0_port, 
                           ZN => n314);
   U483 : OAI211_X1 port map( C1 => n578, C2 => n55, A => n607, B => n314, ZN 
                           => n365);
   U484 : NOR2_X1 port map( A1 => OP_A_3_port, A2 => n1160, ZN => n301);
   U485 : AOI21_X1 port map( B1 => n576, B2 => OP_B_2_port, A => n301, ZN => 
                           n363);
   U486 : INV_X1 port map( A => n301, ZN => n316);
   U487 : NOR2_X1 port map( A1 => n576, A2 => OP_B_2_port, ZN => n224);
   U488 : AOI22_X1 port map( A1 => n365, A2 => n363, B1 => n316, B2 => n224, ZN
                           => n226);
   U489 : INV_X1 port map( A => OP_A_4_port, ZN => n367);
   U490 : NOR2_X1 port map( A1 => n367, A2 => OP_B_4_port, ZN => n225);
   U491 : NOR2_X1 port map( A1 => n606, A2 => OP_B_5_port, ZN => n370);
   U492 : AOI21_X1 port map( B1 => n368, B2 => n225, A => n370, ZN => n318);
   U493 : OAI221_X1 port map( B1 => n315, B2 => n319, C1 => n226, C2 => n319, A
                           => n318, ZN => n232);
   U494 : NAND2_X1 port map( A1 => n377, A2 => OP_A_6_port, ZN => n227);
   U495 : NOR2_X1 port map( A1 => n294, A2 => OP_A_7_port, ZN => n378);
   U496 : NAND2_X1 port map( A1 => n294, A2 => OP_A_7_port, ZN => n379);
   U497 : OAI21_X1 port map( B1 => n227, B2 => n378, A => n379, ZN => n321);
   U498 : INV_X1 port map( A => OP_A_6_port, ZN => n371);
   U499 : AOI21_X1 port map( B1 => n371, B2 => OP_B_6_port, A => n378, ZN => 
                           n323);
   U500 : INV_X1 port map( A => OP_A_12_port, ZN => n233);
   U501 : NAND2_X1 port map( A1 => n233, A2 => OP_B_12_port, ZN => n332);
   U502 : INV_X1 port map( A => OP_A_13_port, ZN => n234);
   U503 : INV_X1 port map( A => OP_B_14_port, ZN => n228);
   U504 : NAND2_X1 port map( A1 => n1080, A2 => OP_B_15_port, ZN => n348);
   U505 : OAI21_X1 port map( B1 => n228, B2 => OP_A_14_port, A => n348, ZN => 
                           n229);
   U506 : AOI21_X1 port map( B1 => n234, B2 => OP_B_13_port, A => n229, ZN => 
                           n240);
   U507 : AND2_X1 port map( A1 => n332, A2 => n240, ZN => n230);
   U508 : INV_X1 port map( A => OP_A_10_port, ZN => n335);
   U509 : INV_X1 port map( A => OP_A_11_port, ZN => n235);
   U510 : NAND2_X1 port map( A1 => n235, A2 => OP_B_11_port, ZN => n342);
   U511 : INV_X1 port map( A => n342, ZN => n239);
   U512 : AOI21_X1 port map( B1 => OP_B_10_port, B2 => n335, A => n239, ZN => 
                           n237);
   U513 : INV_X1 port map( A => OP_A_9_port, ZN => n302);
   U514 : INV_X1 port map( A => OP_A_8_port, ZN => n236);
   U515 : AOI22_X1 port map( A1 => OP_B_9_port, A2 => n302, B1 => OP_B_8_port, 
                           B2 => n236, ZN => n338);
   U516 : NAND3_X1 port map( A1 => n230, A2 => n237, A3 => n338, ZN => n325);
   U517 : INV_X1 port map( A => n325, ZN => n231);
   U518 : OAI221_X1 port map( B1 => n232, B2 => n321, C1 => n323, C2 => n321, A
                           => n231, ZN => n248_port);
   U519 : INV_X1 port map( A => OP_A_14_port, ZN => n331);
   U520 : NOR2_X1 port map( A1 => n331, A2 => OP_B_14_port, ZN => n345);
   U521 : OAI22_X1 port map( A1 => OP_B_13_port, A2 => n234, B1 => OP_B_12_port
                           , B2 => n233, ZN => n334);
   U522 : OR2_X1 port map( A1 => n335, A2 => OP_B_10_port, ZN => n336);
   U523 : NOR2_X1 port map( A1 => n235, A2 => OP_B_11_port, ZN => n344);
   U524 : INV_X1 port map( A => n344, ZN => n337);
   U525 : INV_X1 port map( A => OP_B_9_port, ZN => n339);
   U526 : OAI22_X1 port map( A1 => OP_B_8_port, A2 => n236, B1 => OP_B_9_port, 
                           B2 => n302, ZN => n356);
   U527 : OAI211_X1 port map( C1 => OP_A_9_port, C2 => n339, A => n237, B => 
                           n356, ZN => n238);
   U528 : OAI211_X1 port map( C1 => n239, C2 => n336, A => n337, B => n238, ZN 
                           => n241);
   U529 : OAI221_X1 port map( B1 => n334, B2 => n332, C1 => n334, C2 => n241, A
                           => n240, ZN => n242);
   U530 : INV_X1 port map( A => n242, ZN => n243);
   U531 : NOR2_X1 port map( A1 => n1080, A2 => OP_B_15_port, ZN => n351);
   U532 : AOI211_X1 port map( C1 => n348, C2 => n345, A => n243, B => n351, ZN 
                           => n326);
   U533 : INV_X1 port map( A => OP_B_17_port, ZN => n255_port);
   U534 : NOR2_X1 port map( A1 => OP_A_17_port, A2 => n255_port, ZN => n393);
   U535 : INV_X1 port map( A => OP_B_16_port, ZN => n256_port);
   U536 : NOR2_X1 port map( A1 => OP_A_16_port, A2 => n256_port, ZN => n394);
   U537 : INV_X1 port map( A => OP_B_18_port, ZN => n357);
   U538 : INV_X1 port map( A => OP_A_19_port, ZN => n254_port);
   U539 : NAND2_X1 port map( A1 => OP_B_19_port, A2 => n254_port, ZN => n396);
   U540 : OAI21_X1 port map( B1 => OP_A_18_port, B2 => n357, A => n396, ZN => 
                           n257_port);
   U541 : INV_X1 port map( A => OP_A_21_port, ZN => n245);
   U542 : INV_X1 port map( A => OP_B_22_port, ZN => n389);
   U543 : INV_X1 port map( A => OP_A_23_port, ZN => n252_port);
   U544 : NAND2_X1 port map( A1 => OP_B_23_port, A2 => n252_port, ZN => n407);
   U545 : OAI21_X1 port map( B1 => OP_A_22_port, B2 => n389, A => n407, ZN => 
                           n244);
   U546 : AOI21_X1 port map( B1 => OP_B_21_port, B2 => n245, A => n244, ZN => 
                           n246_port);
   U547 : INV_X1 port map( A => n246_port, ZN => n260_port);
   U548 : INV_X1 port map( A => OP_B_20_port, ZN => n253_port);
   U549 : NOR2_X1 port map( A1 => n253_port, A2 => OP_A_20_port, ZN => n399);
   U550 : OR2_X1 port map( A1 => n260_port, A2 => n399, ZN => n247_port);
   U551 : OR4_X1 port map( A1 => n393, A2 => n394, A3 => n257_port, A4 => 
                           n247_port, ZN => n324);
   U552 : AOI21_X1 port map( B1 => n248_port, B2 => n326, A => n324, ZN => 
                           n249_port);
   U553 : INV_X1 port map( A => n249_port, ZN => n284_port);
   U554 : INV_X1 port map( A => OP_B_24_port, ZN => n416);
   U555 : INV_X1 port map( A => OP_A_25_port, ZN => n265_port);
   U556 : NAND2_X1 port map( A1 => n265_port, A2 => OP_B_25_port, ZN => n417);
   U557 : INV_X1 port map( A => OP_A_26_port, ZN => n422);
   U558 : INV_X1 port map( A => OP_A_27_port, ZN => n1248);
   U559 : NAND2_X1 port map( A1 => OP_B_27_port, A2 => n1248, ZN => n424);
   U560 : INV_X1 port map( A => n424, ZN => n270_port);
   U561 : AOI21_X1 port map( B1 => n422, B2 => OP_B_26_port, A => n270_port, ZN
                           => n266_port);
   U562 : OAI211_X1 port map( C1 => n416, C2 => OP_A_24_port, A => n417, B => 
                           n266_port, ZN => n276_port);
   U563 : INV_X1 port map( A => OP_B_28_port, ZN => n274_port);
   U564 : INV_X1 port map( A => OP_A_29_port, ZN => n1297);
   U565 : NAND2_X1 port map( A1 => n1297, A2 => OP_B_29_port, ZN => n412);
   U566 : NOR2_X1 port map( A1 => OP_B_31_port, A2 => n1370, ZN => n427);
   U567 : INV_X1 port map( A => OP_A_30_port, ZN => n251_port);
   U568 : NAND2_X1 port map( A1 => OP_B_30_port, A2 => n251_port, ZN => n451);
   U569 : INV_X1 port map( A => n451, ZN => n410);
   U570 : NOR2_X1 port map( A1 => n427, A2 => n410, ZN => n271_port);
   U571 : OAI211_X1 port map( C1 => n274_port, C2 => OP_A_28_port, A => n412, B
                           => n271_port, ZN => n250_port);
   U572 : OR2_X1 port map( A1 => n276_port, A2 => n250_port, ZN => n462);
   U573 : NOR2_X1 port map( A1 => OP_B_30_port, A2 => n251_port, ZN => n439);
   U574 : INV_X1 port map( A => n427, ZN => n449);
   U575 : NAND2_X1 port map( A1 => n1370, A2 => OP_B_31_port, ZN => n305);
   U576 : INV_X1 port map( A => n305, ZN => n452);
   U577 : AND2_X1 port map( A1 => n389, A2 => OP_A_22_port, ZN => n263_port);
   U578 : NOR2_X1 port map( A1 => OP_B_23_port, A2 => n252_port, ZN => n408);
   U579 : INV_X1 port map( A => OP_B_21_port, ZN => n401);
   U580 : AOI22_X1 port map( A1 => OP_A_21_port, A2 => n401, B1 => OP_A_20_port
                           , B2 => n253_port, ZN => n403);
   U581 : INV_X1 port map( A => OP_A_18_port, ZN => n390);
   U582 : NOR2_X1 port map( A1 => OP_B_18_port, A2 => n390, ZN => n259_port);
   U583 : NOR2_X1 port map( A1 => OP_B_19_port, A2 => n254_port, ZN => n397);
   U584 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n255_port, ZN => n392);
   U585 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n256_port, ZN => n359);
   U586 : AOI211_X1 port map( C1 => n392, C2 => n359, A => n393, B => n257_port
                           , ZN => n258_port);
   U587 : AOI211_X1 port map( C1 => n259_port, C2 => n396, A => n397, B => 
                           n258_port, ZN => n261_port);
   U588 : AOI221_X1 port map( B1 => n399, B2 => n403, C1 => n261_port, C2 => 
                           n403, A => n260_port, ZN => n262_port);
   U589 : AOI211_X1 port map( C1 => n263_port, C2 => n407, A => n408, B => 
                           n262_port, ZN => n282_port);
   U590 : INV_X1 port map( A => n412, ZN => n288_port);
   U591 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n274_port, ZN => 
                           n264_port);
   U592 : NOR2_X1 port map( A1 => OP_B_29_port, A2 => n1297, ZN => n414);
   U593 : INV_X1 port map( A => n414, ZN => n361);
   U594 : OAI21_X1 port map( B1 => n288_port, B2 => n264_port, A => n361, ZN =>
                           n280_port);
   U595 : INV_X1 port map( A => OP_A_28_port, ZN => n411);
   U596 : AOI21_X1 port map( B1 => OP_B_28_port, B2 => n411, A => n288_port, ZN
                           => n279_port);
   U597 : OR2_X1 port map( A1 => n422, A2 => OP_B_26_port, ZN => n269_port);
   U598 : NOR2_X1 port map( A1 => OP_B_25_port, A2 => n265_port, ZN => n418);
   U599 : AND2_X1 port map( A1 => n416, A2 => OP_A_24_port, ZN => n267_port);
   U600 : OAI211_X1 port map( C1 => n418, C2 => n267_port, A => n417, B => 
                           n266_port, ZN => n268_port);
   U601 : OR2_X1 port map( A1 => n1248, A2 => OP_B_27_port, ZN => n421);
   U602 : OAI211_X1 port map( C1 => n270_port, C2 => n269_port, A => n268_port,
                           B => n421, ZN => n278_port);
   U603 : OAI221_X1 port map( B1 => n280_port, B2 => n279_port, C1 => n280_port
                           , C2 => n278_port, A => n271_port, ZN => n272_port);
   U604 : OAI21_X1 port map( B1 => n282_port, B2 => n462, A => n272_port, ZN =>
                           n273_port);
   U605 : AOI211_X1 port map( C1 => n439, C2 => n449, A => n452, B => n273_port
                           , ZN => n460);
   U606 : OAI21_X1 port map( B1 => n284_port, B2 => n462, A => n460, ZN => 
                           n286_port);
   U607 : NOR2_X1 port map( A1 => OP_COMPARE_1_port, A2 => OP_COMPARE_2_port, 
                           ZN => n437);
   U608 : NOR2_X1 port map( A1 => n452, A2 => n410, ZN => n277_port);
   U609 : OAI211_X1 port map( C1 => n274_port, C2 => OP_A_28_port, A => n412, B
                           => n277_port, ZN => n275_port);
   U610 : OR2_X1 port map( A1 => n276_port, A2 => n275_port, ZN => n329);
   U611 : OAI221_X1 port map( B1 => n280_port, B2 => n279_port, C1 => n280_port
                           , C2 => n278_port, A => n277_port, ZN => n281_port);
   U612 : OAI21_X1 port map( B1 => n282_port, B2 => n329, A => n281_port, ZN =>
                           n283_port);
   U613 : AOI211_X1 port map( C1 => n439, C2 => n305, A => n427, B => n283_port
                           , ZN => n328);
   U614 : OAI211_X1 port map( C1 => n329, C2 => n284_port, A => 
                           OP_COMPARE_0_port, B => n328, ZN => n285_port);
   U615 : OAI211_X1 port map( C1 => OP_COMPARE_0_port, C2 => n286_port, A => 
                           n437, B => n285_port, ZN => n473);
   U616 : INV_X1 port map( A => OP_COMPARE_3_port, ZN => n472);
   U617 : NAND2_X1 port map( A1 => n424, A2 => n421, ZN => n1241);
   U618 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => OP_B_19_port, ZN => n975
                           );
   U619 : OR2_X1 port map( A1 => OP_A_19_port, A2 => OP_B_19_port, ZN => n991);
   U620 : NAND2_X1 port map( A1 => n975, A2 => n991, ZN => n974);
   U621 : INV_X1 port map( A => n974, ZN => n983);
   U622 : NOR2_X1 port map( A1 => OP_A_23_port, A2 => OP_B_23_port, ZN => n1108
                           );
   U623 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => OP_B_23_port, ZN => 
                           n1123);
   U624 : INV_X1 port map( A => n1123, ZN => n287_port);
   U625 : NOR2_X1 port map( A1 => n1108, A2 => n287_port, ZN => n1106);
   U626 : AND2_X1 port map( A1 => OP_A_15_port, A2 => OP_B_15_port, ZN => n877)
                           ;
   U627 : NOR2_X1 port map( A1 => OP_A_15_port, A2 => OP_B_15_port, ZN => n862)
                           ;
   U628 : NOR2_X1 port map( A1 => n877, A2 => n862, ZN => n873);
   U629 : OR4_X1 port map( A1 => n1241, A2 => n983, A3 => n1106, A4 => n873, ZN
                           => n300);
   U630 : NOR2_X1 port map( A1 => n288_port, A2 => n414, ZN => n1302);
   U631 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => OP_B_26_port, ZN => 
                           n1237);
   U632 : OAI21_X1 port map( B1 => OP_A_26_port, B2 => OP_B_26_port, A => n1237
                           , ZN => n1200);
   U633 : NOR2_X1 port map( A1 => OP_A_30_port, A2 => OP_B_30_port, ZN => n1375
                           );
   U634 : NAND2_X1 port map( A1 => OP_A_30_port, A2 => OP_B_30_port, ZN => 
                           n1377);
   U635 : INV_X1 port map( A => n1377, ZN => n289_port);
   U636 : NOR2_X1 port map( A1 => n1375, A2 => n289_port, ZN => n1343);
   U637 : INV_X1 port map( A => n1343, ZN => n1333);
   U638 : NOR2_X1 port map( A1 => OP_A_28_port, A2 => OP_B_28_port, ZN => n1299
                           );
   U639 : INV_X1 port map( A => n1299, ZN => n290);
   U640 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => OP_B_28_port, ZN => 
                           n1301);
   U641 : NAND2_X1 port map( A1 => n290, A2 => n1301, ZN => n1267);
   U642 : NAND4_X1 port map( A1 => n1302, A2 => n1200, A3 => n1333, A4 => n1267
                           , ZN => n299);
   U643 : NAND2_X1 port map( A1 => n1363, A2 => n367, ZN => n597);
   U644 : NAND2_X1 port map( A1 => OP_B_4_port, A2 => OP_A_4_port, ZN => n570);
   U645 : NAND2_X1 port map( A1 => n597, A2 => n570, ZN => n573);
   U646 : NAND2_X1 port map( A1 => n581, A2 => n576, ZN => n546);
   U647 : NOR2_X1 port map( A1 => n581, A2 => n576, ZN => n506);
   U648 : INV_X1 port map( A => n506, ZN => n291);
   U649 : NAND2_X1 port map( A1 => n546, A2 => n291, ZN => n523);
   U650 : NOR2_X1 port map( A1 => OP_B_1_port, A2 => OP_A_1_port, ZN => n520);
   U651 : INV_X1 port map( A => n520, ZN => n502);
   U652 : NAND2_X1 port map( A1 => OP_B_1_port, A2 => OP_A_1_port, ZN => n519);
   U653 : NAND2_X1 port map( A1 => n502, A2 => n519, ZN => n505);
   U654 : NAND2_X1 port map( A1 => n292, A2 => n487, ZN => n475);
   U655 : NAND4_X1 port map( A1 => n573, A2 => n523, A3 => n505, A4 => n475, ZN
                           => n298);
   U656 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => OP_B_11_port, ZN => n749
                           );
   U657 : OR2_X1 port map( A1 => OP_A_11_port, A2 => OP_B_11_port, ZN => n773);
   U658 : NAND2_X1 port map( A1 => n749, A2 => n773, ZN => n754);
   U659 : NAND2_X1 port map( A1 => OP_B_7_port, A2 => OP_A_7_port, ZN => n645);
   U660 : INV_X1 port map( A => OP_A_7_port, ZN => n293);
   U661 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => n678);
   U662 : NAND2_X1 port map( A1 => n645, A2 => n678, ZN => n653);
   U663 : NAND2_X1 port map( A1 => OP_B_6_port, A2 => OP_A_6_port, ZN => n649);
   U664 : NOR2_X1 port map( A1 => OP_B_6_port, A2 => OP_A_6_port, ZN => n651);
   U665 : INV_X1 port map( A => n651, ZN => n295);
   U666 : NAND2_X1 port map( A1 => n649, A2 => n295, ZN => n636);
   U667 : NAND2_X1 port map( A1 => OP_B_5_port, A2 => OP_A_5_port, ZN => n593);
   U668 : NAND2_X1 port map( A1 => n296, A2 => n606, ZN => n632);
   U669 : NAND2_X1 port map( A1 => n593, A2 => n632, ZN => n600);
   U670 : NAND4_X1 port map( A1 => n754, A2 => n653, A3 => n636, A4 => n600, ZN
                           => n297);
   U671 : NOR4_X1 port map( A1 => n300, A2 => n299, A3 => n298, A4 => n297, ZN 
                           => n313);
   U672 : NOR2_X1 port map( A1 => n364, A2 => n301, ZN => n557);
   U673 : NOR2_X1 port map( A1 => OP_A_13_port, A2 => OP_B_13_port, ZN => n831)
                           ;
   U674 : INV_X1 port map( A => n831, ZN => n793);
   U675 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => OP_B_13_port, ZN => n829
                           );
   U676 : NAND2_X1 port map( A1 => n793, A2 => n829, ZN => n798);
   U677 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => OP_B_8_port, ZN => n711);
   U678 : NOR2_X1 port map( A1 => OP_A_8_port, A2 => OP_B_8_port, ZN => n715);
   U679 : INV_X1 port map( A => n715, ZN => n671);
   U680 : NAND2_X1 port map( A1 => n711, A2 => n671, ZN => n680);
   U681 : NOR2_X1 port map( A1 => OP_A_9_port, A2 => OP_B_9_port, ZN => n714);
   U682 : NOR2_X1 port map( A1 => n302, A2 => n339, ZN => n698);
   U683 : NOR2_X1 port map( A1 => n714, A2 => n698, ZN => n702);
   U684 : INV_X1 port map( A => n702, ZN => n303);
   U685 : NAND4_X1 port map( A1 => n557, A2 => n798, A3 => n680, A4 => n303, ZN
                           => n311);
   U686 : NOR2_X1 port map( A1 => OP_A_21_port, A2 => OP_B_21_port, ZN => n1050
                           );
   U687 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => OP_B_21_port, ZN => 
                           n1048);
   U688 : INV_X1 port map( A => n1048, ZN => n1021);
   U689 : NOR2_X1 port map( A1 => n1050, A2 => n1021, ZN => n1020);
   U690 : NOR2_X1 port map( A1 => OP_A_25_port, A2 => OP_B_25_port, ZN => n1196
                           );
   U691 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => OP_B_25_port, ZN => 
                           n1194);
   U692 : INV_X1 port map( A => n1194, ZN => n304);
   U693 : NOR2_X1 port map( A1 => n1196, A2 => n304, ZN => n1165);
   U694 : NOR2_X1 port map( A1 => OP_A_17_port, A2 => OP_B_17_port, ZN => n953)
                           ;
   U695 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => OP_B_17_port, ZN => n951
                           );
   U696 : INV_X1 port map( A => n951, ZN => n928);
   U697 : NOR2_X1 port map( A1 => n953, A2 => n928, ZN => n918);
   U698 : NAND2_X1 port map( A1 => n305, A2 => n449, ZN => n1371);
   U699 : OR4_X1 port map( A1 => n1020, A2 => n1165, A3 => n918, A4 => n1371, 
                           ZN => n310);
   U700 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => OP_B_18_port, ZN => n980
                           );
   U701 : INV_X1 port map( A => n980, ZN => n948);
   U702 : NOR2_X1 port map( A1 => OP_A_18_port, A2 => OP_B_18_port, ZN => n982)
                           ;
   U703 : NOR2_X1 port map( A1 => n948, A2 => n982, ZN => n958);
   U704 : INV_X1 port map( A => n958, ZN => n306);
   U705 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => OP_B_20_port, ZN => 
                           n1046);
   U706 : NOR2_X1 port map( A1 => OP_A_20_port, A2 => OP_B_20_port, ZN => n1049
                           );
   U707 : INV_X1 port map( A => n1049, ZN => n1007);
   U708 : NAND2_X1 port map( A1 => n1046, A2 => n1007, ZN => n1018);
   U709 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => OP_B_22_port, ZN => 
                           n1124);
   U710 : OAI21_X1 port map( B1 => OP_A_22_port, B2 => OP_B_22_port, A => n1124
                           , ZN => n1125);
   U711 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => OP_B_24_port, ZN => 
                           n1193);
   U712 : NOR2_X1 port map( A1 => OP_A_24_port, A2 => OP_B_24_port, ZN => n1195
                           );
   U713 : INV_X1 port map( A => n1195, ZN => n1142);
   U714 : NAND2_X1 port map( A1 => n1193, A2 => n1142, ZN => n1129);
   U715 : NAND4_X1 port map( A1 => n306, A2 => n1018, A3 => n1125, A4 => n1129,
                           ZN => n309);
   U716 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => OP_B_10_port, ZN => n755
                           );
   U717 : OAI21_X1 port map( B1 => OP_A_10_port, B2 => OP_B_10_port, A => n755,
                           ZN => n719);
   U718 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => OP_B_12_port, ZN => n827
                           );
   U719 : NOR2_X1 port map( A1 => OP_A_12_port, A2 => OP_B_12_port, ZN => n830)
                           ;
   U720 : INV_X1 port map( A => n830, ZN => n780);
   U721 : NAND2_X1 port map( A1 => n827, A2 => n780, ZN => n779);
   U722 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => OP_B_14_port, ZN => n870
                           );
   U723 : OAI21_X1 port map( B1 => OP_A_14_port, B2 => OP_B_14_port, A => n870,
                           ZN => n835);
   U724 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => OP_B_16_port, ZN => n949
                           );
   U725 : NOR2_X1 port map( A1 => OP_A_16_port, A2 => OP_B_16_port, ZN => n952)
                           ;
   U726 : INV_X1 port map( A => n952, ZN => n307);
   U727 : NAND2_X1 port map( A1 => n949, A2 => n307, ZN => n904);
   U728 : NAND4_X1 port map( A1 => n719, A2 => n779, A3 => n835, A4 => n904, ZN
                           => n308);
   U729 : NOR4_X1 port map( A1 => n311, A2 => n310, A3 => n309, A4 => n308, ZN 
                           => n312);
   U730 : AOI211_X1 port map( C1 => n313, C2 => n312, A => OP_COMPARE_1_port, B
                           => OP_COMPARE_2_port, ZN => n469);
   U731 : OAI22_X1 port map( A1 => OP_B_0_port, A2 => n314, B1 => OP_B_1_port, 
                           B2 => n578, ZN => n317);
   U732 : OAI21_X1 port map( B1 => OP_B_2_port, B2 => n576, A => n315, ZN => 
                           n366);
   U733 : AOI22_X1 port map( A1 => n363, A2 => n317, B1 => n316, B2 => n366, ZN
                           => n320);
   U734 : OAI21_X1 port map( B1 => n320, B2 => n319, A => n318, ZN => n322);
   U735 : AOI21_X1 port map( B1 => n323, B2 => n322, A => n321, ZN => n360);
   U736 : AOI221_X1 port map( B1 => n360, B2 => n326, C1 => n325, C2 => n326, A
                           => n324, ZN => n327);
   U737 : INV_X1 port map( A => n327, ZN => n461);
   U738 : INV_X1 port map( A => OP_COMPARE_1_port, ZN => n459);
   U739 : OAI211_X1 port map( C1 => n329, C2 => n461, A => n459, B => n328, ZN 
                           => n330);
   U740 : INV_X1 port map( A => n330, ZN => n436);
   U741 : NAND2_X1 port map( A1 => OP_B_14_port, A2 => n331, ZN => n350);
   U742 : INV_X1 port map( A => OP_B_13_port, ZN => n333);
   U743 : AOI222_X1 port map( A1 => OP_A_13_port, A2 => n333, B1 => 
                           OP_A_13_port, B2 => n332, C1 => n333, C2 => n332, ZN
                           => n347);
   U744 : INV_X1 port map( A => n334, ZN => n353);
   U745 : NAND2_X1 port map( A1 => OP_B_10_port, A2 => n335, ZN => n343);
   U746 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n354);
   U747 : AOI211_X1 port map( C1 => n339, C2 => OP_A_9_port, A => n354, B => 
                           n338, ZN => n340);
   U748 : INV_X1 port map( A => n340, ZN => n341);
   U749 : OAI211_X1 port map( C1 => n344, C2 => n343, A => n342, B => n341, ZN 
                           => n346);
   U750 : NOR2_X1 port map( A1 => n351, A2 => n345, ZN => n352);
   U751 : OAI221_X1 port map( B1 => n347, B2 => n353, C1 => n347, C2 => n346, A
                           => n352, ZN => n349);
   U752 : OAI211_X1 port map( C1 => n351, C2 => n350, A => n349, B => n348, ZN 
                           => n387);
   U753 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n355);
   U754 : NOR3_X1 port map( A1 => n356, A2 => n355, A3 => n354, ZN => n381);
   U755 : AOI21_X1 port map( B1 => OP_A_22_port, B2 => n389, A => n408, ZN => 
                           n402);
   U756 : AND2_X1 port map( A1 => n403, A2 => n402, ZN => n358);
   U757 : AOI21_X1 port map( B1 => n357, B2 => OP_A_18_port, A => n397, ZN => 
                           n391);
   U758 : AND4_X1 port map( A1 => n392, A2 => n359, A3 => n358, A4 => n391, ZN 
                           => n385);
   U759 : OAI221_X1 port map( B1 => n387, B2 => n381, C1 => n387, C2 => n360, A
                           => n385, ZN => n443);
   U760 : OAI21_X1 port map( B1 => OP_B_26_port, B2 => n422, A => n421, ZN => 
                           n425);
   U761 : AOI211_X1 port map( C1 => OP_A_24_port, C2 => n416, A => n418, B => 
                           n425, ZN => n438);
   U762 : OAI21_X1 port map( B1 => OP_B_28_port, B2 => n411, A => n361, ZN => 
                           n415);
   U763 : NOR3_X1 port map( A1 => n427, A2 => n439, A3 => n415, ZN => n362);
   U764 : NAND2_X1 port map( A1 => n438, A2 => n362, ZN => n431);
   U765 : OAI21_X1 port map( B1 => n443, B2 => n431, A => OP_COMPARE_1_port, ZN
                           => n434);
   U766 : OAI22_X1 port map( A1 => n366, A2 => n365, B1 => n364, B2 => n363, ZN
                           => n376);
   U767 : NAND2_X1 port map( A1 => OP_B_4_port, A2 => n367, ZN => n369);
   U768 : OAI21_X1 port map( B1 => n370, B2 => n369, A => n368, ZN => n375);
   U769 : AOI21_X1 port map( B1 => OP_A_4_port, B2 => n1363, A => n370, ZN => 
                           n374);
   U770 : OAI21_X1 port map( B1 => OP_B_6_port, B2 => n371, A => n379, ZN => 
                           n372);
   U771 : INV_X1 port map( A => n372, ZN => n373);
   U772 : OAI221_X1 port map( B1 => n376, B2 => n375, C1 => n374, C2 => n375, A
                           => n373, ZN => n384);
   U773 : NOR2_X1 port map( A1 => OP_A_6_port, A2 => n377, ZN => n380);
   U774 : AOI21_X1 port map( B1 => n380, B2 => n379, A => n378, ZN => n383);
   U775 : INV_X1 port map( A => n381, ZN => n382);
   U776 : AOI21_X1 port map( B1 => n384, B2 => n383, A => n382, ZN => n386);
   U777 : OAI21_X1 port map( B1 => n387, B2 => n386, A => n385, ZN => n388);
   U778 : INV_X1 port map( A => n388, ZN => n442);
   U779 : OR2_X1 port map( A1 => OP_A_22_port, A2 => n389, ZN => n409);
   U780 : NAND2_X1 port map( A1 => n390, A2 => OP_B_18_port, ZN => n398);
   U781 : OAI211_X1 port map( C1 => n394, C2 => n393, A => n392, B => n391, ZN 
                           => n395);
   U782 : OAI211_X1 port map( C1 => n398, C2 => n397, A => n396, B => n395, ZN 
                           => n405);
   U783 : INV_X1 port map( A => n399, ZN => n400);
   U784 : OAI222_X1 port map( A1 => n401, A2 => n400, B1 => n401, B2 => 
                           OP_A_21_port, C1 => n400, C2 => OP_A_21_port, ZN => 
                           n404);
   U785 : OAI221_X1 port map( B1 => n405, B2 => n404, C1 => n403, C2 => n404, A
                           => n402, ZN => n406);
   U786 : OAI211_X1 port map( C1 => n409, C2 => n408, A => n407, B => n406, ZN 
                           => n454);
   U787 : INV_X1 port map( A => n454, ZN => n432);
   U788 : AOI21_X1 port map( B1 => n410, B2 => n449, A => n452, ZN => n430);
   U789 : NAND2_X1 port map( A1 => OP_B_28_port, A2 => n411, ZN => n413);
   U790 : OAI21_X1 port map( B1 => n414, B2 => n413, A => n412, ZN => n448);
   U791 : INV_X1 port map( A => n415, ZN => n447);
   U792 : OR2_X1 port map( A1 => OP_A_24_port, A2 => n416, ZN => n419);
   U793 : OAI21_X1 port map( B1 => n419, B2 => n418, A => n417, ZN => n420);
   U794 : INV_X1 port map( A => n420, ZN => n426);
   U795 : NAND3_X1 port map( A1 => OP_B_26_port, A2 => n422, A3 => n421, ZN => 
                           n423);
   U796 : OAI211_X1 port map( C1 => n426, C2 => n425, A => n424, B => n423, ZN 
                           => n446);
   U797 : NOR2_X1 port map( A1 => n427, A2 => n439, ZN => n428);
   U798 : OAI221_X1 port map( B1 => n448, B2 => n447, C1 => n448, C2 => n446, A
                           => n428, ZN => n429);
   U799 : OAI211_X1 port map( C1 => n432, C2 => n431, A => n430, B => n429, ZN 
                           => n433);
   U800 : AOI221_X1 port map( B1 => OP_COMPARE_2_port, B2 => n434, C1 => n442, 
                           C2 => n434, A => n433, ZN => n435);
   U801 : OAI21_X1 port map( B1 => n436, B2 => n435, A => OP_COMPARE_0_port, ZN
                           => n468);
   U802 : INV_X1 port map( A => n437, ZN => n466);
   U803 : INV_X1 port map( A => n438, ZN => n441);
   U804 : NOR2_X1 port map( A1 => n452, A2 => n439, ZN => n445);
   U805 : NAND2_X1 port map( A1 => n447, A2 => n445, ZN => n440);
   U806 : NOR2_X1 port map( A1 => n441, A2 => n440, ZN => n455);
   U807 : AOI21_X1 port map( B1 => n442, B2 => n455, A => OP_COMPARE_2_port, ZN
                           => n458);
   U808 : INV_X1 port map( A => n443, ZN => n444);
   U809 : AOI21_X1 port map( B1 => n444, B2 => n455, A => n459, ZN => n457);
   U810 : OAI221_X1 port map( B1 => n448, B2 => n447, C1 => n448, C2 => n446, A
                           => n445, ZN => n450);
   U811 : OAI211_X1 port map( C1 => n452, C2 => n451, A => n450, B => n449, ZN 
                           => n453);
   U812 : AOI21_X1 port map( B1 => n455, B2 => n454, A => n453, ZN => n456);
   U813 : OAI21_X1 port map( B1 => n458, B2 => n457, A => n456, ZN => n464);
   U814 : OAI211_X1 port map( C1 => n462, C2 => n461, A => n460, B => n459, ZN 
                           => n463);
   U815 : AOI21_X1 port map( B1 => n464, B2 => n463, A => OP_COMPARE_0_port, ZN
                           => n465);
   U816 : OAI21_X1 port map( B1 => n469, B2 => n466, A => n465, ZN => n467);
   U817 : OAI21_X1 port map( B1 => n469, B2 => n468, A => n467, ZN => n471);
   U818 : INV_X1 port map( A => N285, ZN => n470);
   U819 : AOI221_X1 port map( B1 => OP_COMPARE_3_port, B2 => n473, C1 => n472, 
                           C2 => n471, A => n470, ZN => n478);
   U820 : INV_X1 port map( A => N279, ZN => n1398);
   U821 : XOR2_X1 port map( A => n475, B => OP_Ci, Z => n476);
   U822 : NAND2_X1 port map( A1 => OP_LOGIC_1_port, A2 => n474, ZN => n1372);
   U823 : OAI22_X1 port map( A1 => n1398, A2 => n476, B1 => n1372, B2 => n475, 
                           ZN => n477);
   U824 : AOI211_X1 port map( C1 => n1367, C2 => n487, A => n478, B => n477, ZN
                           => n479);
   U825 : OAI211_X1 port map( C1 => n1159, C2 => n481, A => n480, B => n479, ZN
                           => Y(0));
   U826 : INV_X1 port map( A => n507, ZN => n482);
   U827 : AOI21_X1 port map( B1 => OP_B_1_port, B2 => C428_DATA4_1, A => n482, 
                           ZN => n484);
   U828 : OAI22_X1 port map( A1 => n1396, A2 => n484, B1 => n1139, B2 => n483, 
                           ZN => n486);
   U829 : AOI22_X1 port map( A1 => n542, A2 => OP_A_0_port, B1 => OP_A_1_port, 
                           B2 => n56, ZN => n920);
   U830 : OAI22_X1 port map( A1 => n920, A2 => n1061, B1 => n519, B2 => n1369, 
                           ZN => n485);
   U831 : AOI211_X1 port map( C1 => n1330, C2 => OP1(1), A => n486, B => n485, 
                           ZN => n504);
   U832 : AOI22_X1 port map( A1 => OP_B_0_port, A2 => OP_A_0_port, B1 => OP_Ci,
                           B2 => n487, ZN => n521);
   U833 : INV_X1 port map( A => n521, ZN => n489);
   U834 : INV_X1 port map( A => n505, ZN => n488);
   U835 : AOI221_X1 port map( B1 => n521, B2 => n505, C1 => n489, C2 => n488, A
                           => n1398, ZN => n501);
   U836 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n55, ZN => n1353);
   U837 : NAND2_X1 port map( A1 => n491, A2 => OP_A_26_port, ZN => n1226);
   U838 : NAND2_X1 port map( A1 => OP_A_27_port, A2 => n553, ZN => n1289);
   U839 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => n56, ZN => n1166);
   U840 : NAND4_X1 port map( A1 => n1353, A2 => n1226, A3 => n1289, A4 => n1166
                           , ZN => n791);
   U841 : NAND2_X1 port map( A1 => n491, A2 => OP_A_30_port, ZN => n1354);
   U842 : NAND2_X1 port map( A1 => OP_A_29_port, A2 => n56, ZN => n1290);
   U843 : OAI211_X1 port map( C1 => n575, C2 => n1370, A => n1354, B => n1290, 
                           ZN => n490);
   U844 : AOI21_X1 port map( B1 => OP_SHIFT, B2 => n55, A => n490, ZN => n1298)
                           ;
   U845 : INV_X1 port map( A => n1298, ZN => n797);
   U846 : AOI22_X1 port map( A1 => n855, A2 => n791, B1 => n510, B2 => n797, ZN
                           => n493);
   U847 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => n55, ZN => n1225);
   U848 : NAND2_X1 port map( A1 => n491, A2 => OP_A_22_port, ZN => n1098);
   U849 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => n553, ZN => n1169);
   U850 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => n56, ZN => n1033);
   U851 : NAND4_X1 port map( A1 => n1225, A2 => n1098, A3 => n1169, A4 => n1033
                           , ZN => n792);
   U852 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => n55, ZN => n1097);
   U853 : NAND2_X1 port map( A1 => n542, A2 => OP_A_18_port, ZN => n971);
   U854 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => n553, ZN => n1036);
   U855 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n56, ZN => n912);
   U856 : NAND4_X1 port map( A1 => n1097, A2 => n971, A3 => n1036, A4 => n912, 
                           ZN => n794);
   U857 : AOI22_X1 port map( A1 => n63, A2 => n792, B1 => n894, B2 => n794, ZN 
                           => n492);
   U858 : NAND2_X1 port map( A1 => n493, A2 => n492, ZN => n922);
   U859 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => n55, ZN => n738);
   U860 : NAND2_X1 port map( A1 => OP_A_7_port, A2 => n553, ZN => n693);
   U861 : NAND2_X1 port map( A1 => OP_A_5_port, A2 => n56, ZN => n494);
   U862 : NAND4_X1 port map( A1 => n738, A2 => n658, A3 => n693, A4 => n494, ZN
                           => n596);
   U863 : AOI22_X1 port map( A1 => OP_B_4_port, A2 => n922, B1 => n1358, B2 => 
                           n596, ZN => n499);
   U864 : NAND2_X1 port map( A1 => OP_A_4_port, A2 => n55, ZN => n656);
   U865 : NAND2_X1 port map( A1 => OP_A_1_port, A2 => n56, ZN => n495);
   U866 : OAI211_X1 port map( C1 => n575, C2 => n550, A => n656, B => n495, ZN 
                           => n497);
   U867 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n55, ZN => n970);
   U868 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => n56, ZN => n802);
   U869 : NAND2_X1 port map( A1 => OP_A_15_port, A2 => n553, ZN => n915);
   U870 : NAND4_X1 port map( A1 => n852, A2 => n970, A3 => n802, A4 => n915, ZN
                           => n609);
   U871 : INV_X1 port map( A => n609, ZN => n795);
   U872 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => n55, ZN => n850);
   U873 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => n553, ZN => n803);
   U874 : NAND2_X1 port map( A1 => OP_A_9_port, A2 => n56, ZN => n694);
   U875 : AND4_X1 port map( A1 => n850, A2 => n740, A3 => n803, A4 => n694, ZN 
                           => n699);
   U876 : OAI22_X1 port map( A1 => n795, A2 => n891, B1 => n699, B2 => n566, ZN
                           => n496);
   U877 : AOI221_X1 port map( B1 => n552, B2 => n1360, C1 => n497, C2 => n1360,
                           A => n496, ZN => n498);
   U878 : AOI21_X1 port map( B1 => n499, B2 => n498, A => n1159, ZN => n500);
   U879 : AOI211_X1 port map( C1 => n1367, C2 => n502, A => n501, B => n500, ZN
                           => n503);
   U880 : OAI211_X1 port map( C1 => n1372, C2 => n505, A => n504, B => n503, ZN
                           => Y(1));
   U881 : INV_X1 port map( A => n523, ZN => n522);
   U882 : AOI22_X1 port map( A1 => n506, A2 => n1245, B1 => n1344, B2 => n522, 
                           ZN => n533);
   U883 : INV_X1 port map( A => n1139, ZN => n1348);
   U884 : NAND2_X1 port map( A1 => OP_A_2_port, A2 => n56, ZN => n515);
   U885 : OAI211_X1 port map( C1 => n575, C2 => n549, A => n507, B => n515, ZN 
                           => n820);
   U886 : AOI22_X1 port map( A1 => n1348, A2 => OP2(2), B1 => n1228, B2 => n820
                           , ZN => n532);
   U887 : AOI22_X1 port map( A1 => OP1(2), A2 => n1330, B1 => n1367, B2 => n546
                           , ZN => n531);
   U888 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => n56, ZN => n816);
   U889 : NAND2_X1 port map( A1 => OP_A_16_port, A2 => n603, ZN => n938);
   U890 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n55, ZN => n1003);
   U891 : NAND4_X1 port map( A1 => n890, A2 => n816, A3 => n938, A4 => n1003, 
                           ZN => n841);
   U892 : INV_X1 port map( A => n841, ZN => n728);
   U893 : NAND2_X1 port map( A1 => OP_A_8_port, A2 => n603, ZN => n723);
   U894 : NAND2_X1 port map( A1 => OP_A_6_port, A2 => n56, ZN => n625);
   U895 : NAND2_X1 port map( A1 => OP_A_9_port, A2 => n55, ZN => n766);
   U896 : NAND4_X1 port map( A1 => n723, A2 => n625, A3 => n766, A4 => n675, ZN
                           => n618);
   U897 : NAND2_X1 port map( A1 => OP_A_12_port, A2 => n603, ZN => n818);
   U898 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => n56, ZN => n724);
   U899 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => n55, ZN => n888);
   U900 : NAND4_X1 port map( A1 => n818, A2 => n724, A3 => n769, A4 => n888, ZN
                           => n721);
   U901 : AOI22_X1 port map( A1 => n1358, A2 => n618, B1 => n1350, B2 => n721, 
                           ZN => n518);
   U902 : NAND2_X1 port map( A1 => OP_A_24_port, A2 => n603, ZN => n1206);
   U903 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => n56, ZN => n1056);
   U904 : NAND2_X1 port map( A1 => n542, A2 => OP_A_23_port, ZN => n1132);
   U905 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => n55, ZN => n1270);
   U906 : AND4_X1 port map( A1 => n1206, A2 => n1056, A3 => n1132, A4 => n1270,
                           ZN => n824);
   U907 : AOI22_X1 port map( A1 => OP_B_1_port, A2 => OP_SHIFT, B1 => 
                           OP_A_30_port, B2 => n56, ZN => n508);
   U908 : OAI21_X1 port map( B1 => n509, B2 => n1370, A => n508, ZN => n1328);
   U909 : NAND2_X1 port map( A1 => OP_A_20_port, A2 => n603, ZN => n1059);
   U910 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => n56, ZN => n935);
   U911 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => n55, ZN => n1131);
   U912 : NAND2_X1 port map( A1 => n542, A2 => OP_A_19_port, ZN => n1004);
   U913 : NAND4_X1 port map( A1 => n1059, A2 => n935, A3 => n1131, A4 => n1004,
                           ZN => n826);
   U914 : AOI22_X1 port map( A1 => n510, A2 => n1328, B1 => n894, B2 => n826, 
                           ZN => n513);
   U915 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => n56, ZN => n1203);
   U916 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n553, ZN => n1320);
   U917 : NAND2_X1 port map( A1 => n542, A2 => OP_A_27_port, ZN => n1271);
   U918 : NAND2_X1 port map( A1 => OP_A_29_port, A2 => n55, ZN => n511);
   U919 : NAND4_X1 port map( A1 => n1203, A2 => n1320, A3 => n1271, A4 => n511,
                           ZN => n837);
   U920 : NAND2_X1 port map( A1 => n855, A2 => n837, ZN => n512);
   U921 : OAI211_X1 port map( C1 => n824, C2 => n742, A => n513, B => n512, ZN 
                           => n934);
   U922 : NAND2_X1 port map( A1 => OP_A_4_port, A2 => n553, ZN => n627);
   U923 : INV_X1 port map( A => n580, ZN => n514);
   U924 : NAND2_X1 port map( A1 => OP_A_5_port, A2 => n55, ZN => n673);
   U925 : NAND4_X1 port map( A1 => n627, A2 => n515, A3 => n514, A4 => n673, ZN
                           => n516);
   U926 : AOI22_X1 port map( A1 => OP_B_4_port, A2 => n934, B1 => n1360, B2 => 
                           n516, ZN => n517);
   U927 : OAI211_X1 port map( C1 => n728, C2 => n891, A => n518, B => n517, ZN 
                           => n529);
   U928 : OAI21_X1 port map( B1 => n521, B2 => n520, A => n519, ZN => n547);
   U929 : INV_X1 port map( A => n547, ZN => n524);
   U930 : AOI221_X1 port map( B1 => n524, B2 => n523, C1 => n547, C2 => n522, A
                           => n1398, ZN => n528);
   U931 : AOI211_X1 port map( C1 => n526, C2 => n525, A => n537, B => n1396, ZN
                           => n527);
   U932 : AOI211_X1 port map( C1 => N284, C2 => n529, A => n528, B => n527, ZN 
                           => n530);
   U933 : NAND4_X1 port map( A1 => n533, A2 => n532, A3 => n531, A4 => n530, ZN
                           => Y(2));
   U934 : XNOR2_X1 port map( A => n535, B => n534, ZN => n536);
   U935 : XNOR2_X1 port map( A => n537, B => n536, ZN => n563);
   U936 : INV_X1 port map( A => n1396, ZN => n986);
   U937 : INV_X1 port map( A => n986, ZN => n1284);
   U938 : NAND2_X1 port map( A1 => OP_A_25_port, A2 => n553, ZN => n1227);
   U939 : NAND2_X1 port map( A1 => OP_A_23_port, A2 => n56, ZN => n1096);
   U940 : NAND2_X1 port map( A1 => OP_A_26_port, A2 => n55, ZN => n1287);
   U941 : NAND2_X1 port map( A1 => n542, A2 => OP_A_24_port, ZN => n1168);
   U942 : NAND4_X1 port map( A1 => n1227, A2 => n1096, A3 => n1287, A4 => n1168
                           , ZN => n863);
   U943 : NAND2_X1 port map( A1 => OP_A_29_port, A2 => n553, ZN => n1355);
   U944 : NAND2_X1 port map( A1 => OP_A_27_port, A2 => n56, ZN => n1224);
   U945 : NAND2_X1 port map( A1 => n542, A2 => OP_A_28_port, ZN => n1288);
   U946 : NAND3_X1 port map( A1 => n1355, A2 => n1224, A3 => n1288, ZN => n538)
                           ;
   U947 : AOI21_X1 port map( B1 => OP_A_30_port, B2 => n55, A => n538, ZN => 
                           n869);
   U948 : NOR2_X1 port map( A1 => n869, A2 => n741, ZN => n540);
   U949 : AOI22_X1 port map( A1 => n56, A2 => OP_A_31_port, B1 => OP_SHIFT, B2 
                           => n607, ZN => n1374);
   U950 : NAND2_X1 port map( A1 => OP_A_21_port, A2 => n553, ZN => n1099);
   U951 : NAND2_X1 port map( A1 => OP_A_19_port, A2 => n56, ZN => n969);
   U952 : NAND2_X1 port map( A1 => OP_A_22_port, A2 => n55, ZN => n1167);
   U953 : NAND2_X1 port map( A1 => n542, A2 => OP_A_20_port, ZN => n1035);
   U954 : NAND4_X1 port map( A1 => n1099, A2 => n969, A3 => n1167, A4 => n1035,
                           ZN => n865);
   U955 : INV_X1 port map( A => n865, ZN => n748);
   U956 : OAI22_X1 port map( A1 => n1374, A2 => n857, B1 => n748, B2 => n765, 
                           ZN => n539);
   U957 : NAND2_X1 port map( A1 => OP_A_9_port, A2 => n553, ZN => n737);
   U958 : NAND2_X1 port map( A1 => OP_A_7_port, A2 => n56, ZN => n655);
   U959 : NAND2_X1 port map( A1 => OP_A_10_port, A2 => n55, ZN => n801);
   U960 : NAND4_X1 port map( A1 => n737, A2 => n655, A3 => n801, A4 => n696, ZN
                           => n648);
   U961 : NAND2_X1 port map( A1 => OP_A_13_port, A2 => n553, ZN => n851);
   U962 : NAND2_X1 port map( A1 => OP_A_11_port, A2 => n56, ZN => n739);
   U963 : NAND2_X1 port map( A1 => OP_A_14_port, A2 => n55, ZN => n913);
   U964 : NAND4_X1 port map( A1 => n851, A2 => n739, A3 => n804, A4 => n913, ZN
                           => n644);
   U965 : AOI22_X1 port map( A1 => n1358, A2 => n648, B1 => n1350, B2 => n644, 
                           ZN => n545);
   U966 : NAND2_X1 port map( A1 => OP_A_5_port, A2 => n553, ZN => n657);
   U967 : NAND2_X1 port map( A1 => OP_A_3_port, A2 => n56, ZN => n541);
   U968 : NAND2_X1 port map( A1 => OP_A_6_port, A2 => n55, ZN => n695);
   U969 : NAND4_X1 port map( A1 => n657, A2 => n541, A3 => n695, A4 => n604, ZN
                           => n543);
   U970 : NAND2_X1 port map( A1 => OP_A_15_port, A2 => n56, ZN => n849);
   U971 : NAND2_X1 port map( A1 => OP_A_17_port, A2 => n553, ZN => n972);
   U972 : NAND2_X1 port map( A1 => OP_A_18_port, A2 => n55, ZN => n1034);
   U973 : NAND2_X1 port map( A1 => n542, A2 => OP_A_16_port, ZN => n914);
   U974 : NAND4_X1 port map( A1 => n849, A2 => n972, A3 => n1034, A4 => n914, 
                           ZN => n874);
   U975 : AOI22_X1 port map( A1 => n1360, A2 => n543, B1 => n1352, B2 => n874, 
                           ZN => n544);
   U976 : OAI211_X1 port map( C1 => n964, C2 => n1363, A => n545, B => n544, ZN
                           => n560);
   U977 : AOI22_X1 port map( A1 => OP_B_2_port, A2 => OP_A_2_port, B1 => n547, 
                           B2 => n546, ZN => n548);
   U978 : NOR2_X1 port map( A1 => n557, A2 => n548, ZN => n571);
   U979 : AOI211_X1 port map( C1 => n557, C2 => n548, A => n1398, B => n571, ZN
                           => n559);
   U980 : AOI22_X1 port map( A1 => n1348, A2 => OP2(3), B1 => n1347, B2 => 
                           OP1(3), ZN => n556);
   U981 : OAI22_X1 port map( A1 => n550, A2 => n607, B1 => n549, B2 => n577, ZN
                           => n551);
   U982 : AOI211_X1 port map( C1 => n553, C2 => OP_A_1_port, A => n552, B => 
                           n551, ZN => n966);
   U983 : INV_X1 port map( A => n966, ZN => n554);
   U984 : AOI22_X1 port map( A1 => OP_B_3_port, A2 => n1367, B1 => n1228, B2 =>
                           n554, ZN => n555);
   U985 : OAI211_X1 port map( C1 => n557, C2 => n1372, A => n556, B => n555, ZN
                           => n558);
   U986 : AOI211_X1 port map( C1 => N284, C2 => n560, A => n559, B => n558, ZN 
                           => n562);
   U987 : OAI221_X1 port map( B1 => n1367, B2 => OP_B_3_port, C1 => n1367, C2 
                           => n1245, A => OP_A_3_port, ZN => n561);
   U988 : OAI211_X1 port map( C1 => n563, C2 => n1284, A => n562, B => n561, ZN
                           => Y(3));
   U989 : NAND2_X1 port map( A1 => n1352, A2 => N284, ZN => n868);
   U990 : INV_X1 port map( A => n868, ZN => n838);
   U991 : AOI211_X1 port map( C1 => n565, C2 => intadd_0_SUM_0_port, A => n564,
                           B => n1396, ZN => n568);
   U992 : NOR2_X1 port map( A1 => n1159, A2 => n566, ZN => n864);
   U993 : INV_X1 port map( A => n864, ZN => n823);
   U994 : NOR2_X1 port map( A1 => n1159, A2 => n899, ZN => n866);
   U995 : INV_X1 port map( A => n866, ZN => n727);
   U996 : OAI22_X1 port map( A1 => n771, A2 => n823, B1 => n681, B2 => n727, ZN
                           => n567);
   U997 : AOI211_X1 port map( C1 => n838, C2 => n777, A => n568, B => n567, ZN 
                           => n589);
   U998 : INV_X1 port map( A => n573, ZN => n572);
   U999 : NAND2_X1 port map( A1 => OP_B_4_port, A2 => N284, ZN => n764);
   U1000 : INV_X1 port map( A => n764, ZN => n744);
   U1001 : AOI22_X1 port map( A1 => n855, A2 => n1265, B1 => n62, B2 => n781, 
                           ZN => n569);
   U1002 : INV_X1 port map( A => OP_SHIFT, ZN => n1158);
   U1003 : NOR2_X1 port map( A1 => n857, A2 => n1158, ZN => n660);
   U1004 : INV_X1 port map( A => n660, ZN => n623);
   U1005 : OAI211_X1 port map( C1 => n784, C2 => n765, A => n569, B => n623, ZN
                           => n1008);
   U1006 : AOI22_X1 port map( A1 => n1344, A2 => n572, B1 => n744, B2 => n1008,
                           ZN => n588);
   U1007 : INV_X1 port map( A => n570, ZN => n598);
   U1008 : AOI22_X1 port map( A1 => n1245, A2 => n598, B1 => n1367, B2 => n597,
                           ZN => n587);
   U1009 : AOI21_X1 port map( B1 => OP_A_3_port, B2 => OP_B_3_port, A => n571, 
                           ZN => n574);
   U1010 : INV_X1 port map( A => n574, ZN => n599);
   U1011 : AOI221_X1 port map( B1 => n574, B2 => n573, C1 => n599, C2 => n572, 
                           A => n1398, ZN => n585);
   U1012 : OAI22_X1 port map( A1 => n578, A2 => n577, B1 => n576, B2 => n575, 
                           ZN => n579);
   U1013 : AOI211_X1 port map( C1 => n56, C2 => OP_A_4_port, A => n580, B => 
                           n579, ZN => n892);
   U1014 : AOI22_X1 port map( A1 => OP_B_2_port, A2 => n895, B1 => n892, B2 => 
                           n581, ZN => n770);
   U1015 : NAND2_X1 port map( A1 => n770, A2 => n1160, ZN => n1011);
   U1016 : NAND2_X1 port map( A1 => n1363, A2 => n1366, ZN => n885);
   U1017 : NOR2_X1 port map( A1 => OP_B_4_port, A2 => n1159, ZN => n1252);
   U1018 : NAND2_X1 port map( A1 => n894, A2 => n1252, ZN => n1373);
   U1019 : INV_X1 port map( A => n1373, ZN => n1329);
   U1020 : AOI22_X1 port map( A1 => n1330, A2 => OP1(4), B1 => n1329, B2 => 
                           n582, ZN => n583);
   U1021 : OAI21_X1 port map( B1 => n1011, B2 => n885, A => n583, ZN => n584);
   U1022 : AOI211_X1 port map( C1 => n1348, C2 => OP2(4), A => n585, B => n584,
                           ZN => n586);
   U1023 : NAND4_X1 port map( A1 => n589, A2 => n588, A3 => n587, A4 => n586, 
                           ZN => Y(4));
   U1024 : XNOR2_X1 port map( A => n591, B => n590, ZN => n592);
   U1025 : XNOR2_X1 port map( A => intadd_0_SUM_1_port, B => n592, ZN => n617);
   U1026 : INV_X1 port map( A => n794, ZN => n703);
   U1027 : OAI22_X1 port map( A1 => n703, A2 => n868, B1 => n699, B2 => n727, 
                           ZN => n595);
   U1028 : OAI22_X1 port map( A1 => n593, A2 => n1369, B1 => n1372, B2 => n600,
                           ZN => n594);
   U1029 : AOI211_X1 port map( C1 => n1329, C2 => n596, A => n595, B => n594, 
                           ZN => n616);
   U1030 : OAI21_X1 port map( B1 => n599, B2 => n598, A => n597, ZN => n601);
   U1031 : INV_X1 port map( A => n601, ZN => n633);
   U1032 : INV_X1 port map( A => n600, ZN => n602);
   U1033 : AOI221_X1 port map( B1 => n633, B2 => n602, C1 => n601, C2 => n600, 
                           A => n1398, ZN => n614);
   U1034 : INV_X1 port map( A => n885, ZN => n743);
   U1035 : AOI22_X1 port map( A1 => OP_A_3_port, A2 => n603, B1 => OP_A_2_port,
                           B2 => n55, ZN => n605);
   U1036 : OAI211_X1 port map( C1 => n607, C2 => n606, A => n605, B => n604, ZN
                           => n919);
   U1037 : INV_X1 port map( A => n919, ZN => n697);
   U1038 : OAI22_X1 port map( A1 => n697, A2 => n765, B1 => n920, B2 => n742, 
                           ZN => n1029);
   U1039 : AOI22_X1 port map( A1 => n1330, A2 => OP1(5), B1 => n743, B2 => 
                           n1029, ZN => n611);
   U1040 : AOI22_X1 port map( A1 => n853, A2 => n791, B1 => n894, B2 => n792, 
                           ZN => n608);
   U1041 : OAI211_X1 port map( C1 => n1298, C2 => n741, A => n608, B => n623, 
                           ZN => n1038);
   U1042 : AOI22_X1 port map( A1 => n744, A2 => n1038, B1 => n864, B2 => n609, 
                           ZN => n610);
   U1043 : OAI211_X1 port map( C1 => n1139, C2 => n612, A => n611, B => n610, 
                           ZN => n613);
   U1044 : AOI211_X1 port map( C1 => n1367, C2 => n632, A => n614, B => n613, 
                           ZN => n615);
   U1045 : OAI211_X1 port map( C1 => n1284, C2 => n617, A => n616, B => n615, 
                           ZN => Y(5));
   U1046 : INV_X1 port map( A => n636, ZN => n634);
   U1047 : AOI22_X1 port map( A1 => n1329, A2 => n618, B1 => n1344, B2 => n634,
                           ZN => n640);
   U1048 : AOI211_X1 port map( C1 => n620, C2 => intadd_1_SUM_0_port, A => n619
                           , B => n1396, ZN => n622);
   U1049 : OAI22_X1 port map( A1 => n651, A2 => n1368, B1 => n728, B2 => n823, 
                           ZN => n621);
   U1050 : AOI211_X1 port map( C1 => n866, C2 => n721, A => n622, B => n621, ZN
                           => n639);
   U1051 : AOI22_X1 port map( A1 => n855, A2 => n1328, B1 => n63, B2 => n837, 
                           ZN => n624);
   U1052 : OAI211_X1 port map( C1 => n824, C2 => n765, A => n624, B => n623, ZN
                           => n1065);
   U1053 : NAND4_X1 port map( A1 => n628, A2 => n627, A3 => n626, A4 => n625, 
                           ZN => n940);
   U1054 : AOI22_X1 port map( A1 => n62, A2 => n820, B1 => n894, B2 => n940, ZN
                           => n1062);
   U1055 : AOI22_X1 port map( A1 => n1348, A2 => OP2(6), B1 => n1330, B2 => 
                           OP1(6), ZN => n629);
   U1056 : OAI21_X1 port map( B1 => n1062, B2 => n885, A => n629, ZN => n631);
   U1057 : INV_X1 port map( A => n826, ZN => n729);
   U1058 : OAI22_X1 port map( A1 => n729, A2 => n868, B1 => n649, B2 => n1369, 
                           ZN => n630);
   U1059 : AOI211_X1 port map( C1 => n744, C2 => n1065, A => n631, B => n630, 
                           ZN => n638);
   U1060 : AOI22_X1 port map( A1 => OP_B_5_port, A2 => OP_A_5_port, B1 => n633,
                           B2 => n632, ZN => n650);
   U1061 : INV_X1 port map( A => n650, ZN => n635);
   U1062 : OAI221_X1 port map( B1 => n650, B2 => n636, C1 => n635, C2 => n634, 
                           A => N279, ZN => n637);
   U1063 : NAND4_X1 port map( A1 => n640, A2 => n639, A3 => n638, A4 => n637, 
                           ZN => Y(6));
   U1064 : XNOR2_X1 port map( A => n642, B => n641, ZN => n643);
   U1065 : XNOR2_X1 port map( A => intadd_1_SUM_1_port, B => n643, ZN => n669);
   U1066 : INV_X1 port map( A => n644, ZN => n747);
   U1067 : OAI22_X1 port map( A1 => n748, A2 => n868, B1 => n747, B2 => n727, 
                           ZN => n647);
   U1068 : OAI22_X1 port map( A1 => n645, A2 => n1369, B1 => n1372, B2 => n653,
                           ZN => n646);
   U1069 : AOI211_X1 port map( C1 => n1329, C2 => n648, A => n647, B => n646, 
                           ZN => n668);
   U1070 : OAI21_X1 port map( B1 => n651, B2 => n650, A => n649, ZN => n677);
   U1071 : INV_X1 port map( A => n677, ZN => n654);
   U1072 : INV_X1 port map( A => n653, ZN => n652);
   U1073 : AOI221_X1 port map( B1 => n654, B2 => n653, C1 => n677, C2 => n652, 
                           A => n1398, ZN => n666);
   U1074 : NAND4_X1 port map( A1 => n658, A2 => n657, A3 => n656, A4 => n655, 
                           ZN => n854);
   U1075 : INV_X1 port map( A => n854, ZN => n963);
   U1076 : OAI22_X1 port map( A1 => n963, A2 => n765, B1 => n966, B2 => n742, 
                           ZN => n1100);
   U1077 : AOI22_X1 port map( A1 => n1330, A2 => OP1(7), B1 => n743, B2 => 
                           n1100, ZN => n663);
   U1078 : OAI22_X1 port map( A1 => n1374, A2 => n741, B1 => n869, B2 => n742, 
                           ZN => n659);
   U1079 : AOI211_X1 port map( C1 => n894, C2 => n863, A => n660, B => n659, ZN
                           => n1107);
   U1080 : INV_X1 port map( A => n1107, ZN => n661);
   U1081 : AOI22_X1 port map( A1 => n744, A2 => n661, B1 => n864, B2 => n874, 
                           ZN => n662);
   U1082 : OAI211_X1 port map( C1 => n1139, C2 => n664, A => n663, B => n662, 
                           ZN => n665);
   U1083 : AOI211_X1 port map( C1 => n1367, C2 => n678, A => n666, B => n665, 
                           ZN => n667);
   U1084 : OAI211_X1 port map( C1 => n1284, C2 => n669, A => n668, B => n667, 
                           ZN => Y(7));
   U1085 : AOI22_X1 port map( A1 => n63, A2 => n1265, B1 => n894, B2 => n781, 
                           ZN => n670);
   U1086 : OAI21_X1 port map( B1 => n1160, B2 => n1158, A => n670, ZN => n1135)
                           ;
   U1087 : AOI22_X1 port map( A1 => n744, A2 => n1135, B1 => n1367, B2 => n671,
                           ZN => n690);
   U1088 : INV_X1 port map( A => n711, ZN => n676);
   U1089 : NAND4_X1 port map( A1 => n675, A2 => n674, A3 => n673, A4 => n672, 
                           ZN => n1006);
   U1090 : INV_X1 port map( A => n1006, ZN => n905);
   U1091 : OAI222_X1 port map( A1 => n895, A2 => n741, B1 => n765, B2 => n905, 
                           C1 => n742, C2 => n892, ZN => n1134);
   U1092 : AOI22_X1 port map( A1 => n676, A2 => n1245, B1 => n743, B2 => n1134,
                           ZN => n689);
   U1093 : AOI22_X1 port map( A1 => OP_B_7_port, A2 => OP_A_7_port, B1 => n678,
                           B2 => n677, ZN => n712);
   U1094 : NOR2_X1 port map( A1 => n712, A2 => n680, ZN => n679);
   U1095 : AOI211_X1 port map( C1 => n712, C2 => n680, A => n1398, B => n679, 
                           ZN => n687);
   U1096 : OAI22_X1 port map( A1 => n681, A2 => n1373, B1 => n680, B2 => n1372,
                           ZN => n686);
   U1097 : AOI22_X1 port map( A1 => n1348, A2 => OP2(8), B1 => n1330, B2 => 
                           OP1(8), ZN => n684);
   U1098 : OAI22_X1 port map( A1 => n784, A2 => n868, B1 => n771, B2 => n727, 
                           ZN => n682);
   U1099 : AOI21_X1 port map( B1 => n864, B2 => n777, A => n682, ZN => n683);
   U1100 : OAI211_X1 port map( C1 => intadd_2_SUM_0_port, C2 => n1284, A => 
                           n684, B => n683, ZN => n685);
   U1101 : NOR3_X1 port map( A1 => n687, A2 => n686, A3 => n685, ZN => n688);
   U1102 : NAND3_X1 port map( A1 => n690, A2 => n689, A3 => n688, ZN => Y(8));
   U1103 : OAI22_X1 port map( A1 => intadd_2_SUM_1_port, A2 => n1284, B1 => 
                           n1139, B2 => n691, ZN => n692);
   U1104 : AOI21_X1 port map( B1 => n702, B2 => n1344, A => n692, ZN => n710);
   U1105 : NAND4_X1 port map( A1 => n696, A2 => n695, A3 => n694, A4 => n693, 
                           ZN => n1037);
   U1106 : INV_X1 port map( A => n1037, ZN => n931);
   U1107 : OAI222_X1 port map( A1 => n742, A2 => n697, B1 => n765, B2 => n931, 
                           C1 => n741, C2 => n920, ZN => n1161);
   U1108 : AOI22_X1 port map( A1 => n1330, A2 => OP1(9), B1 => n743, B2 => 
                           n1161, ZN => n709);
   U1109 : NOR2_X1 port map( A1 => n1158, A2 => n764, ZN => n1121);
   U1110 : INV_X1 port map( A => n1121, ZN => n1109);
   U1111 : NOR2_X1 port map( A1 => n1160, A2 => n1109, ZN => n753);
   U1112 : INV_X1 port map( A => n698, ZN => n713);
   U1113 : OAI22_X1 port map( A1 => n699, A2 => n1373, B1 => n713, B2 => n1369,
                           ZN => n700);
   U1114 : AOI211_X1 port map( C1 => n838, C2 => n792, A => n753, B => n700, ZN
                           => n708);
   U1115 : AOI21_X1 port map( B1 => n712, B2 => n711, A => n715, ZN => n701);
   U1116 : XOR2_X1 port map( A => n702, B => n701, Z => n706);
   U1117 : OAI22_X1 port map( A1 => n703, A2 => n823, B1 => n714, B2 => n1368, 
                           ZN => n705);
   U1118 : AOI22_X1 port map( A1 => n853, A2 => n797, B1 => n894, B2 => n791, 
                           ZN => n1174);
   U1119 : OAI22_X1 port map( A1 => n1174, A2 => n764, B1 => n795, B2 => n727, 
                           ZN => n704);
   U1120 : AOI211_X1 port map( C1 => n706, C2 => N279, A => n705, B => n704, ZN
                           => n707);
   U1121 : NAND4_X1 port map( A1 => n710, A2 => n709, A3 => n708, A4 => n707, 
                           ZN => Y(9));
   U1122 : NAND2_X1 port map( A1 => n713, A2 => n711, ZN => n718);
   U1123 : INV_X1 port map( A => n712, ZN => n717);
   U1124 : OAI21_X1 port map( B1 => n715, B2 => n714, A => n713, ZN => n716);
   U1125 : OAI21_X1 port map( B1 => n718, B2 => n717, A => n716, ZN => n756);
   U1126 : XNOR2_X1 port map( A => n719, B => n756, ZN => n736);
   U1127 : NOR2_X1 port map( A1 => OP_A_10_port, A2 => OP_B_10_port, ZN => n757
                           );
   U1128 : OAI22_X1 port map( A1 => n757, A2 => n1368, B1 => n1372, B2 => n719,
                           ZN => n720);
   U1129 : AOI211_X1 port map( C1 => n1329, C2 => n721, A => n753, B => n720, 
                           ZN => n735);
   U1130 : AOI22_X1 port map( A1 => n1348, A2 => OP2(10), B1 => n1347, B2 => 
                           OP1(10), ZN => n722);
   U1131 : OAI21_X1 port map( B1 => n755, B2 => n1369, A => n722, ZN => n733);
   U1132 : OAI22_X1 port map( A1 => n824, A2 => n868, B1 => intadd_2_SUM_2_port
                           , B2 => n1284, ZN => n732);
   U1133 : NAND4_X1 port map( A1 => n726, A2 => n725, A3 => n724, A4 => n723, 
                           ZN => n939);
   U1134 : AOI222_X1 port map( A1 => n820, A2 => n855, B1 => n940, B2 => n853, 
                           C1 => n939, C2 => n894, ZN => n1212);
   U1135 : AOI22_X1 port map( A1 => n62, A2 => n1328, B1 => n894, B2 => n837, 
                           ZN => n1182);
   U1136 : OAI22_X1 port map( A1 => n1212, A2 => n885, B1 => n1182, B2 => n764,
                           ZN => n731);
   U1137 : OAI22_X1 port map( A1 => n729, A2 => n823, B1 => n728, B2 => n727, 
                           ZN => n730);
   U1138 : NOR4_X1 port map( A1 => n733, A2 => n732, A3 => n731, A4 => n730, ZN
                           => n734);
   U1139 : OAI211_X1 port map( C1 => n1398, C2 => n736, A => n735, B => n734, 
                           ZN => Y(10));
   U1140 : AOI22_X1 port map( A1 => n866, A2 => n874, B1 => n838, B2 => n863, 
                           ZN => n763);
   U1141 : OAI22_X1 port map( A1 => n1374, A2 => n742, B1 => n869, B2 => n765, 
                           ZN => n1251);
   U1142 : NAND4_X1 port map( A1 => n740, A2 => n739, A3 => n738, A4 => n737, 
                           ZN => n973);
   U1143 : INV_X1 port map( A => n973, ZN => n1112);
   U1144 : OAI222_X1 port map( A1 => n742, A2 => n963, B1 => n765, B2 => n1112,
                           C1 => n741, C2 => n966, ZN => n1243);
   U1145 : AOI22_X1 port map( A1 => n744, A2 => n1251, B1 => n743, B2 => n1243,
                           ZN => n762);
   U1146 : AOI22_X1 port map( A1 => OP1(11), A2 => n1330, B1 => n1367, B2 => 
                           n773, ZN => n746);
   U1147 : NAND2_X1 port map( A1 => n1348, A2 => OP2(11), ZN => n745);
   U1148 : OAI211_X1 port map( C1 => intadd_2_SUM_3_port, C2 => n1284, A => 
                           n746, B => n745, ZN => n752);
   U1149 : OAI22_X1 port map( A1 => n748, A2 => n823, B1 => n747, B2 => n1373, 
                           ZN => n751);
   U1150 : OAI22_X1 port map( A1 => n749, A2 => n1369, B1 => n1372, B2 => n754,
                           ZN => n750);
   U1151 : NOR4_X1 port map( A1 => n753, A2 => n752, A3 => n751, A4 => n750, ZN
                           => n761);
   U1152 : INV_X1 port map( A => n754, ZN => n759);
   U1153 : OAI21_X1 port map( B1 => n757, B2 => n756, A => n755, ZN => n774);
   U1154 : AOI21_X1 port map( B1 => n759, B2 => n774, A => n1398, ZN => n758);
   U1155 : OAI21_X1 port map( B1 => n759, B2 => n774, A => n758, ZN => n760);
   U1156 : NAND4_X1 port map( A1 => n763, A2 => n762, A3 => n761, A4 => n760, 
                           ZN => Y(11));
   U1157 : NOR2_X1 port map( A1 => n765, A2 => n764, ZN => n876);
   U1158 : NAND4_X1 port map( A1 => n769, A2 => n768, A3 => n767, A4 => n766, 
                           ZN => n1119);
   U1159 : AOI222_X1 port map( A1 => n1006, A2 => n62, B1 => OP_B_3_port, B2 =>
                           n770, C1 => n1119, C2 => n894, ZN => n1278);
   U1160 : OAI22_X1 port map( A1 => n1278, A2 => n885, B1 => n771, B2 => n1373,
                           ZN => n772);
   U1161 : AOI21_X1 port map( B1 => n876, B2 => n1265, A => n772, ZN => n790);
   U1162 : AOI22_X1 port map( A1 => OP_A_11_port, A2 => OP_B_11_port, B1 => 
                           n774, B2 => n773, ZN => n828);
   U1163 : NOR2_X1 port map( A1 => n828, A2 => n779, ZN => n775);
   U1164 : AOI211_X1 port map( C1 => n828, C2 => n779, A => n1398, B => n775, 
                           ZN => n788);
   U1165 : OAI22_X1 port map( A1 => intadd_2_SUM_4_port, A2 => n1284, B1 => 
                           n1139, B2 => n776, ZN => n787);
   U1166 : AOI22_X1 port map( A1 => n1330, A2 => OP1(12), B1 => n866, B2 => 
                           n777, ZN => n778);
   U1167 : OAI21_X1 port map( B1 => n779, B2 => n1372, A => n778, ZN => n786);
   U1168 : AOI22_X1 port map( A1 => n838, A2 => n781, B1 => n1367, B2 => n780, 
                           ZN => n783);
   U1169 : NOR2_X1 port map( A1 => n894, A2 => n1109, ZN => n861);
   U1170 : INV_X1 port map( A => n861, ZN => n782);
   U1171 : OAI211_X1 port map( C1 => n784, C2 => n823, A => n783, B => n782, ZN
                           => n785);
   U1172 : NOR4_X1 port map( A1 => n788, A2 => n787, A3 => n786, A4 => n785, ZN
                           => n789);
   U1173 : OAI211_X1 port map( C1 => n827, C2 => n1369, A => n790, B => n789, 
                           ZN => Y(12));
   U1174 : AOI22_X1 port map( A1 => n864, A2 => n792, B1 => n838, B2 => n791, 
                           ZN => n815);
   U1175 : AOI22_X1 port map( A1 => n866, A2 => n794, B1 => n1367, B2 => n793, 
                           ZN => n814);
   U1176 : OAI22_X1 port map( A1 => n795, A2 => n1373, B1 => n829, B2 => n1369,
                           ZN => n796);
   U1177 : AOI211_X1 port map( C1 => n876, C2 => n797, A => n861, B => n796, ZN
                           => n813);
   U1178 : INV_X1 port map( A => n798, ZN => n807);
   U1179 : AOI21_X1 port map( B1 => n828, B2 => n827, A => n830, ZN => n799);
   U1180 : XOR2_X1 port map( A => n807, B => n799, Z => n811);
   U1181 : OAI22_X1 port map( A1 => intadd_2_SUM_5_port, A2 => n1284, B1 => 
                           n1139, B2 => n800, ZN => n810);
   U1182 : NAND4_X1 port map( A1 => n804, A2 => n803, A3 => n802, A4 => n801, 
                           ZN => n1170);
   U1183 : AOI22_X1 port map( A1 => n855, A2 => n919, B1 => n853, B2 => n1037, 
                           ZN => n805);
   U1184 : OAI21_X1 port map( B1 => n920, B2 => n857, A => n805, ZN => n806);
   U1185 : AOI21_X1 port map( B1 => n894, B2 => n1170, A => n806, ZN => n1295);
   U1186 : AOI22_X1 port map( A1 => n807, A2 => n1344, B1 => n1347, B2 => 
                           OP1(13), ZN => n808);
   U1187 : OAI21_X1 port map( B1 => n1295, B2 => n885, A => n808, ZN => n809);
   U1188 : AOI211_X1 port map( C1 => n811, C2 => N279, A => n810, B => n809, ZN
                           => n812);
   U1189 : NAND4_X1 port map( A1 => n815, A2 => n814, A3 => n813, A4 => n812, 
                           ZN => Y(13));
   U1190 : NOR2_X1 port map( A1 => OP_A_14_port, A2 => OP_B_14_port, ZN => n872
                           );
   U1191 : NAND4_X1 port map( A1 => n819, A2 => n818, A3 => n817, A4 => n816, 
                           ZN => n1207);
   U1192 : INV_X1 port map( A => n820, ZN => n932);
   U1193 : AOI22_X1 port map( A1 => n855, A2 => n940, B1 => n62, B2 => n939, ZN
                           => n821);
   U1194 : OAI21_X1 port map( B1 => n932, B2 => n857, A => n821, ZN => n822);
   U1195 : AOI21_X1 port map( B1 => n894, B2 => n1207, A => n822, ZN => n1326);
   U1196 : OAI22_X1 port map( A1 => n824, A2 => n823, B1 => n1326, B2 => n885, 
                           ZN => n825);
   U1197 : AOI21_X1 port map( B1 => n866, B2 => n826, A => n825, ZN => n848);
   U1198 : INV_X1 port map( A => n835, ZN => n842);
   U1199 : NAND2_X1 port map( A1 => n829, A2 => n827, ZN => n834);
   U1200 : INV_X1 port map( A => n828, ZN => n833);
   U1201 : OAI21_X1 port map( B1 => n831, B2 => n830, A => n829, ZN => n832);
   U1202 : OAI21_X1 port map( B1 => n834, B2 => n833, A => n832, ZN => n871);
   U1203 : INV_X1 port map( A => n871, ZN => n836);
   U1204 : AOI221_X1 port map( B1 => n842, B2 => n836, C1 => n835, C2 => n871, 
                           A => n1398, ZN => n846);
   U1205 : AOI22_X1 port map( A1 => n1348, A2 => OP2(14), B1 => n1347, B2 => 
                           OP1(14), ZN => n840);
   U1206 : AOI22_X1 port map( A1 => n838, A2 => n837, B1 => n876, B2 => n1328, 
                           ZN => n839);
   U1207 : OAI211_X1 port map( C1 => intadd_2_SUM_6_port, C2 => n1284, A => 
                           n840, B => n839, ZN => n845);
   U1208 : AOI22_X1 port map( A1 => n842, A2 => n1344, B1 => n1329, B2 => n841,
                           ZN => n843);
   U1209 : OAI21_X1 port map( B1 => n870, B2 => n1369, A => n843, ZN => n844);
   U1210 : NOR4_X1 port map( A1 => n861, A2 => n846, A3 => n845, A4 => n844, ZN
                           => n847);
   U1211 : OAI211_X1 port map( C1 => n872, C2 => n1368, A => n848, B => n847, 
                           ZN => Y(14));
   U1212 : NAND4_X1 port map( A1 => n852, A2 => n851, A3 => n850, A4 => n849, 
                           ZN => n1229);
   U1213 : AOI22_X1 port map( A1 => n855, A2 => n854, B1 => n63, B2 => n973, ZN
                           => n856);
   U1214 : OAI21_X1 port map( B1 => n966, B2 => n857, A => n856, ZN => n858);
   U1215 : AOI21_X1 port map( B1 => n894, B2 => n1229, A => n858, ZN => n1364);
   U1216 : OAI22_X1 port map( A1 => intadd_2_SUM_7_port, A2 => n1284, B1 => 
                           n1139, B2 => n859, ZN => n860);
   U1217 : AOI211_X1 port map( C1 => n1330, C2 => OP1(15), A => n861, B => n860
                           , ZN => n884);
   U1218 : INV_X1 port map( A => n862, ZN => n901);
   U1219 : AOI22_X1 port map( A1 => n866, A2 => n865, B1 => n864, B2 => n863, 
                           ZN => n867);
   U1220 : OAI21_X1 port map( B1 => n869, B2 => n868, A => n867, ZN => n882);
   U1221 : OAI21_X1 port map( B1 => n872, B2 => n871, A => n870, ZN => n902);
   U1222 : XNOR2_X1 port map( A => n873, B => n902, ZN => n880);
   U1223 : AOI22_X1 port map( A1 => n1329, A2 => n874, B1 => n1344, B2 => n873,
                           ZN => n879);
   U1224 : INV_X1 port map( A => n1374, ZN => n875);
   U1225 : AOI22_X1 port map( A1 => n877, A2 => n1245, B1 => n876, B2 => n875, 
                           ZN => n878);
   U1226 : OAI211_X1 port map( C1 => n1398, C2 => n880, A => n879, B => n878, 
                           ZN => n881);
   U1227 : AOI211_X1 port map( C1 => n1367, C2 => n901, A => n882, B => n881, 
                           ZN => n883);
   U1228 : OAI211_X1 port map( C1 => n1364, C2 => n885, A => n884, B => n883, 
                           ZN => Y(15));
   U1229 : AOI22_X1 port map( A1 => n1348, A2 => OP2(16), B1 => n1347, B2 => 
                           OP1(16), ZN => n911);
   U1230 : OAI22_X1 port map( A1 => intadd_2_SUM_8_port, A2 => n1284, B1 => 
                           n949, B2 => n1369, ZN => n886);
   U1231 : NOR2_X1 port map( A1 => n1121, A2 => n886, ZN => n910);
   U1232 : NAND4_X1 port map( A1 => n890, A2 => n889, A3 => n888, A4 => n887, 
                           ZN => n1268);
   U1233 : INV_X1 port map( A => n1268, ZN => n893);
   U1234 : NOR2_X1 port map( A1 => n900, A2 => n891, ZN => n1230);
   U1235 : INV_X1 port map( A => n1230, ZN => n1111);
   U1236 : OAI22_X1 port map( A1 => n893, A2 => n1061, B1 => n892, B2 => n1111,
                           ZN => n897);
   U1237 : NOR2_X1 port map( A1 => n900, A2 => n1363, ZN => n1244);
   U1238 : NAND2_X1 port map( A1 => n894, A2 => n1244, ZN => n965);
   U1239 : OAI22_X1 port map( A1 => n952, A2 => n1368, B1 => n965, B2 => n895, 
                           ZN => n896);
   U1240 : AOI211_X1 port map( C1 => n1252, C2 => n898, A => n897, B => n896, 
                           ZN => n909);
   U1241 : NOR2_X1 port map( A1 => n900, A2 => n899, ZN => n1242);
   U1242 : AOI22_X1 port map( A1 => OP_A_15_port, A2 => OP_B_15_port, B1 => 
                           n902, B2 => n901, ZN => n950);
   U1243 : NOR2_X1 port map( A1 => n950, A2 => n904, ZN => n903);
   U1244 : AOI211_X1 port map( C1 => n950, C2 => n904, A => n1398, B => n903, 
                           ZN => n907);
   U1245 : NAND2_X1 port map( A1 => n1350, A2 => n1366, ZN => n1233);
   U1246 : OAI22_X1 port map( A1 => n905, A2 => n1233, B1 => n904, B2 => n1372,
                           ZN => n906);
   U1247 : AOI211_X1 port map( C1 => n1242, C2 => n1119, A => n907, B => n906, 
                           ZN => n908);
   U1248 : NAND4_X1 port map( A1 => n911, A2 => n910, A3 => n909, A4 => n908, 
                           ZN => Y(16));
   U1249 : NAND4_X1 port map( A1 => n915, A2 => n914, A3 => n913, A4 => n912, 
                           ZN => n1285);
   U1250 : AOI22_X1 port map( A1 => n918, A2 => n1344, B1 => n1228, B2 => n1285
                           , ZN => n930);
   U1251 : AOI22_X1 port map( A1 => n1348, A2 => OP2(17), B1 => n1347, B2 => 
                           OP1(17), ZN => n916);
   U1252 : OAI211_X1 port map( C1 => intadd_2_SUM_9_port, C2 => n1284, A => 
                           n916, B => n1109, ZN => n927);
   U1253 : AOI21_X1 port map( B1 => n950, B2 => n949, A => n952, ZN => n917);
   U1254 : XNOR2_X1 port map( A => n918, B => n917, ZN => n925);
   U1255 : AOI22_X1 port map( A1 => n1230, A2 => n919, B1 => n1242, B2 => n1170
                           , ZN => n924);
   U1256 : OAI22_X1 port map( A1 => n920, A2 => n965, B1 => n953, B2 => n1368, 
                           ZN => n921);
   U1257 : AOI21_X1 port map( B1 => n1252, B2 => n922, A => n921, ZN => n923);
   U1258 : OAI211_X1 port map( C1 => n1398, C2 => n925, A => n924, B => n923, 
                           ZN => n926);
   U1259 : AOI211_X1 port map( C1 => n928, C2 => n1245, A => n927, B => n926, 
                           ZN => n929);
   U1260 : OAI211_X1 port map( C1 => n931, C2 => n1233, A => n930, B => n929, 
                           ZN => Y(17));
   U1261 : OAI22_X1 port map( A1 => n932, A2 => n965, B1 => n982, B2 => n1368, 
                           ZN => n933);
   U1262 : AOI211_X1 port map( C1 => n1252, C2 => n934, A => n1121, B => n933, 
                           ZN => n961);
   U1263 : NAND4_X1 port map( A1 => n938, A2 => n937, A3 => n936, A4 => n935, 
                           ZN => n1316);
   U1264 : INV_X1 port map( A => n1316, ZN => n1210);
   U1265 : INV_X1 port map( A => n939, ZN => n1068);
   U1266 : OAI22_X1 port map( A1 => n1210, A2 => n1061, B1 => n1068, B2 => 
                           n1233, ZN => n947);
   U1267 : INV_X1 port map( A => n940, ZN => n945);
   U1268 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_18, B1 => 
                           OP_A_12_port, B2 => n60, C1 => OP_A_11_port, C2 => 
                           n1027, ZN => n978);
   U1269 : XOR2_X1 port map( A => n978, B => intadd_1_SUM_12_port, Z => n941);
   U1270 : XNOR2_X1 port map( A => intadd_2_n1, B => n941, ZN => n942);
   U1271 : AOI22_X1 port map( A1 => n986, A2 => n942, B1 => n1242, B2 => n1207,
                           ZN => n944);
   U1272 : AOI22_X1 port map( A1 => n1348, A2 => OP2(18), B1 => n1347, B2 => 
                           OP1(18), ZN => n943);
   U1273 : OAI211_X1 port map( C1 => n945, C2 => n1111, A => n944, B => n943, 
                           ZN => n946);
   U1274 : AOI211_X1 port map( C1 => n948, C2 => n1245, A => n947, B => n946, 
                           ZN => n960);
   U1275 : NAND2_X1 port map( A1 => n951, A2 => n949, ZN => n956);
   U1276 : INV_X1 port map( A => n950, ZN => n955);
   U1277 : OAI21_X1 port map( B1 => n953, B2 => n952, A => n951, ZN => n954);
   U1278 : OAI21_X1 port map( B1 => n956, B2 => n955, A => n954, ZN => n981);
   U1279 : XNOR2_X1 port map( A => n958, B => n981, ZN => n957);
   U1280 : AOI22_X1 port map( A1 => n958, A2 => n1344, B1 => N279, B2 => n957, 
                           ZN => n959);
   U1281 : NAND3_X1 port map( A1 => n961, A2 => n960, A3 => n959, ZN => Y(18));
   U1282 : AOI22_X1 port map( A1 => n1348, A2 => OP2(19), B1 => n1347, B2 => 
                           OP1(19), ZN => n962);
   U1283 : OAI21_X1 port map( B1 => n963, B2 => n1111, A => n962, ZN => n968);
   U1284 : INV_X1 port map( A => n1252, ZN => n1181);
   U1285 : OAI22_X1 port map( A1 => n966, A2 => n965, B1 => n964, B2 => n1181, 
                           ZN => n967);
   U1286 : AOI211_X1 port map( C1 => n1367, C2 => n991, A => n968, B => n967, 
                           ZN => n990);
   U1287 : NAND4_X1 port map( A1 => n972, A2 => n971, A3 => n970, A4 => n969, 
                           ZN => n1351);
   U1288 : INV_X1 port map( A => n1233, ZN => n1122);
   U1289 : AOI22_X1 port map( A1 => n1228, A2 => n1351, B1 => n1122, B2 => n973
                           , ZN => n989);
   U1290 : OAI22_X1 port map( A1 => n975, A2 => n1369, B1 => n1372, B2 => n974,
                           ZN => n976);
   U1291 : AOI211_X1 port map( C1 => n1242, C2 => n1229, A => n1121, B => n976,
                           ZN => n988);
   U1292 : AND2_X1 port map( A1 => intadd_1_SUM_12_port, A2 => intadd_2_n1, ZN 
                           => n977);
   U1293 : OAI22_X1 port map( A1 => n978, A2 => n977, B1 => 
                           intadd_1_SUM_12_port, B2 => intadd_2_n1, ZN => n994)
                           ;
   U1294 : AOI222_X1 port map( A1 => n1083, A2 => C429_DATA4_19, B1 => 
                           OP_A_12_port, B2 => n1027, C1 => n60, C2 => 
                           OP_A_13_port, ZN => n997);
   U1295 : XNOR2_X1 port map( A => intadd_1_SUM_13_port, B => n997, ZN => n979)
                           ;
   U1296 : XNOR2_X1 port map( A => n994, B => n979, ZN => n985);
   U1297 : OAI21_X1 port map( B1 => n982, B2 => n981, A => n980, ZN => n992);
   U1298 : XOR2_X1 port map( A => n983, B => n992, Z => n984);
   U1299 : AOI22_X1 port map( A1 => n986, A2 => n985, B1 => n984, B2 => N279, 
                           ZN => n987);
   U1300 : NAND4_X1 port map( A1 => n990, A2 => n989, A3 => n988, A4 => n987, 
                           ZN => Y(19));
   U1301 : AOI22_X1 port map( A1 => n1242, A2 => n1268, B1 => n1122, B2 => 
                           n1119, ZN => n1017);
   U1302 : AOI22_X1 port map( A1 => OP_A_19_port, A2 => OP_B_19_port, B1 => 
                           n992, B2 => n991, ZN => n1047);
   U1303 : NOR2_X1 port map( A1 => n1047, A2 => n1018, ZN => n993);
   U1304 : AOI211_X1 port map( C1 => n1047, C2 => n1018, A => n1398, B => n993,
                           ZN => n1015);
   U1305 : INV_X1 port map( A => n994, ZN => n998);
   U1306 : INV_X1 port map( A => intadd_1_SUM_13_port, ZN => n995);
   U1307 : NAND2_X1 port map( A1 => n995, A2 => n994, ZN => n996);
   U1308 : AOI22_X1 port map( A1 => intadd_1_SUM_13_port, A2 => n998, B1 => 
                           n997, B2 => n996, ZN => n1026);
   U1309 : AOI222_X1 port map( A1 => n1414, A2 => C429_DATA4_20, B1 => n60, B2 
                           => OP_A_14_port, C1 => n1027, C2 => OP_A_13_port, ZN
                           => n1022);
   U1310 : INV_X1 port map( A => intadd_1_SUM_14_port, ZN => n1025);
   U1311 : XNOR2_X1 port map( A => n1022, B => n1025, ZN => n999);
   U1312 : XNOR2_X1 port map( A => n1026, B => n999, ZN => n1000);
   U1313 : NOR2_X1 port map( A1 => n1000, A2 => n1284, ZN => n1014);
   U1314 : AOI22_X1 port map( A1 => n1348, A2 => OP2(20), B1 => n1347, B2 => 
                           OP1(20), ZN => n1001);
   U1315 : OAI211_X1 port map( C1 => n1369, C2 => n1046, A => n1001, B => n1109
                           , ZN => n1013);
   U1316 : INV_X1 port map( A => n1244, ZN => n1211);
   U1317 : NAND4_X1 port map( A1 => n1005, A2 => n1004, A3 => n1003, A4 => 
                           n1002, ZN => n1269);
   U1318 : AOI22_X1 port map( A1 => n1228, A2 => n1269, B1 => n1230, B2 => 
                           n1006, ZN => n1010);
   U1319 : AOI22_X1 port map( A1 => n1252, A2 => n1008, B1 => n1367, B2 => 
                           n1007, ZN => n1009);
   U1320 : OAI211_X1 port map( C1 => n1211, C2 => n1011, A => n1010, B => n1009
                           , ZN => n1012);
   U1321 : NOR4_X1 port map( A1 => n1015, A2 => n1014, A3 => n1013, A4 => n1012
                           , ZN => n1016);
   U1322 : OAI211_X1 port map( C1 => n1018, C2 => n1372, A => n1017, B => n1016
                           , ZN => Y(20));
   U1323 : AOI21_X1 port map( B1 => n1047, B2 => n1046, A => n1049, ZN => n1019
                           );
   U1324 : XNOR2_X1 port map( A => n1020, B => n1019, ZN => n1045);
   U1325 : AOI22_X1 port map( A1 => n1021, A2 => n1245, B1 => n1020, B2 => 
                           n1344, ZN => n1044);
   U1326 : INV_X1 port map( A => n1026, ZN => n1023);
   U1327 : OAI21_X1 port map( B1 => intadd_1_SUM_14_port, B2 => n1023, A => 
                           n1022, ZN => n1024);
   U1328 : OAI21_X1 port map( B1 => n1026, B2 => n1025, A => n1024, ZN => n1076
                           );
   U1329 : INV_X1 port map( A => n1076, ZN => n1073);
   U1330 : CLKBUF_X1 port map( A => n1414, Z => n1083);
   U1331 : AOI222_X1 port map( A1 => OP_A_15_port, A2 => n60, B1 => n1083, B2 
                           => C429_DATA4_21, C1 => n1027, C2 => OP_A_14_port, 
                           ZN => n1075);
   U1332 : INV_X1 port map( A => intadd_1_SUM_15_port, ZN => n1072);
   U1333 : XNOR2_X1 port map( A => n1075, B => n1072, ZN => n1028);
   U1334 : XNOR2_X1 port map( A => n1073, B => n1028, ZN => n1032);
   U1335 : AOI22_X1 port map( A1 => n1348, A2 => OP2(21), B1 => n1330, B2 => 
                           OP1(21), ZN => n1031);
   U1336 : AOI22_X1 port map( A1 => n1244, A2 => n1029, B1 => n1242, B2 => 
                           n1285, ZN => n1030);
   U1337 : OAI211_X1 port map( C1 => n1032, C2 => n1284, A => n1031, B => n1030
                           , ZN => n1042);
   U1338 : NAND4_X1 port map( A1 => n1036, A2 => n1035, A3 => n1034, A4 => 
                           n1033, ZN => n1286);
   U1339 : AOI22_X1 port map( A1 => n1228, A2 => n1286, B1 => n1230, B2 => 
                           n1037, ZN => n1040);
   U1340 : AOI21_X1 port map( B1 => n1252, B2 => n1038, A => n1121, ZN => n1039
                           );
   U1341 : OAI211_X1 port map( C1 => n1050, C2 => n1368, A => n1040, B => n1039
                           , ZN => n1041);
   U1342 : AOI211_X1 port map( C1 => n1122, C2 => n1170, A => n1042, B => n1041
                           , ZN => n1043);
   U1343 : OAI211_X1 port map( C1 => n1398, C2 => n1045, A => n1044, B => n1043
                           , ZN => Y(21));
   U1344 : INV_X1 port map( A => n1125, ZN => n1055);
   U1345 : NAND2_X1 port map( A1 => n1048, A2 => n1046, ZN => n1053);
   U1346 : INV_X1 port map( A => n1047, ZN => n1052);
   U1347 : OAI21_X1 port map( B1 => n1050, B2 => n1049, A => n1048, ZN => n1051
                           );
   U1348 : OAI21_X1 port map( B1 => n1053, B2 => n1052, A => n1051, ZN => n1126
                           );
   U1349 : INV_X1 port map( A => n1126, ZN => n1054);
   U1350 : AOI221_X1 port map( B1 => n1055, B2 => n1054, C1 => n1125, C2 => 
                           n1126, A => n1398, ZN => n1071);
   U1351 : NOR2_X1 port map( A1 => OP_A_22_port, A2 => OP_B_22_port, ZN => 
                           n1104);
   U1352 : OAI22_X1 port map( A1 => n1104, A2 => n1368, B1 => n1124, B2 => 
                           n1369, ZN => n1070);
   U1353 : AOI22_X1 port map( A1 => n1348, A2 => OP2(22), B1 => n1330, B2 => 
                           OP1(22), ZN => n1067);
   U1354 : NAND4_X1 port map( A1 => n1059, A2 => n1058, A3 => n1057, A4 => 
                           n1056, ZN => n1317);
   U1355 : INV_X1 port map( A => n1317, ZN => n1184);
   U1356 : INV_X1 port map( A => n1207, ZN => n1060);
   U1357 : OAI22_X1 port map( A1 => n1184, A2 => n1061, B1 => n1060, B2 => 
                           n1233, ZN => n1064);
   U1358 : INV_X1 port map( A => n1242, ZN => n1183);
   U1359 : OAI22_X1 port map( A1 => n1210, A2 => n1183, B1 => n1062, B2 => 
                           n1211, ZN => n1063);
   U1360 : AOI211_X1 port map( C1 => n1252, C2 => n1065, A => n1064, B => n1063
                           , ZN => n1066);
   U1361 : OAI211_X1 port map( C1 => n1068, C2 => n1111, A => n1067, B => n1066
                           , ZN => n1069);
   U1362 : NOR4_X1 port map( A1 => n1121, A2 => n1071, A3 => n1070, A4 => n1069
                           , ZN => n1088);
   U1363 : NAND2_X1 port map( A1 => n1073, A2 => n1072, ZN => n1074);
   U1364 : AOI22_X1 port map( A1 => intadd_1_SUM_15_port, A2 => n1076, B1 => 
                           n1075, B2 => n1074, ZN => n1091);
   U1365 : OAI21_X1 port map( B1 => OP_A_15_port, B2 => n1078, A => n1077, ZN 
                           => n1079);
   U1366 : INV_X1 port map( A => n1079, ZN => n1092);
   U1367 : XNOR2_X1 port map( A => DP_OP_446J3_125_4819_n12, B => n1092, ZN => 
                           n1082);
   U1368 : AOI21_X1 port map( B1 => n1083, B2 => n1082, A => n1380, ZN => n1084
                           );
   U1369 : INV_X1 port map( A => n1084, ZN => n1090);
   U1370 : XNOR2_X1 port map( A => n1091, B => n1090, ZN => n1086);
   U1371 : AOI21_X1 port map( B1 => intadd_1_SUM_16_port, B2 => n1086, A => 
                           n1284, ZN => n1085);
   U1372 : OAI21_X1 port map( B1 => intadd_1_SUM_16_port, B2 => n1086, A => 
                           n1085, ZN => n1087);
   U1373 : OAI211_X1 port map( C1 => n1372, C2 => n1125, A => n1088, B => n1087
                           , ZN => Y(22));
   U1374 : INV_X1 port map( A => intadd_1_SUM_16_port, ZN => n1089);
   U1375 : FA_X1 port map( A => n1091, B => n1090, CI => n1089, CO => n1093, S 
                           => n_1170);
   U1376 : NOR3_X1 port map( A1 => n1093, A2 => n65, A3 => n1380, ZN => n1143);
   U1377 : INV_X1 port map( A => n1143, ZN => n1094);
   U1378 : OAI21_X1 port map( B1 => n1380, B2 => n65, A => n1093, ZN => n1144);
   U1379 : NAND2_X1 port map( A1 => n1094, A2 => n1144, ZN => n1095);
   U1380 : XNOR2_X1 port map( A => intadd_1_SUM_17_port, B => n1095, ZN => 
                           n1118);
   U1381 : NAND4_X1 port map( A1 => n1099, A2 => n1098, A3 => n1097, A4 => 
                           n1096, ZN => n1349);
   U1382 : AOI22_X1 port map( A1 => n1228, A2 => n1349, B1 => n1122, B2 => 
                           n1229, ZN => n1102);
   U1383 : AOI22_X1 port map( A1 => n1244, A2 => n1100, B1 => n1242, B2 => 
                           n1351, ZN => n1101);
   U1384 : OAI211_X1 port map( C1 => n1123, C2 => n1369, A => n1102, B => n1101
                           , ZN => n1103);
   U1385 : AOI21_X1 port map( B1 => n1344, B2 => n1106, A => n1103, ZN => n1117
                           );
   U1386 : OAI21_X1 port map( B1 => n1104, B2 => n1126, A => n1124, ZN => n1105
                           );
   U1387 : XOR2_X1 port map( A => n1106, B => n1105, Z => n1115);
   U1388 : OAI22_X1 port map( A1 => n1108, A2 => n1368, B1 => n1107, B2 => 
                           n1181, ZN => n1114);
   U1389 : AOI22_X1 port map( A1 => n1348, A2 => OP2(23), B1 => n1330, B2 => 
                           OP1(23), ZN => n1110);
   U1390 : OAI211_X1 port map( C1 => n1112, C2 => n1111, A => n1110, B => n1109
                           , ZN => n1113);
   U1391 : AOI211_X1 port map( C1 => n1115, C2 => N279, A => n1114, B => n1113,
                           ZN => n1116);
   U1392 : OAI211_X1 port map( C1 => n1284, C2 => n1118, A => n1117, B => n1116
                           , ZN => Y(23));
   U1393 : AOI22_X1 port map( A1 => n1242, A2 => n1269, B1 => n1230, B2 => 
                           n1119, ZN => n1152);
   U1394 : OAI22_X1 port map( A1 => n1193, A2 => n1369, B1 => n1129, B2 => 
                           n1372, ZN => n1120);
   U1395 : AOI211_X1 port map( C1 => n1122, C2 => n1268, A => n1121, B => n1120
                           , ZN => n1151);
   U1396 : OAI211_X1 port map( C1 => n1126, C2 => n1125, A => n1124, B => n1123
                           , ZN => n1127);
   U1397 : OAI21_X1 port map( B1 => OP_A_23_port, B2 => OP_B_23_port, A => 
                           n1127, ZN => n1192);
   U1398 : NOR2_X1 port map( A1 => n1192, A2 => n1129, ZN => n1128);
   U1399 : AOI211_X1 port map( C1 => n1192, C2 => n1129, A => n1398, B => n1128
                           , ZN => n1141);
   U1400 : NAND4_X1 port map( A1 => n1133, A2 => n1132, A3 => n1131, A4 => 
                           n1130, ZN => n1274);
   U1401 : AOI22_X1 port map( A1 => n1330, A2 => OP1(24), B1 => n1228, B2 => 
                           n1274, ZN => n1137);
   U1402 : AOI22_X1 port map( A1 => n1252, A2 => n1135, B1 => n1244, B2 => 
                           n1134, ZN => n1136);
   U1403 : OAI211_X1 port map( C1 => n1139, C2 => n1138, A => n1137, B => n1136
                           , ZN => n1140);
   U1404 : AOI211_X1 port map( C1 => n1367, C2 => n1142, A => n1141, B => n1140
                           , ZN => n1150);
   U1405 : AOI21_X1 port map( B1 => intadd_1_SUM_17_port, B2 => n1144, A => 
                           n1143, ZN => n1145);
   U1406 : NOR3_X1 port map( A1 => n1145, A2 => n65, A3 => n1380, ZN => n1153);
   U1407 : INV_X1 port map( A => n1153, ZN => n1146);
   U1408 : OAI21_X1 port map( B1 => n1380, B2 => n65, A => n1145, ZN => n1154);
   U1409 : NAND2_X1 port map( A1 => n1146, A2 => n1154, ZN => n1148);
   U1410 : AOI21_X1 port map( B1 => intadd_1_SUM_18_port, B2 => n1148, A => 
                           n1284, ZN => n1147);
   U1411 : OAI21_X1 port map( B1 => intadd_1_SUM_18_port, B2 => n1148, A => 
                           n1147, ZN => n1149);
   U1412 : NAND4_X1 port map( A1 => n1152, A2 => n1151, A3 => n1150, A4 => 
                           n1149, ZN => Y(24));
   U1413 : AOI21_X1 port map( B1 => intadd_1_SUM_18_port, B2 => n1154, A => 
                           n1153, ZN => n1155);
   U1414 : NOR3_X1 port map( A1 => n1155, A2 => n65, A3 => n1380, ZN => n1186);
   U1415 : INV_X1 port map( A => n1186, ZN => n1156);
   U1416 : OAI21_X1 port map( B1 => n1380, B2 => n65, A => n1155, ZN => n1187);
   U1417 : NAND2_X1 port map( A1 => n1156, A2 => n1187, ZN => n1157);
   U1418 : XNOR2_X1 port map( A => intadd_1_SUM_19_port, B => n1157, ZN => 
                           n1180);
   U1419 : AOI211_X1 port map( C1 => n1160, C2 => n1363, A => n1159, B => n1158
                           , ZN => n1236);
   U1420 : AOI22_X1 port map( A1 => n1244, A2 => n1161, B1 => n1242, B2 => 
                           n1286, ZN => n1162);
   U1421 : OAI21_X1 port map( B1 => n1194, B2 => n1369, A => n1162, ZN => n1163
                           );
   U1422 : AOI211_X1 port map( C1 => n1165, C2 => n1344, A => n1236, B => n1163
                           , ZN => n1179);
   U1423 : AOI21_X1 port map( B1 => n1192, B2 => n1193, A => n1195, ZN => n1164
                           );
   U1424 : XOR2_X1 port map( A => n1165, B => n1164, Z => n1177);
   U1425 : INV_X1 port map( A => n1285, ZN => n1173);
   U1426 : NAND4_X1 port map( A1 => n1169, A2 => n1168, A3 => n1167, A4 => 
                           n1166, ZN => n1291);
   U1427 : AOI22_X1 port map( A1 => n1230, A2 => n1170, B1 => n1228, B2 => 
                           n1291, ZN => n1172);
   U1428 : AOI22_X1 port map( A1 => n1348, A2 => OP2(25), B1 => n1330, B2 => 
                           OP1(25), ZN => n1171);
   U1429 : OAI211_X1 port map( C1 => n1173, C2 => n1233, A => n1172, B => n1171
                           , ZN => n1176);
   U1430 : OAI22_X1 port map( A1 => n1196, A2 => n1368, B1 => n1174, B2 => 
                           n1181, ZN => n1175);
   U1431 : AOI211_X1 port map( C1 => n1177, C2 => N279, A => n1176, B => n1175,
                           ZN => n1178);
   U1432 : OAI211_X1 port map( C1 => n1284, C2 => n1180, A => n1179, B => n1178
                           , ZN => Y(25));
   U1433 : INV_X1 port map( A => n1200, ZN => n1202);
   U1434 : OAI22_X1 port map( A1 => n1184, A2 => n1183, B1 => n1182, B2 => 
                           n1181, ZN => n1185);
   U1435 : AOI211_X1 port map( C1 => n1202, C2 => n1344, A => n1236, B => n1185
                           , ZN => n1218);
   U1436 : AOI21_X1 port map( B1 => intadd_1_SUM_19_port, B2 => n1187, A => 
                           n1186, ZN => n1188);
   U1437 : NOR3_X1 port map( A1 => n1188, A2 => n65, A3 => n1380, ZN => n1219);
   U1438 : INV_X1 port map( A => n1219, ZN => n1189);
   U1439 : OAI21_X1 port map( B1 => n1380, B2 => n65, A => n1188, ZN => n1220);
   U1440 : NAND2_X1 port map( A1 => n1189, A2 => n1220, ZN => n1191);
   U1441 : NOR2_X1 port map( A1 => intadd_1_SUM_20_port, A2 => n1191, ZN => 
                           n1190);
   U1442 : AOI211_X1 port map( C1 => intadd_1_SUM_20_port, C2 => n1191, A => 
                           n1284, B => n1190, ZN => n1216);
   U1443 : INV_X1 port map( A => n1192, ZN => n1199);
   U1444 : NAND2_X1 port map( A1 => n1194, A2 => n1193, ZN => n1198);
   U1445 : OAI21_X1 port map( B1 => n1196, B2 => n1195, A => n1194, ZN => n1197
                           );
   U1446 : OAI21_X1 port map( B1 => n1199, B2 => n1198, A => n1197, ZN => n1238
                           );
   U1447 : INV_X1 port map( A => n1238, ZN => n1201);
   U1448 : AOI221_X1 port map( B1 => n1202, B2 => n1201, C1 => n1200, C2 => 
                           n1238, A => n1398, ZN => n1215);
   U1449 : NAND4_X1 port map( A1 => n1206, A2 => n1205, A3 => n1204, A4 => 
                           n1203, ZN => n1322);
   U1450 : AOI22_X1 port map( A1 => n1230, A2 => n1207, B1 => n1228, B2 => 
                           n1322, ZN => n1209);
   U1451 : AOI22_X1 port map( A1 => n1348, A2 => OP2(26), B1 => n1330, B2 => 
                           OP1(26), ZN => n1208);
   U1452 : OAI211_X1 port map( C1 => n1210, C2 => n1233, A => n1209, B => n1208
                           , ZN => n1214);
   U1453 : NOR2_X1 port map( A1 => OP_A_26_port, A2 => OP_B_26_port, ZN => 
                           n1239);
   U1454 : OAI22_X1 port map( A1 => n1239, A2 => n1368, B1 => n1212, B2 => 
                           n1211, ZN => n1213);
   U1455 : NOR4_X1 port map( A1 => n1216, A2 => n1215, A3 => n1214, A4 => n1213
                           , ZN => n1217);
   U1456 : OAI211_X1 port map( C1 => n1237, C2 => n1369, A => n1218, B => n1217
                           , ZN => Y(26));
   U1457 : AOI21_X1 port map( B1 => intadd_1_SUM_20_port, B2 => n1220, A => 
                           n1219, ZN => n1221);
   U1458 : NOR3_X1 port map( A1 => n1221, A2 => n65, A3 => n1380, ZN => n1256);
   U1459 : INV_X1 port map( A => n1256, ZN => n1222);
   U1460 : OAI21_X1 port map( B1 => n1380, B2 => n65, A => n1221, ZN => n1257);
   U1461 : NAND2_X1 port map( A1 => n1222, A2 => n1257, ZN => n1223);
   U1462 : XNOR2_X1 port map( A => intadd_1_SUM_21_port, B => n1223, ZN => 
                           n1255);
   U1463 : INV_X1 port map( A => n1351, ZN => n1234);
   U1464 : NAND4_X1 port map( A1 => n1227, A2 => n1226, A3 => n1225, A4 => 
                           n1224, ZN => n1357);
   U1465 : AOI22_X1 port map( A1 => n1230, A2 => n1229, B1 => n1228, B2 => 
                           n1357, ZN => n1232);
   U1466 : AOI22_X1 port map( A1 => n1348, A2 => OP2(27), B1 => n1330, B2 => 
                           OP1(27), ZN => n1231);
   U1467 : OAI211_X1 port map( C1 => n1234, C2 => n1233, A => n1232, B => n1231
                           , ZN => n1235);
   U1468 : AOI211_X1 port map( C1 => n1344, C2 => n1241, A => n1236, B => n1235
                           , ZN => n1254);
   U1469 : OAI21_X1 port map( B1 => n1239, B2 => n1238, A => n1237, ZN => n1266
                           );
   U1470 : OAI21_X1 port map( B1 => n1241, B2 => n1266, A => N279, ZN => n1240)
                           ;
   U1471 : AOI21_X1 port map( B1 => n1241, B2 => n1266, A => n1240, ZN => n1250
                           );
   U1472 : AOI22_X1 port map( A1 => n1244, A2 => n1243, B1 => n1242, B2 => 
                           n1349, ZN => n1247);
   U1473 : OAI221_X1 port map( B1 => n1367, B2 => n1245, C1 => n1367, C2 => 
                           OP_A_27_port, A => OP_B_27_port, ZN => n1246);
   U1474 : OAI211_X1 port map( C1 => n1368, C2 => n1248, A => n1247, B => n1246
                           , ZN => n1249);
   U1475 : AOI211_X1 port map( C1 => n1252, C2 => n1251, A => n1250, B => n1249
                           , ZN => n1253);
   U1476 : OAI211_X1 port map( C1 => n1284, C2 => n1255, A => n1254, B => n1253
                           , ZN => Y(27));
   U1477 : AOI21_X1 port map( B1 => intadd_1_SUM_21_port, B2 => n1257, A => 
                           n1256, ZN => n1258);
   U1478 : NOR3_X1 port map( A1 => n1258, A2 => n65, A3 => n1380, ZN => n1303);
   U1479 : INV_X1 port map( A => n1303, ZN => n1259);
   U1480 : OAI21_X1 port map( B1 => n1380, B2 => n65, A => n1258, ZN => n1304);
   U1481 : NAND2_X1 port map( A1 => n1259, A2 => n1304, ZN => n1260);
   U1482 : XNOR2_X1 port map( A => intadd_1_SUM_22_port, B => n1260, ZN => 
                           n1283);
   U1483 : AOI22_X1 port map( A1 => n1348, A2 => OP2(28), B1 => n1330, B2 => 
                           OP1(28), ZN => n1262);
   U1484 : NAND3_X1 port map( A1 => OP_SHIFT, A2 => N284, A3 => n1261, ZN => 
                           n1402);
   U1485 : OAI211_X1 port map( C1 => n1299, C2 => n1368, A => n1262, B => n1402
                           , ZN => n1264);
   U1486 : OAI22_X1 port map( A1 => n1301, A2 => n1369, B1 => n1372, B2 => 
                           n1267, ZN => n1263);
   U1487 : AOI211_X1 port map( C1 => n1329, C2 => n1265, A => n1264, B => n1263
                           , ZN => n1282);
   U1488 : AOI222_X1 port map( A1 => OP_A_27_port, A2 => OP_B_27_port, B1 => 
                           OP_A_27_port, B2 => n1266, C1 => OP_B_27_port, C2 =>
                           n1266, ZN => n1300);
   U1489 : XOR2_X1 port map( A => n1267, B => n1300, Z => n1280);
   U1490 : AOI22_X1 port map( A1 => n1350, A2 => n1269, B1 => n1352, B2 => 
                           n1268, ZN => n1277);
   U1491 : NAND2_X1 port map( A1 => OP_A_28_port, A2 => n56, ZN => n1273);
   U1492 : NAND4_X1 port map( A1 => n1273, A2 => n1272, A3 => n1271, A4 => 
                           n1270, ZN => n1275);
   U1493 : AOI22_X1 port map( A1 => n1360, A2 => n1275, B1 => n1358, B2 => 
                           n1274, ZN => n1276);
   U1494 : OAI211_X1 port map( C1 => n1278, C2 => n1363, A => n1277, B => n1276
                           , ZN => n1279);
   U1495 : AOI22_X1 port map( A1 => n1280, A2 => N279, B1 => n1366, B2 => n1279
                           , ZN => n1281);
   U1496 : OAI211_X1 port map( C1 => n1284, C2 => n1283, A => n1282, B => n1281
                           , ZN => Y(28));
   U1497 : AOI22_X1 port map( A1 => n1348, A2 => OP2(29), B1 => n1330, B2 => 
                           OP1(29), ZN => n1315);
   U1498 : AOI22_X1 port map( A1 => n1350, A2 => n1286, B1 => n1352, B2 => 
                           n1285, ZN => n1294);
   U1499 : NAND4_X1 port map( A1 => n1290, A2 => n1289, A3 => n1288, A4 => 
                           n1287, ZN => n1292);
   U1500 : AOI22_X1 port map( A1 => n1360, A2 => n1292, B1 => n1358, B2 => 
                           n1291, ZN => n1293);
   U1501 : OAI211_X1 port map( C1 => n1295, C2 => n1363, A => n1294, B => n1293
                           , ZN => n1296);
   U1502 : AOI22_X1 port map( A1 => OP_A_29_port, A2 => n1367, B1 => n1366, B2 
                           => n1296, ZN => n1314);
   U1503 : OAI21_X1 port map( B1 => n1297, B2 => n1369, A => n1368, ZN => n1312
                           );
   U1504 : OAI22_X1 port map( A1 => n1302, A2 => n1372, B1 => n1298, B2 => 
                           n1373, ZN => n1311);
   U1505 : AOI21_X1 port map( B1 => n1301, B2 => n1300, A => n1299, ZN => n1332
                           );
   U1506 : XOR2_X1 port map( A => n1332, B => n1302, Z => n1309);
   U1507 : AOI21_X1 port map( B1 => intadd_1_SUM_22_port, B2 => n1304, A => 
                           n1303, ZN => n1305);
   U1508 : NOR3_X1 port map( A1 => n1305, A2 => n65, A3 => n1380, ZN => n1334);
   U1509 : INV_X1 port map( A => n1334, ZN => n1306);
   U1510 : OAI21_X1 port map( B1 => n1380, B2 => n65, A => n1305, ZN => n1335);
   U1511 : NAND2_X1 port map( A1 => n1306, A2 => n1335, ZN => n1307);
   U1512 : XNOR2_X1 port map( A => intadd_1_SUM_23_port, B => n1307, ZN => 
                           n1308);
   U1513 : OAI22_X1 port map( A1 => n1398, A2 => n1309, B1 => n1396, B2 => 
                           n1308, ZN => n1310);
   U1514 : AOI211_X1 port map( C1 => OP_B_29_port, C2 => n1312, A => n1311, B 
                           => n1310, ZN => n1313);
   U1515 : NAND4_X1 port map( A1 => n1315, A2 => n1314, A3 => n1313, A4 => 
                           n1402, ZN => Y(29));
   U1516 : AOI22_X1 port map( A1 => n1350, A2 => n1317, B1 => n1352, B2 => 
                           n1316, ZN => n1325);
   U1517 : NAND2_X1 port map( A1 => OP_A_30_port, A2 => n56, ZN => n1321);
   U1518 : NAND4_X1 port map( A1 => n1321, A2 => n1320, A3 => n1319, A4 => 
                           n1318, ZN => n1323);
   U1519 : AOI22_X1 port map( A1 => n1360, A2 => n1323, B1 => n1358, B2 => 
                           n1322, ZN => n1324);
   U1520 : OAI211_X1 port map( C1 => n1326, C2 => n1363, A => n1325, B => n1324
                           , ZN => n1327);
   U1521 : AOI22_X1 port map( A1 => n1329, A2 => n1328, B1 => n1366, B2 => 
                           n1327, ZN => n1346);
   U1522 : AOI22_X1 port map( A1 => n1348, A2 => OP2(30), B1 => n1330, B2 => 
                           OP1(30), ZN => n1331);
   U1523 : OAI211_X1 port map( C1 => n1375, C2 => n1368, A => n1331, B => n1402
                           , ZN => n1342);
   U1524 : AOI222_X1 port map( A1 => OP_B_29_port, A2 => OP_A_29_port, B1 => 
                           OP_B_29_port, B2 => n1332, C1 => OP_A_29_port, C2 =>
                           n1332, ZN => n1376);
   U1525 : XNOR2_X1 port map( A => n1376, B => n1333, ZN => n1340);
   U1526 : AOI21_X1 port map( B1 => intadd_1_SUM_23_port, B2 => n1335, A => 
                           n1334, ZN => n1336);
   U1527 : NOR3_X1 port map( A1 => n1336, A2 => n65, A3 => n1380, ZN => n1386);
   U1528 : INV_X1 port map( A => n1386, ZN => n1337);
   U1529 : OAI21_X1 port map( B1 => n1380, B2 => n65, A => n1336, ZN => n1387);
   U1530 : NAND2_X1 port map( A1 => n1337, A2 => n1387, ZN => n1338);
   U1531 : XNOR2_X1 port map( A => intadd_1_SUM_24_port, B => n1338, ZN => 
                           n1339);
   U1532 : OAI22_X1 port map( A1 => n1398, A2 => n1340, B1 => n1396, B2 => 
                           n1339, ZN => n1341);
   U1533 : AOI211_X1 port map( C1 => n1344, C2 => n1343, A => n1342, B => n1341
                           , ZN => n1345);
   U1534 : OAI211_X1 port map( C1 => n1377, C2 => n1369, A => n1346, B => n1345
                           , ZN => Y(30));
   U1535 : AOI22_X1 port map( A1 => n1348, A2 => OP2(31), B1 => OP1(31), B2 => 
                           n1347, ZN => n1405);
   U1536 : AOI22_X1 port map( A1 => n1352, A2 => n1351, B1 => n1350, B2 => 
                           n1349, ZN => n1362);
   U1537 : NAND2_X1 port map( A1 => OP_A_31_port, A2 => n56, ZN => n1356);
   U1538 : NAND4_X1 port map( A1 => n1356, A2 => n1355, A3 => n1354, A4 => 
                           n1353, ZN => n1359);
   U1539 : AOI22_X1 port map( A1 => n1360, A2 => n1359, B1 => n1358, B2 => 
                           n1357, ZN => n1361);
   U1540 : OAI211_X1 port map( C1 => n1364, C2 => n1363, A => n1362, B => n1361
                           , ZN => n1365);
   U1541 : AOI22_X1 port map( A1 => OP_A_31_port, A2 => n1367, B1 => n1366, B2 
                           => n1365, ZN => n1404);
   U1542 : OAI21_X1 port map( B1 => n1370, B2 => n1369, A => n1368, ZN => n1401
                           );
   U1543 : INV_X1 port map( A => n1371, ZN => n1378);
   U1544 : OAI22_X1 port map( A1 => n1374, A2 => n1373, B1 => n1378, B2 => 
                           n1372, ZN => n1400);
   U1545 : AOI21_X1 port map( B1 => n1377, B2 => n1376, A => n1375, ZN => n1379
                           );
   U1546 : XOR2_X1 port map( A => n1379, B => n1378, Z => n1397);
   U1547 : NOR2_X1 port map( A1 => n65, A2 => n1380, ZN => n1385);
   U1548 : INV_X1 port map( A => n1381, ZN => n1382);
   U1549 : AOI21_X1 port map( B1 => n1383, B2 => n1382, A => n1385, ZN => n1384
                           );
   U1550 : AOI21_X1 port map( B1 => n1385, B2 => intadd_1_B_18_port, A => n1384
                           , ZN => n1389);
   U1551 : AOI21_X1 port map( B1 => intadd_1_SUM_24_port, B2 => n1387, A => 
                           n1386, ZN => n1388);
   U1552 : XOR2_X1 port map( A => n1389, B => n1388, Z => n1390);
   U1553 : MUX2_X1 port map( A => n61, B => n58, S => n1390, Z => n1394);
   U1554 : INV_X1 port map( A => intadd_0_A_16_port, ZN => n1391);
   U1555 : MUX2_X1 port map( A => intadd_0_A_16_port, B => n1391, S => 
                           intadd_0_n1, Z => n1392);
   U1556 : XOR2_X1 port map( A => intadd_1_n1, B => n1392, Z => n1393);
   U1557 : XNOR2_X1 port map( A => n1394, B => n1393, ZN => n1395);
   U1558 : OAI22_X1 port map( A1 => n1398, A2 => n1397, B1 => n1396, B2 => 
                           n1395, ZN => n1399);
   U1559 : AOI211_X1 port map( C1 => OP_B_31_port, C2 => n1401, A => n1400, B 
                           => n1399, ZN => n1403);
   U1560 : NAND4_X1 port map( A1 => n1405, A2 => n1404, A3 => n1403, A4 => 
                           n1402, ZN => Y(31));
   U1561 : OAI22_X1 port map( A1 => OPC(6), A2 => n1407, B1 => n1406, B2 => 
                           n1411, ZN => N282);
   U1562 : OAI22_X1 port map( A1 => n1411, A2 => n1410, B1 => n1409, B2 => 
                           n1408, ZN => N283);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( CLK, RST : in std_logic);

end DLX;

architecture SYN_DLX_RTL of DLX is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component RF_N32_NA5
      port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
            ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component ALU_N32_NB8
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
            std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);
            Z : out std_logic);
   end component;
   
   component DLX_DRAM_N256_NW32
      port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector 
            (31 downto 0);  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component DLX_IRAM_RAM_DEPTH256_I_SIZE32
      port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  
            DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, 
      IR_26_port, IR_10_port, IR_9_port, IR_8_port, IR_7_port, IR_6_port, 
      IR_5_port, IR_4_port, IR_3_port, IR_2_port, IR_1_port, IR_0_port, 
      ALU_OPCODE_i_0_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_4_port, ALU_OPCODE_i_5_port, 
      ALU_OPCODE_i_6_port, IR_BUS_31_port, IR_BUS_30_port, IR_BUS_29_port, 
      IR_BUS_28_port, IR_BUS_27_port, IR_BUS_26_port, IR_BUS_25_port, 
      IR_BUS_24_port, IR_BUS_23_port, IR_BUS_22_port, IR_BUS_21_port, 
      IR_BUS_20_port, IR_BUS_19_port, IR_BUS_18_port, IR_BUS_17_port, 
      IR_BUS_16_port, IR_BUS_15_port, IR_BUS_14_port, IR_BUS_13_port, 
      IR_BUS_12_port, IR_BUS_11_port, IR_BUS_10_port, IR_BUS_9_port, 
      IR_BUS_8_port, IR_BUS_7_port, IR_BUS_6_port, IR_BUS_5_port, IR_BUS_4_port
      , IR_BUS_3_port, IR_BUS_2_port, IR_BUS_1_port, IR_BUS_0_port, 
      DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, DATA_OUT_28_port, 
      DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, DATA_OUT_24_port, 
      DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, 
      DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, 
      DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, 
      DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, 
      DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, 
      DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port, 
      DATA_ADDR_31_port, DATA_ADDR_30_port, DATA_ADDR_29_port, 
      DATA_ADDR_28_port, DATA_ADDR_27_port, DATA_ADDR_26_port, 
      DATA_ADDR_25_port, DATA_ADDR_24_port, DATA_ADDR_23_port, 
      DATA_ADDR_22_port, DATA_ADDR_21_port, DATA_ADDR_20_port, 
      DATA_ADDR_19_port, DATA_ADDR_18_port, DATA_ADDR_17_port, 
      DATA_ADDR_16_port, DATA_ADDR_15_port, DATA_ADDR_14_port, 
      DATA_ADDR_13_port, DATA_ADDR_12_port, DATA_ADDR_11_port, 
      DATA_ADDR_10_port, DATA_ADDR_9_port, DATA_ADDR_8_port, DATA_ADDR_7_port, 
      DATA_ADDR_6_port, DATA_ADDR_5_port, DATA_ADDR_4_port, DATA_ADDR_3_port, 
      DATA_ADDR_2_port, DATA_ADDR_1_port, DATA_ADDR_0_port, DATA_IN_31_port, 
      DATA_IN_30_port, DATA_IN_29_port, DATA_IN_28_port, DATA_IN_27_port, 
      DATA_IN_26_port, DATA_IN_25_port, DATA_IN_24_port, DATA_IN_23_port, 
      DATA_IN_22_port, DATA_IN_21_port, DATA_IN_20_port, DATA_IN_19_port, 
      DATA_IN_18_port, DATA_IN_17_port, DATA_IN_16_port, DATA_IN_15_port, 
      DATA_IN_14_port, DATA_IN_13_port, DATA_IN_12_port, DATA_IN_11_port, 
      DATA_IN_10_port, DATA_IN_9_port, DATA_IN_8_port, DATA_IN_7_port, 
      DATA_IN_6_port, DATA_IN_5_port, DATA_IN_4_port, DATA_IN_3_port, 
      DATA_IN_2_port, DATA_IN_1_port, DATA_IN_0_port, CU_I_aluOpcode2_0_port, 
      CU_I_aluOpcode2_1_port, CU_I_aluOpcode2_2_port, CU_I_aluOpcode2_3_port, 
      CU_I_aluOpcode2_4_port, CU_I_aluOpcode2_5_port, CU_I_aluOpcode2_6_port, 
      CU_I_aluOpcode1_0_port, CU_I_aluOpcode1_1_port, CU_I_aluOpcode1_2_port, 
      CU_I_aluOpcode1_3_port, CU_I_aluOpcode1_4_port, CU_I_aluOpcode1_5_port, 
      CU_I_aluOpcode1_6_port, DATAPATH_I_ALU_OUTPUT_0_port, 
      DATAPATH_I_ALU_OUTPUT_1_port, DATAPATH_I_ALU_OUTPUT_2_port, 
      DATAPATH_I_ALU_OUTPUT_3_port, DATAPATH_I_ALU_OUTPUT_4_port, 
      DATAPATH_I_ALU_OUTPUT_5_port, DATAPATH_I_ALU_OUTPUT_6_port, 
      DATAPATH_I_ALU_OUTPUT_7_port, DATAPATH_I_ALU_OUTPUT_8_port, 
      DATAPATH_I_ALU_OUTPUT_9_port, DATAPATH_I_ALU_OUTPUT_10_port, 
      DATAPATH_I_ALU_OUTPUT_11_port, DATAPATH_I_ALU_OUTPUT_12_port, 
      DATAPATH_I_ALU_OUTPUT_13_port, DATAPATH_I_ALU_OUTPUT_14_port, 
      DATAPATH_I_ALU_OUTPUT_15_port, DATAPATH_I_ALU_OUTPUT_16_port, 
      DATAPATH_I_ALU_OUTPUT_17_port, DATAPATH_I_ALU_OUTPUT_18_port, 
      DATAPATH_I_ALU_OUTPUT_19_port, DATAPATH_I_ALU_OUTPUT_20_port, 
      DATAPATH_I_ALU_OUTPUT_21_port, DATAPATH_I_ALU_OUTPUT_22_port, 
      DATAPATH_I_ALU_OUTPUT_23_port, DATAPATH_I_ALU_OUTPUT_24_port, 
      DATAPATH_I_ALU_OUTPUT_25_port, DATAPATH_I_ALU_OUTPUT_26_port, 
      DATAPATH_I_ALU_OUTPUT_27_port, DATAPATH_I_ALU_OUTPUT_28_port, 
      DATAPATH_I_ALU_OUTPUT_29_port, DATAPATH_I_ALU_OUTPUT_30_port, 
      DATAPATH_I_ALU_OUTPUT_31_port, DATAPATH_I_RF_OUT2_0_port, 
      DATAPATH_I_RF_OUT2_1_port, DATAPATH_I_RF_OUT2_2_port, 
      DATAPATH_I_RF_OUT2_3_port, DATAPATH_I_RF_OUT2_4_port, 
      DATAPATH_I_RF_OUT2_5_port, DATAPATH_I_RF_OUT2_6_port, 
      DATAPATH_I_RF_OUT2_7_port, DATAPATH_I_RF_OUT2_8_port, 
      DATAPATH_I_RF_OUT2_9_port, DATAPATH_I_RF_OUT2_10_port, 
      DATAPATH_I_RF_OUT2_11_port, DATAPATH_I_RF_OUT2_12_port, 
      DATAPATH_I_RF_OUT2_13_port, DATAPATH_I_RF_OUT2_14_port, 
      DATAPATH_I_RF_OUT2_15_port, DATAPATH_I_RF_OUT2_16_port, 
      DATAPATH_I_RF_OUT2_17_port, DATAPATH_I_RF_OUT2_18_port, 
      DATAPATH_I_RF_OUT2_19_port, DATAPATH_I_RF_OUT2_20_port, 
      DATAPATH_I_RF_OUT2_21_port, DATAPATH_I_RF_OUT2_22_port, 
      DATAPATH_I_RF_OUT2_23_port, DATAPATH_I_RF_OUT2_24_port, 
      DATAPATH_I_RF_OUT2_25_port, DATAPATH_I_RF_OUT2_26_port, 
      DATAPATH_I_RF_OUT2_27_port, DATAPATH_I_RF_OUT2_28_port, 
      DATAPATH_I_RF_OUT2_29_port, DATAPATH_I_RF_OUT2_30_port, 
      DATAPATH_I_RF_OUT2_31_port, DATAPATH_I_RF_OUT1_0_port, 
      DATAPATH_I_RF_OUT1_1_port, DATAPATH_I_RF_OUT1_2_port, 
      DATAPATH_I_RF_OUT1_3_port, DATAPATH_I_RF_OUT1_4_port, 
      DATAPATH_I_RF_OUT1_5_port, DATAPATH_I_RF_OUT1_6_port, 
      DATAPATH_I_RF_OUT1_7_port, DATAPATH_I_RF_OUT1_8_port, 
      DATAPATH_I_RF_OUT1_9_port, DATAPATH_I_RF_OUT1_10_port, 
      DATAPATH_I_RF_OUT1_11_port, DATAPATH_I_RF_OUT1_12_port, 
      DATAPATH_I_RF_OUT1_13_port, DATAPATH_I_RF_OUT1_14_port, 
      DATAPATH_I_RF_OUT1_15_port, DATAPATH_I_RF_OUT1_16_port, 
      DATAPATH_I_RF_OUT1_17_port, DATAPATH_I_RF_OUT1_18_port, 
      DATAPATH_I_RF_OUT1_19_port, DATAPATH_I_RF_OUT1_20_port, 
      DATAPATH_I_RF_OUT1_21_port, DATAPATH_I_RF_OUT1_22_port, 
      DATAPATH_I_RF_OUT1_23_port, DATAPATH_I_RF_OUT1_24_port, 
      DATAPATH_I_RF_OUT1_25_port, DATAPATH_I_RF_OUT1_26_port, 
      DATAPATH_I_RF_OUT1_27_port, DATAPATH_I_RF_OUT1_28_port, 
      DATAPATH_I_RF_OUT1_29_port, DATAPATH_I_RF_OUT1_30_port, 
      DATAPATH_I_RF_OUT1_31_port, DATAPATH_I_N414, DATAPATH_I_N413, 
      DATAPATH_I_N412, DATAPATH_I_N411, DATAPATH_I_N410, DATAPATH_I_N409, 
      DATAPATH_I_N408, DATAPATH_I_N407, DATAPATH_I_N406, DATAPATH_I_N405, 
      DATAPATH_I_N404, DATAPATH_I_N403, DATAPATH_I_N402, DATAPATH_I_N401, 
      DATAPATH_I_N400, DATAPATH_I_N399, DATAPATH_I_N398, DATAPATH_I_N397, 
      DATAPATH_I_N396, DATAPATH_I_N395, DATAPATH_I_N394, DATAPATH_I_N393, 
      DATAPATH_I_N392, DATAPATH_I_N391, DATAPATH_I_N390, DATAPATH_I_N389, 
      DATAPATH_I_N388, DATAPATH_I_N387, DATAPATH_I_N386, DATAPATH_I_N385, 
      DATAPATH_I_N384, DATAPATH_I_N383, DATAPATH_I_N382, DATAPATH_I_N381, 
      DATAPATH_I_N380, DATAPATH_I_N379, DATAPATH_I_N378, DATAPATH_I_N312, 
      DATAPATH_I_N311, DATAPATH_I_N310, DATAPATH_I_N309, DATAPATH_I_N308, 
      DATAPATH_I_N306, DATAPATH_I_N305, DATAPATH_I_N304, DATAPATH_I_N303, 
      DATAPATH_I_N302, DATAPATH_I_N301, DATAPATH_I_N300, DATAPATH_I_N299, 
      DATAPATH_I_N298, DATAPATH_I_N297, DATAPATH_I_N296, DATAPATH_I_N295, 
      DATAPATH_I_N294, DATAPATH_I_N293, DATAPATH_I_N292, DATAPATH_I_N291, 
      DATAPATH_I_N290, DATAPATH_I_N289, DATAPATH_I_N288, DATAPATH_I_N287, 
      DATAPATH_I_N286, DATAPATH_I_N285, DATAPATH_I_N284, DATAPATH_I_N283, 
      DATAPATH_I_N282, DATAPATH_I_N281, DATAPATH_I_N280, DATAPATH_I_N279, 
      DATAPATH_I_N278, DATAPATH_I_N277, DATAPATH_I_N276, DATAPATH_I_N275, 
      DATAPATH_I_N274, DATAPATH_I_N273, DATAPATH_I_N272, DATAPATH_I_N271, 
      DATAPATH_I_N270, DATAPATH_I_N269, DATAPATH_I_N268, DATAPATH_I_N267, 
      DATAPATH_I_N266, DATAPATH_I_N265, DATAPATH_I_N264, DATAPATH_I_N263, 
      DATAPATH_I_N262, DATAPATH_I_N261, DATAPATH_I_N260, DATAPATH_I_N259, 
      DATAPATH_I_N258, DATAPATH_I_N257, DATAPATH_I_N256, DATAPATH_I_N255, 
      DATAPATH_I_N254, DATAPATH_I_N253, DATAPATH_I_N252, DATAPATH_I_N251, 
      DATAPATH_I_N250, DATAPATH_I_N249, DATAPATH_I_N248, DATAPATH_I_N247, 
      DATAPATH_I_N246, DATAPATH_I_N245, DATAPATH_I_N244, DATAPATH_I_N243, 
      DATAPATH_I_N177, DATAPATH_I_N176, DATAPATH_I_N175, DATAPATH_I_N174, 
      DATAPATH_I_N173, DATAPATH_I_N172, DATAPATH_I_N171, DATAPATH_I_N170, 
      DATAPATH_I_N169, DATAPATH_I_N168, DATAPATH_I_N167, DATAPATH_I_N166, 
      DATAPATH_I_N165, DATAPATH_I_N164, DATAPATH_I_N163, DATAPATH_I_N162, 
      DATAPATH_I_N161, DATAPATH_I_N160, DATAPATH_I_N159, DATAPATH_I_N158, 
      DATAPATH_I_N157, DATAPATH_I_N156, DATAPATH_I_N155, DATAPATH_I_N154, 
      DATAPATH_I_N153, DATAPATH_I_N152, DATAPATH_I_N151, DATAPATH_I_N150, 
      DATAPATH_I_N149, DATAPATH_I_N148, DATAPATH_I_N147, DATAPATH_I_N146, 
      DATAPATH_I_N145, DATAPATH_I_N144, DATAPATH_I_N143, DATAPATH_I_N142, 
      DATAPATH_I_N141, DATAPATH_I_N140, DATAPATH_I_N139, DATAPATH_I_N138, 
      DATAPATH_I_N137, DATAPATH_I_N136, DATAPATH_I_N135, DATAPATH_I_N134, 
      DATAPATH_I_N133, DATAPATH_I_N132, DATAPATH_I_N131, DATAPATH_I_N130, 
      DATAPATH_I_N129, DATAPATH_I_N128, DATAPATH_I_N127, DATAPATH_I_N126, 
      DATAPATH_I_N125, DATAPATH_I_N124, DATAPATH_I_N123, DATAPATH_I_N122, 
      DATAPATH_I_N121, DATAPATH_I_N120, DATAPATH_I_N119, DATAPATH_I_N118, 
      DATAPATH_I_N117, DATAPATH_I_N116, DATAPATH_I_N115, DATAPATH_I_N114, 
      DATAPATH_I_N113, DATAPATH_I_N112, DATAPATH_I_N111, DATAPATH_I_N110, 
      DATAPATH_I_N109, DATAPATH_I_N65, DATAPATH_I_N64, DATAPATH_I_N63, 
      DATAPATH_I_N62, DATAPATH_I_N61, DATAPATH_I_N60, DATAPATH_I_N59, 
      DATAPATH_I_N58, DATAPATH_I_N57, DATAPATH_I_N56, DATAPATH_I_N55, 
      DATAPATH_I_N54, DATAPATH_I_N53, DATAPATH_I_N52, DATAPATH_I_N51, 
      DATAPATH_I_N50, DATAPATH_I_N49, DATAPATH_I_N48, DATAPATH_I_N47, 
      DATAPATH_I_N46, DATAPATH_I_N45, DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_0_port
      , DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_1_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_2_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_3_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_4_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_5_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_6_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_7_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_8_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_9_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_10_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_11_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_12_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_13_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_14_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_15_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_16_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_17_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_18_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_19_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_20_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_21_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_22_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_23_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_24_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_25_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_26_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_27_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_28_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_29_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_30_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_31_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_0_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_1_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_2_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_3_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_4_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_5_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_6_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_7_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_8_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_9_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_10_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_11_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_12_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_13_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_14_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_15_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_16_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_17_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_18_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_19_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_20_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_21_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_22_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_23_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_24_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_25_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_26_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_27_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_28_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_29_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_30_port, 
      DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_31_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_0_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_1_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_2_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_3_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_4_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_5_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_6_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_7_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_8_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_9_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_10_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_11_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_12_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_13_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_14_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_15_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_16_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_17_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_18_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_19_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_20_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_21_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_22_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_23_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_24_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_25_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_26_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_27_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_28_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_29_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_30_port, 
      DATAPATH_I_ID_EX_RF_OUT2_NEXT_31_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_0_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_1_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_2_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_3_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_4_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_5_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_6_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_7_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_8_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_9_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_10_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_11_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_12_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_13_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_14_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_15_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_16_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_17_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_18_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_19_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_20_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_21_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_22_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_23_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_24_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_25_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_26_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_27_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_28_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_29_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_30_port, 
      DATAPATH_I_ID_EX_RF_OUT1_NEXT_31_port, DATAPATH_I_ID_EX_RS2_NEXT_0_port, 
      DATAPATH_I_ID_EX_RS2_NEXT_1_port, DATAPATH_I_ID_EX_RS2_NEXT_2_port, 
      DATAPATH_I_ID_EX_RS2_NEXT_3_port, DATAPATH_I_ID_EX_RS2_NEXT_4_port, 
      DATAPATH_I_ID_EX_RS1_NEXT_0_port, DATAPATH_I_ID_EX_RS1_NEXT_1_port, 
      DATAPATH_I_ID_EX_RS1_NEXT_2_port, DATAPATH_I_ID_EX_RS1_NEXT_3_port, 
      DATAPATH_I_ID_EX_RS1_NEXT_4_port, DATAPATH_I_MEM_WB_RD_0_port, 
      DATAPATH_I_MEM_WB_RD_1_port, DATAPATH_I_MEM_WB_RD_2_port, 
      DATAPATH_I_MEM_WB_RD_3_port, DATAPATH_I_MEM_WB_RD_4_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_0_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_1_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_2_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_3_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_4_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_5_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_6_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_7_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_8_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_9_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_10_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_11_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_12_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_13_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_14_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_15_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_16_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_17_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_18_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_19_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_20_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_21_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_22_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_23_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_24_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_25_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_26_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_27_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_28_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_29_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_30_port, 
      DATAPATH_I_MEM_WB_DRAM_OUTPUT_31_port, DATAPATH_I_MEM_WB_RF_WE, 
      DATAPATH_I_EX_MEM_RD_0_port, DATAPATH_I_EX_MEM_RD_1_port, 
      DATAPATH_I_EX_MEM_RD_2_port, DATAPATH_I_EX_MEM_RD_3_port, 
      DATAPATH_I_EX_MEM_RD_4_port, DATAPATH_I_ID_EX_RF_OUT2_0_port, 
      DATAPATH_I_ID_EX_RF_OUT2_1_port, DATAPATH_I_ID_EX_RF_OUT2_2_port, 
      DATAPATH_I_ID_EX_RF_OUT2_3_port, DATAPATH_I_ID_EX_RF_OUT2_4_port, 
      DATAPATH_I_ID_EX_RF_OUT2_5_port, DATAPATH_I_ID_EX_RF_OUT2_6_port, 
      DATAPATH_I_ID_EX_RF_OUT2_7_port, DATAPATH_I_ID_EX_RF_OUT2_8_port, 
      DATAPATH_I_ID_EX_RF_OUT2_9_port, DATAPATH_I_ID_EX_RF_OUT2_10_port, 
      DATAPATH_I_ID_EX_RF_OUT2_11_port, DATAPATH_I_ID_EX_RF_OUT2_12_port, 
      DATAPATH_I_ID_EX_RF_OUT2_13_port, DATAPATH_I_ID_EX_RF_OUT2_14_port, 
      DATAPATH_I_ID_EX_RF_OUT2_15_port, DATAPATH_I_ID_EX_RF_OUT2_16_port, 
      DATAPATH_I_ID_EX_RF_OUT2_17_port, DATAPATH_I_ID_EX_RF_OUT2_18_port, 
      DATAPATH_I_ID_EX_RF_OUT2_19_port, DATAPATH_I_ID_EX_RF_OUT2_20_port, 
      DATAPATH_I_ID_EX_RF_OUT2_21_port, DATAPATH_I_ID_EX_RF_OUT2_22_port, 
      DATAPATH_I_ID_EX_RF_OUT2_23_port, DATAPATH_I_ID_EX_RF_OUT2_24_port, 
      DATAPATH_I_ID_EX_RF_OUT2_25_port, DATAPATH_I_ID_EX_RF_OUT2_26_port, 
      DATAPATH_I_ID_EX_RF_OUT2_27_port, DATAPATH_I_ID_EX_RF_OUT2_28_port, 
      DATAPATH_I_ID_EX_RF_OUT2_29_port, DATAPATH_I_ID_EX_RF_OUT2_30_port, 
      DATAPATH_I_ID_EX_RF_OUT2_31_port, DATAPATH_I_ID_EX_RF_OUT1_0_port, 
      DATAPATH_I_ID_EX_RF_OUT1_1_port, DATAPATH_I_ID_EX_RF_OUT1_2_port, 
      DATAPATH_I_ID_EX_RF_OUT1_3_port, DATAPATH_I_ID_EX_RF_OUT1_4_port, 
      DATAPATH_I_ID_EX_RF_OUT1_5_port, DATAPATH_I_ID_EX_RF_OUT1_6_port, 
      DATAPATH_I_ID_EX_RF_OUT1_7_port, DATAPATH_I_ID_EX_RF_OUT1_8_port, 
      DATAPATH_I_ID_EX_RF_OUT1_9_port, DATAPATH_I_ID_EX_RF_OUT1_10_port, 
      DATAPATH_I_ID_EX_RF_OUT1_11_port, DATAPATH_I_ID_EX_RF_OUT1_12_port, 
      DATAPATH_I_ID_EX_RF_OUT1_13_port, DATAPATH_I_ID_EX_RF_OUT1_14_port, 
      DATAPATH_I_ID_EX_RF_OUT1_15_port, DATAPATH_I_ID_EX_RF_OUT1_16_port, 
      DATAPATH_I_ID_EX_RF_OUT1_17_port, DATAPATH_I_ID_EX_RF_OUT1_18_port, 
      DATAPATH_I_ID_EX_RF_OUT1_19_port, DATAPATH_I_ID_EX_RF_OUT1_20_port, 
      DATAPATH_I_ID_EX_RF_OUT1_21_port, DATAPATH_I_ID_EX_RF_OUT1_22_port, 
      DATAPATH_I_ID_EX_RF_OUT1_23_port, DATAPATH_I_ID_EX_RF_OUT1_24_port, 
      DATAPATH_I_ID_EX_RF_OUT1_25_port, DATAPATH_I_ID_EX_RF_OUT1_26_port, 
      DATAPATH_I_ID_EX_RF_OUT1_27_port, DATAPATH_I_ID_EX_RF_OUT1_28_port, 
      DATAPATH_I_ID_EX_RF_OUT1_29_port, DATAPATH_I_ID_EX_RF_OUT1_30_port, 
      DATAPATH_I_ID_EX_RF_OUT1_31_port, DATAPATH_I_ID_EX_RD_0_port, 
      DATAPATH_I_ID_EX_RD_1_port, DATAPATH_I_ID_EX_RD_2_port, 
      DATAPATH_I_ID_EX_RD_3_port, DATAPATH_I_ID_EX_RD_4_port, 
      DATAPATH_I_IF_ID_IR_11_port, DATAPATH_I_IF_ID_IR_12_port, 
      DATAPATH_I_IF_ID_IR_13_port, DATAPATH_I_IF_ID_IR_14_port, 
      DATAPATH_I_IF_ID_IR_15_port, DATAPATH_I_IF_ID_IR_16_port, 
      DATAPATH_I_IF_ID_IR_17_port, DATAPATH_I_IF_ID_IR_18_port, 
      DATAPATH_I_IF_ID_IR_19_port, DATAPATH_I_IF_ID_IR_20_port, 
      DATAPATH_I_IF_ID_IR_21_port, DATAPATH_I_IF_ID_IR_22_port, 
      DATAPATH_I_IF_ID_IR_23_port, DATAPATH_I_IF_ID_IR_24_port, 
      DATAPATH_I_IF_ID_IR_25_port, DATAPATH_I_IF_ID_IR_26_port, 
      DATAPATH_I_IF_ID_IR_27_port, DATAPATH_I_IF_ID_IR_28_port, 
      DATAPATH_I_IF_ID_IR_29_port, DATAPATH_I_IF_ID_IR_30_port, 
      DATAPATH_I_IF_ID_IR_31_port, DATAPATH_I_n29, DATAPATH_I_n28, 
      DATAPATH_I_n27, DATAPATH_I_n26, DATAPATH_I_n25, DATAPATH_I_n24, 
      DATAPATH_I_n23, DATAPATH_I_n22, DATAPATH_I_n21, DATAPATH_I_n20, 
      DATAPATH_I_n19, DATAPATH_I_n18, DATAPATH_I_n17, DATAPATH_I_n16, 
      DATAPATH_I_n15, DATAPATH_I_LATCH_LMD_LDI_0_N3, 
      DATAPATH_I_LATCH_LMD_LDI_1_N3, DATAPATH_I_LATCH_LMD_LDI_2_N3, 
      DATAPATH_I_LATCH_LMD_LDI_3_N3, DATAPATH_I_LATCH_LMD_LDI_4_N3, 
      DATAPATH_I_LATCH_LMD_LDI_5_N3, DATAPATH_I_LATCH_LMD_LDI_6_N3, 
      DATAPATH_I_LATCH_LMD_LDI_7_N3, DATAPATH_I_LATCH_LMD_LDI_8_N3, 
      DATAPATH_I_LATCH_LMD_LDI_9_N3, DATAPATH_I_LATCH_LMD_LDI_10_N3, 
      DATAPATH_I_LATCH_LMD_LDI_11_N3, DATAPATH_I_LATCH_LMD_LDI_12_N3, 
      DATAPATH_I_LATCH_LMD_LDI_13_N3, DATAPATH_I_LATCH_LMD_LDI_14_N3, 
      DATAPATH_I_LATCH_LMD_LDI_15_N3, DATAPATH_I_LATCH_LMD_LDI_16_N3, 
      DATAPATH_I_LATCH_LMD_LDI_17_N3, DATAPATH_I_LATCH_LMD_LDI_18_N3, 
      DATAPATH_I_LATCH_LMD_LDI_19_N3, DATAPATH_I_LATCH_LMD_LDI_20_N3, 
      DATAPATH_I_LATCH_LMD_LDI_21_N3, DATAPATH_I_LATCH_LMD_LDI_22_N3, 
      DATAPATH_I_LATCH_LMD_LDI_23_N3, DATAPATH_I_LATCH_LMD_LDI_24_N3, 
      DATAPATH_I_LATCH_LMD_LDI_25_N3, DATAPATH_I_LATCH_LMD_LDI_26_N3, 
      DATAPATH_I_LATCH_LMD_LDI_27_N3, DATAPATH_I_LATCH_LMD_LDI_28_N3, 
      DATAPATH_I_LATCH_LMD_LDI_29_N3, DATAPATH_I_LATCH_LMD_LDI_30_N3, 
      DATAPATH_I_LATCH_LMD_LDI_31_N3, DATAPATH_I_LATCH_ALUOUT_LDI_0_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_1_N3, DATAPATH_I_LATCH_ALUOUT_LDI_2_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_3_N3, DATAPATH_I_LATCH_ALUOUT_LDI_4_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_5_N3, DATAPATH_I_LATCH_ALUOUT_LDI_6_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_7_N3, DATAPATH_I_LATCH_ALUOUT_LDI_8_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_9_N3, DATAPATH_I_LATCH_ALUOUT_LDI_10_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_11_N3, DATAPATH_I_LATCH_ALUOUT_LDI_12_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_13_N3, DATAPATH_I_LATCH_ALUOUT_LDI_14_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_15_N3, DATAPATH_I_LATCH_ALUOUT_LDI_16_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_17_N3, DATAPATH_I_LATCH_ALUOUT_LDI_18_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_19_N3, DATAPATH_I_LATCH_ALUOUT_LDI_20_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_21_N3, DATAPATH_I_LATCH_ALUOUT_LDI_22_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_23_N3, DATAPATH_I_LATCH_ALUOUT_LDI_24_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_25_N3, DATAPATH_I_LATCH_ALUOUT_LDI_26_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_27_N3, DATAPATH_I_LATCH_ALUOUT_LDI_28_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_29_N3, DATAPATH_I_LATCH_ALUOUT_LDI_30_N3, 
      DATAPATH_I_LATCH_ALUOUT_LDI_31_N3, DATAPATH_I_LATCH_RF2_LDI_0_N3, 
      DATAPATH_I_LATCH_RF2_LDI_1_N3, DATAPATH_I_LATCH_RF2_LDI_2_N3, 
      DATAPATH_I_LATCH_RF2_LDI_3_N3, DATAPATH_I_LATCH_RF2_LDI_4_N3, 
      DATAPATH_I_LATCH_RF2_LDI_5_N3, DATAPATH_I_LATCH_RF2_LDI_6_N3, 
      DATAPATH_I_LATCH_RF2_LDI_7_N3, DATAPATH_I_LATCH_RF2_LDI_8_N3, 
      DATAPATH_I_LATCH_RF2_LDI_9_N3, DATAPATH_I_LATCH_RF2_LDI_10_N3, 
      DATAPATH_I_LATCH_RF2_LDI_11_N3, DATAPATH_I_LATCH_RF2_LDI_12_N3, 
      DATAPATH_I_LATCH_RF2_LDI_13_N3, DATAPATH_I_LATCH_RF2_LDI_14_N3, 
      DATAPATH_I_LATCH_RF2_LDI_15_N3, DATAPATH_I_LATCH_RF2_LDI_16_N3, 
      DATAPATH_I_LATCH_RF2_LDI_17_N3, DATAPATH_I_LATCH_RF2_LDI_18_N3, 
      DATAPATH_I_LATCH_RF2_LDI_19_N3, DATAPATH_I_LATCH_RF2_LDI_20_N3, 
      DATAPATH_I_LATCH_RF2_LDI_21_N3, DATAPATH_I_LATCH_RF2_LDI_22_N3, 
      DATAPATH_I_LATCH_RF2_LDI_23_N3, DATAPATH_I_LATCH_RF2_LDI_24_N3, 
      DATAPATH_I_LATCH_RF2_LDI_25_N3, DATAPATH_I_LATCH_RF2_LDI_26_N3, 
      DATAPATH_I_LATCH_RF2_LDI_27_N3, DATAPATH_I_LATCH_RF2_LDI_28_N3, 
      DATAPATH_I_LATCH_RF2_LDI_29_N3, DATAPATH_I_LATCH_RF2_LDI_30_N3, 
      DATAPATH_I_LATCH_RF2_LDI_31_N3, DATAPATH_I_LATCH_RF1_LDI_0_N3, 
      DATAPATH_I_LATCH_RF1_LDI_1_N3, DATAPATH_I_LATCH_RF1_LDI_2_N3, 
      DATAPATH_I_LATCH_RF1_LDI_3_N3, DATAPATH_I_LATCH_RF1_LDI_4_N3, 
      DATAPATH_I_LATCH_RF1_LDI_5_N3, DATAPATH_I_LATCH_RF1_LDI_6_N3, 
      DATAPATH_I_LATCH_RF1_LDI_7_N3, DATAPATH_I_LATCH_RF1_LDI_8_N3, 
      DATAPATH_I_LATCH_RF1_LDI_9_N3, DATAPATH_I_LATCH_RF1_LDI_10_N3, 
      DATAPATH_I_LATCH_RF1_LDI_11_N3, DATAPATH_I_LATCH_RF1_LDI_12_N3, 
      DATAPATH_I_LATCH_RF1_LDI_13_N3, DATAPATH_I_LATCH_RF1_LDI_14_N3, 
      DATAPATH_I_LATCH_RF1_LDI_15_N3, DATAPATH_I_LATCH_RF1_LDI_16_N3, 
      DATAPATH_I_LATCH_RF1_LDI_17_N3, DATAPATH_I_LATCH_RF1_LDI_18_N3, 
      DATAPATH_I_LATCH_RF1_LDI_19_N3, DATAPATH_I_LATCH_RF1_LDI_20_N3, 
      DATAPATH_I_LATCH_RF1_LDI_21_N3, DATAPATH_I_LATCH_RF1_LDI_22_N3, 
      DATAPATH_I_LATCH_RF1_LDI_23_N3, DATAPATH_I_LATCH_RF1_LDI_24_N3, 
      DATAPATH_I_LATCH_RF1_LDI_25_N3, DATAPATH_I_LATCH_RF1_LDI_26_N3, 
      DATAPATH_I_LATCH_RF1_LDI_27_N3, DATAPATH_I_LATCH_RF1_LDI_28_N3, 
      DATAPATH_I_LATCH_RF1_LDI_29_N3, DATAPATH_I_LATCH_RF1_LDI_30_N3, 
      DATAPATH_I_LATCH_RF1_LDI_31_N3, DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_N3,
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_N3, 
      DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_N3, n285, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, 
      n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, 
      n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
      n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, 
      n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, 
      n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, 
      n441, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, 
      n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, 
      n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, 
      n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, 
      n_1377, n_1378, n_1379 : std_logic;

begin
   
   IRAM_I : DLX_IRAM_RAM_DEPTH256_I_SIZE32 port map( RST => RST, ADDR(31) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(30) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(29) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(28) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(27) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(26) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(25) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(24) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(23) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(22) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(21) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(20) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(19) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(18) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(17) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(16) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(15) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(14) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(13) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(12) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(11) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(10) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(9) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(8) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(7) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(6) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(5) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(4) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(3) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(2) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(1) => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(0) => 
                           DATAPATH_I_MEM_WB_RF_WE, DOUT(31) => IR_BUS_31_port,
                           DOUT(30) => IR_BUS_30_port, DOUT(29) => 
                           IR_BUS_29_port, DOUT(28) => IR_BUS_28_port, DOUT(27)
                           => IR_BUS_27_port, DOUT(26) => IR_BUS_26_port, 
                           DOUT(25) => IR_BUS_25_port, DOUT(24) => 
                           IR_BUS_24_port, DOUT(23) => IR_BUS_23_port, DOUT(22)
                           => IR_BUS_22_port, DOUT(21) => IR_BUS_21_port, 
                           DOUT(20) => IR_BUS_20_port, DOUT(19) => 
                           IR_BUS_19_port, DOUT(18) => IR_BUS_18_port, DOUT(17)
                           => IR_BUS_17_port, DOUT(16) => IR_BUS_16_port, 
                           DOUT(15) => IR_BUS_15_port, DOUT(14) => 
                           IR_BUS_14_port, DOUT(13) => IR_BUS_13_port, DOUT(12)
                           => IR_BUS_12_port, DOUT(11) => IR_BUS_11_port, 
                           DOUT(10) => IR_BUS_10_port, DOUT(9) => IR_BUS_9_port
                           , DOUT(8) => IR_BUS_8_port, DOUT(7) => IR_BUS_7_port
                           , DOUT(6) => IR_BUS_6_port, DOUT(5) => IR_BUS_5_port
                           , DOUT(4) => IR_BUS_4_port, DOUT(3) => IR_BUS_3_port
                           , DOUT(2) => IR_BUS_2_port, DOUT(1) => IR_BUS_1_port
                           , DOUT(0) => IR_BUS_0_port);
   DRAM_I : DLX_DRAM_N256_NW32 port map( CLK => CLK, RST => RST, RE => 
                           DATAPATH_I_MEM_WB_RF_WE, WE => 
                           DATAPATH_I_MEM_WB_RF_WE, ADDR(31) => 
                           DATA_ADDR_31_port, ADDR(30) => DATA_ADDR_30_port, 
                           ADDR(29) => DATA_ADDR_29_port, ADDR(28) => 
                           DATA_ADDR_28_port, ADDR(27) => DATA_ADDR_27_port, 
                           ADDR(26) => DATA_ADDR_26_port, ADDR(25) => 
                           DATA_ADDR_25_port, ADDR(24) => DATA_ADDR_24_port, 
                           ADDR(23) => DATA_ADDR_23_port, ADDR(22) => 
                           DATA_ADDR_22_port, ADDR(21) => DATA_ADDR_21_port, 
                           ADDR(20) => DATA_ADDR_20_port, ADDR(19) => 
                           DATA_ADDR_19_port, ADDR(18) => DATA_ADDR_18_port, 
                           ADDR(17) => DATA_ADDR_17_port, ADDR(16) => 
                           DATA_ADDR_16_port, ADDR(15) => DATA_ADDR_15_port, 
                           ADDR(14) => DATA_ADDR_14_port, ADDR(13) => 
                           DATA_ADDR_13_port, ADDR(12) => DATA_ADDR_12_port, 
                           ADDR(11) => DATA_ADDR_11_port, ADDR(10) => 
                           DATA_ADDR_10_port, ADDR(9) => DATA_ADDR_9_port, 
                           ADDR(8) => DATA_ADDR_8_port, ADDR(7) => 
                           DATA_ADDR_7_port, ADDR(6) => DATA_ADDR_6_port, 
                           ADDR(5) => DATA_ADDR_5_port, ADDR(4) => 
                           DATA_ADDR_4_port, ADDR(3) => DATA_ADDR_3_port, 
                           ADDR(2) => DATA_ADDR_2_port, ADDR(1) => 
                           DATA_ADDR_1_port, ADDR(0) => DATA_ADDR_0_port, 
                           DIN(31) => DATA_IN_31_port, DIN(30) => 
                           DATA_IN_30_port, DIN(29) => DATA_IN_29_port, DIN(28)
                           => DATA_IN_28_port, DIN(27) => DATA_IN_27_port, 
                           DIN(26) => DATA_IN_26_port, DIN(25) => 
                           DATA_IN_25_port, DIN(24) => DATA_IN_24_port, DIN(23)
                           => DATA_IN_23_port, DIN(22) => DATA_IN_22_port, 
                           DIN(21) => DATA_IN_21_port, DIN(20) => 
                           DATA_IN_20_port, DIN(19) => DATA_IN_19_port, DIN(18)
                           => DATA_IN_18_port, DIN(17) => DATA_IN_17_port, 
                           DIN(16) => DATA_IN_16_port, DIN(15) => 
                           DATA_IN_15_port, DIN(14) => DATA_IN_14_port, DIN(13)
                           => DATA_IN_13_port, DIN(12) => DATA_IN_12_port, 
                           DIN(11) => DATA_IN_11_port, DIN(10) => 
                           DATA_IN_10_port, DIN(9) => DATA_IN_9_port, DIN(8) =>
                           DATA_IN_8_port, DIN(7) => DATA_IN_7_port, DIN(6) => 
                           DATA_IN_6_port, DIN(5) => DATA_IN_5_port, DIN(4) => 
                           DATA_IN_4_port, DIN(3) => DATA_IN_3_port, DIN(2) => 
                           DATA_IN_2_port, DIN(1) => DATA_IN_1_port, DIN(0) => 
                           DATA_IN_0_port, DOUT(31) => DATA_OUT_31_port, 
                           DOUT(30) => DATA_OUT_30_port, DOUT(29) => 
                           DATA_OUT_29_port, DOUT(28) => DATA_OUT_28_port, 
                           DOUT(27) => DATA_OUT_27_port, DOUT(26) => 
                           DATA_OUT_26_port, DOUT(25) => DATA_OUT_25_port, 
                           DOUT(24) => DATA_OUT_24_port, DOUT(23) => 
                           DATA_OUT_23_port, DOUT(22) => DATA_OUT_22_port, 
                           DOUT(21) => DATA_OUT_21_port, DOUT(20) => 
                           DATA_OUT_20_port, DOUT(19) => DATA_OUT_19_port, 
                           DOUT(18) => DATA_OUT_18_port, DOUT(17) => 
                           DATA_OUT_17_port, DOUT(16) => DATA_OUT_16_port, 
                           DOUT(15) => DATA_OUT_15_port, DOUT(14) => 
                           DATA_OUT_14_port, DOUT(13) => DATA_OUT_13_port, 
                           DOUT(12) => DATA_OUT_12_port, DOUT(11) => 
                           DATA_OUT_11_port, DOUT(10) => DATA_OUT_10_port, 
                           DOUT(9) => DATA_OUT_9_port, DOUT(8) => 
                           DATA_OUT_8_port, DOUT(7) => DATA_OUT_7_port, DOUT(6)
                           => DATA_OUT_6_port, DOUT(5) => DATA_OUT_5_port, 
                           DOUT(4) => DATA_OUT_4_port, DOUT(3) => 
                           DATA_OUT_3_port, DOUT(2) => DATA_OUT_2_port, DOUT(1)
                           => DATA_OUT_1_port, DOUT(0) => DATA_OUT_0_port);
   DATAPATH_I_ARITHMETIC_LOGIC_UNIT : ALU_N32_NB8 port map( OP1(31) => 
                           DATAPATH_I_ID_EX_RF_OUT1_31_port, OP1(30) => 
                           DATAPATH_I_ID_EX_RF_OUT1_30_port, OP1(29) => 
                           DATAPATH_I_ID_EX_RF_OUT1_29_port, OP1(28) => 
                           DATAPATH_I_ID_EX_RF_OUT1_28_port, OP1(27) => 
                           DATAPATH_I_ID_EX_RF_OUT1_27_port, OP1(26) => 
                           DATAPATH_I_ID_EX_RF_OUT1_26_port, OP1(25) => 
                           DATAPATH_I_ID_EX_RF_OUT1_25_port, OP1(24) => 
                           DATAPATH_I_ID_EX_RF_OUT1_24_port, OP1(23) => 
                           DATAPATH_I_ID_EX_RF_OUT1_23_port, OP1(22) => 
                           DATAPATH_I_ID_EX_RF_OUT1_22_port, OP1(21) => 
                           DATAPATH_I_ID_EX_RF_OUT1_21_port, OP1(20) => 
                           DATAPATH_I_ID_EX_RF_OUT1_20_port, OP1(19) => 
                           DATAPATH_I_ID_EX_RF_OUT1_19_port, OP1(18) => 
                           DATAPATH_I_ID_EX_RF_OUT1_18_port, OP1(17) => 
                           DATAPATH_I_ID_EX_RF_OUT1_17_port, OP1(16) => 
                           DATAPATH_I_ID_EX_RF_OUT1_16_port, OP1(15) => 
                           DATAPATH_I_ID_EX_RF_OUT1_15_port, OP1(14) => 
                           DATAPATH_I_ID_EX_RF_OUT1_14_port, OP1(13) => 
                           DATAPATH_I_ID_EX_RF_OUT1_13_port, OP1(12) => 
                           DATAPATH_I_ID_EX_RF_OUT1_12_port, OP1(11) => 
                           DATAPATH_I_ID_EX_RF_OUT1_11_port, OP1(10) => 
                           DATAPATH_I_ID_EX_RF_OUT1_10_port, OP1(9) => 
                           DATAPATH_I_ID_EX_RF_OUT1_9_port, OP1(8) => 
                           DATAPATH_I_ID_EX_RF_OUT1_8_port, OP1(7) => 
                           DATAPATH_I_ID_EX_RF_OUT1_7_port, OP1(6) => 
                           DATAPATH_I_ID_EX_RF_OUT1_6_port, OP1(5) => 
                           DATAPATH_I_ID_EX_RF_OUT1_5_port, OP1(4) => 
                           DATAPATH_I_ID_EX_RF_OUT1_4_port, OP1(3) => 
                           DATAPATH_I_ID_EX_RF_OUT1_3_port, OP1(2) => 
                           DATAPATH_I_ID_EX_RF_OUT1_2_port, OP1(1) => 
                           DATAPATH_I_ID_EX_RF_OUT1_1_port, OP1(0) => 
                           DATAPATH_I_ID_EX_RF_OUT1_0_port, OP2(31) => 
                           DATAPATH_I_ID_EX_RF_OUT2_31_port, OP2(30) => 
                           DATAPATH_I_ID_EX_RF_OUT2_30_port, OP2(29) => 
                           DATAPATH_I_ID_EX_RF_OUT2_29_port, OP2(28) => 
                           DATAPATH_I_ID_EX_RF_OUT2_28_port, OP2(27) => 
                           DATAPATH_I_ID_EX_RF_OUT2_27_port, OP2(26) => 
                           DATAPATH_I_ID_EX_RF_OUT2_26_port, OP2(25) => 
                           DATAPATH_I_ID_EX_RF_OUT2_25_port, OP2(24) => 
                           DATAPATH_I_ID_EX_RF_OUT2_24_port, OP2(23) => 
                           DATAPATH_I_ID_EX_RF_OUT2_23_port, OP2(22) => 
                           DATAPATH_I_ID_EX_RF_OUT2_22_port, OP2(21) => 
                           DATAPATH_I_ID_EX_RF_OUT2_21_port, OP2(20) => 
                           DATAPATH_I_ID_EX_RF_OUT2_20_port, OP2(19) => 
                           DATAPATH_I_ID_EX_RF_OUT2_19_port, OP2(18) => 
                           DATAPATH_I_ID_EX_RF_OUT2_18_port, OP2(17) => 
                           DATAPATH_I_ID_EX_RF_OUT2_17_port, OP2(16) => 
                           DATAPATH_I_ID_EX_RF_OUT2_16_port, OP2(15) => 
                           DATAPATH_I_ID_EX_RF_OUT2_15_port, OP2(14) => 
                           DATAPATH_I_ID_EX_RF_OUT2_14_port, OP2(13) => 
                           DATAPATH_I_ID_EX_RF_OUT2_13_port, OP2(12) => 
                           DATAPATH_I_ID_EX_RF_OUT2_12_port, OP2(11) => 
                           DATAPATH_I_ID_EX_RF_OUT2_11_port, OP2(10) => 
                           DATAPATH_I_ID_EX_RF_OUT2_10_port, OP2(9) => 
                           DATAPATH_I_ID_EX_RF_OUT2_9_port, OP2(8) => 
                           DATAPATH_I_ID_EX_RF_OUT2_8_port, OP2(7) => 
                           DATAPATH_I_ID_EX_RF_OUT2_7_port, OP2(6) => 
                           DATAPATH_I_ID_EX_RF_OUT2_6_port, OP2(5) => 
                           DATAPATH_I_ID_EX_RF_OUT2_5_port, OP2(4) => 
                           DATAPATH_I_ID_EX_RF_OUT2_4_port, OP2(3) => 
                           DATAPATH_I_ID_EX_RF_OUT2_3_port, OP2(2) => 
                           DATAPATH_I_ID_EX_RF_OUT2_2_port, OP2(1) => 
                           DATAPATH_I_ID_EX_RF_OUT2_1_port, OP2(0) => 
                           DATAPATH_I_ID_EX_RF_OUT2_0_port, OPC(0) => 
                           ALU_OPCODE_i_0_port, OPC(1) => ALU_OPCODE_i_1_port, 
                           OPC(2) => ALU_OPCODE_i_2_port, OPC(3) => 
                           ALU_OPCODE_i_3_port, OPC(4) => ALU_OPCODE_i_4_port, 
                           OPC(5) => ALU_OPCODE_i_5_port, OPC(6) => 
                           ALU_OPCODE_i_6_port, Y(31) => 
                           DATAPATH_I_ALU_OUTPUT_31_port, Y(30) => 
                           DATAPATH_I_ALU_OUTPUT_30_port, Y(29) => 
                           DATAPATH_I_ALU_OUTPUT_29_port, Y(28) => 
                           DATAPATH_I_ALU_OUTPUT_28_port, Y(27) => 
                           DATAPATH_I_ALU_OUTPUT_27_port, Y(26) => 
                           DATAPATH_I_ALU_OUTPUT_26_port, Y(25) => 
                           DATAPATH_I_ALU_OUTPUT_25_port, Y(24) => 
                           DATAPATH_I_ALU_OUTPUT_24_port, Y(23) => 
                           DATAPATH_I_ALU_OUTPUT_23_port, Y(22) => 
                           DATAPATH_I_ALU_OUTPUT_22_port, Y(21) => 
                           DATAPATH_I_ALU_OUTPUT_21_port, Y(20) => 
                           DATAPATH_I_ALU_OUTPUT_20_port, Y(19) => 
                           DATAPATH_I_ALU_OUTPUT_19_port, Y(18) => 
                           DATAPATH_I_ALU_OUTPUT_18_port, Y(17) => 
                           DATAPATH_I_ALU_OUTPUT_17_port, Y(16) => 
                           DATAPATH_I_ALU_OUTPUT_16_port, Y(15) => 
                           DATAPATH_I_ALU_OUTPUT_15_port, Y(14) => 
                           DATAPATH_I_ALU_OUTPUT_14_port, Y(13) => 
                           DATAPATH_I_ALU_OUTPUT_13_port, Y(12) => 
                           DATAPATH_I_ALU_OUTPUT_12_port, Y(11) => 
                           DATAPATH_I_ALU_OUTPUT_11_port, Y(10) => 
                           DATAPATH_I_ALU_OUTPUT_10_port, Y(9) => 
                           DATAPATH_I_ALU_OUTPUT_9_port, Y(8) => 
                           DATAPATH_I_ALU_OUTPUT_8_port, Y(7) => 
                           DATAPATH_I_ALU_OUTPUT_7_port, Y(6) => 
                           DATAPATH_I_ALU_OUTPUT_6_port, Y(5) => 
                           DATAPATH_I_ALU_OUTPUT_5_port, Y(4) => 
                           DATAPATH_I_ALU_OUTPUT_4_port, Y(3) => 
                           DATAPATH_I_ALU_OUTPUT_3_port, Y(2) => 
                           DATAPATH_I_ALU_OUTPUT_2_port, Y(1) => 
                           DATAPATH_I_ALU_OUTPUT_1_port, Y(0) => 
                           DATAPATH_I_ALU_OUTPUT_0_port, Z => n_1171);
   DATAPATH_I_REGISTER_FILE : RF_N32_NA5 port map( RST => RST, EN => n285, 
                           EN_RD1 => n285, EN_RD2 => n285, EN_WR => 
                           DATAPATH_I_MEM_WB_RF_WE, ADD_RD1(4) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_4_port, ADD_RD1(3) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_3_port, ADD_RD1(2) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_2_port, ADD_RD1(1) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_1_port, ADD_RD1(0) => 
                           DATAPATH_I_ID_EX_RS1_NEXT_0_port, ADD_RD2(4) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_4_port, ADD_RD2(3) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_3_port, ADD_RD2(2) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_2_port, ADD_RD2(1) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_1_port, ADD_RD2(0) => 
                           DATAPATH_I_ID_EX_RS2_NEXT_0_port, ADD_WR(4) => 
                           DATAPATH_I_MEM_WB_RD_4_port, ADD_WR(3) => 
                           DATAPATH_I_MEM_WB_RD_3_port, ADD_WR(2) => 
                           DATAPATH_I_MEM_WB_RD_2_port, ADD_WR(1) => 
                           DATAPATH_I_MEM_WB_RD_1_port, ADD_WR(0) => 
                           DATAPATH_I_MEM_WB_RD_0_port, DATAIN(31) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_31_port, DATAIN(30) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_30_port, DATAIN(29) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_29_port, DATAIN(28) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_28_port, DATAIN(27) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_27_port, DATAIN(26) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_26_port, DATAIN(25) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_25_port, DATAIN(24) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_24_port, DATAIN(23) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_23_port, DATAIN(22) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_22_port, DATAIN(21) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_21_port, DATAIN(20) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_20_port, DATAIN(19) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_19_port, DATAIN(18) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_18_port, DATAIN(17) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_17_port, DATAIN(16) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_16_port, DATAIN(15) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_15_port, DATAIN(14) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_14_port, DATAIN(13) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_13_port, DATAIN(12) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_12_port, DATAIN(11) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_11_port, DATAIN(10) =>
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_10_port, DATAIN(9) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_9_port, DATAIN(8) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_8_port, DATAIN(7) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_7_port, DATAIN(6) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_6_port, DATAIN(5) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_5_port, DATAIN(4) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_4_port, DATAIN(3) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_3_port, DATAIN(2) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_2_port, DATAIN(1) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_1_port, DATAIN(0) => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_0_port, OUT1(31) => 
                           DATAPATH_I_RF_OUT1_31_port, OUT1(30) => 
                           DATAPATH_I_RF_OUT1_30_port, OUT1(29) => 
                           DATAPATH_I_RF_OUT1_29_port, OUT1(28) => 
                           DATAPATH_I_RF_OUT1_28_port, OUT1(27) => 
                           DATAPATH_I_RF_OUT1_27_port, OUT1(26) => 
                           DATAPATH_I_RF_OUT1_26_port, OUT1(25) => 
                           DATAPATH_I_RF_OUT1_25_port, OUT1(24) => 
                           DATAPATH_I_RF_OUT1_24_port, OUT1(23) => 
                           DATAPATH_I_RF_OUT1_23_port, OUT1(22) => 
                           DATAPATH_I_RF_OUT1_22_port, OUT1(21) => 
                           DATAPATH_I_RF_OUT1_21_port, OUT1(20) => 
                           DATAPATH_I_RF_OUT1_20_port, OUT1(19) => 
                           DATAPATH_I_RF_OUT1_19_port, OUT1(18) => 
                           DATAPATH_I_RF_OUT1_18_port, OUT1(17) => 
                           DATAPATH_I_RF_OUT1_17_port, OUT1(16) => 
                           DATAPATH_I_RF_OUT1_16_port, OUT1(15) => 
                           DATAPATH_I_RF_OUT1_15_port, OUT1(14) => 
                           DATAPATH_I_RF_OUT1_14_port, OUT1(13) => 
                           DATAPATH_I_RF_OUT1_13_port, OUT1(12) => 
                           DATAPATH_I_RF_OUT1_12_port, OUT1(11) => 
                           DATAPATH_I_RF_OUT1_11_port, OUT1(10) => 
                           DATAPATH_I_RF_OUT1_10_port, OUT1(9) => 
                           DATAPATH_I_RF_OUT1_9_port, OUT1(8) => 
                           DATAPATH_I_RF_OUT1_8_port, OUT1(7) => 
                           DATAPATH_I_RF_OUT1_7_port, OUT1(6) => 
                           DATAPATH_I_RF_OUT1_6_port, OUT1(5) => 
                           DATAPATH_I_RF_OUT1_5_port, OUT1(4) => 
                           DATAPATH_I_RF_OUT1_4_port, OUT1(3) => 
                           DATAPATH_I_RF_OUT1_3_port, OUT1(2) => 
                           DATAPATH_I_RF_OUT1_2_port, OUT1(1) => 
                           DATAPATH_I_RF_OUT1_1_port, OUT1(0) => 
                           DATAPATH_I_RF_OUT1_0_port, OUT2(31) => 
                           DATAPATH_I_RF_OUT2_31_port, OUT2(30) => 
                           DATAPATH_I_RF_OUT2_30_port, OUT2(29) => 
                           DATAPATH_I_RF_OUT2_29_port, OUT2(28) => 
                           DATAPATH_I_RF_OUT2_28_port, OUT2(27) => 
                           DATAPATH_I_RF_OUT2_27_port, OUT2(26) => 
                           DATAPATH_I_RF_OUT2_26_port, OUT2(25) => 
                           DATAPATH_I_RF_OUT2_25_port, OUT2(24) => 
                           DATAPATH_I_RF_OUT2_24_port, OUT2(23) => 
                           DATAPATH_I_RF_OUT2_23_port, OUT2(22) => 
                           DATAPATH_I_RF_OUT2_22_port, OUT2(21) => 
                           DATAPATH_I_RF_OUT2_21_port, OUT2(20) => 
                           DATAPATH_I_RF_OUT2_20_port, OUT2(19) => 
                           DATAPATH_I_RF_OUT2_19_port, OUT2(18) => 
                           DATAPATH_I_RF_OUT2_18_port, OUT2(17) => 
                           DATAPATH_I_RF_OUT2_17_port, OUT2(16) => 
                           DATAPATH_I_RF_OUT2_16_port, OUT2(15) => 
                           DATAPATH_I_RF_OUT2_15_port, OUT2(14) => 
                           DATAPATH_I_RF_OUT2_14_port, OUT2(13) => 
                           DATAPATH_I_RF_OUT2_13_port, OUT2(12) => 
                           DATAPATH_I_RF_OUT2_12_port, OUT2(11) => 
                           DATAPATH_I_RF_OUT2_11_port, OUT2(10) => 
                           DATAPATH_I_RF_OUT2_10_port, OUT2(9) => 
                           DATAPATH_I_RF_OUT2_9_port, OUT2(8) => 
                           DATAPATH_I_RF_OUT2_8_port, OUT2(7) => 
                           DATAPATH_I_RF_OUT2_7_port, OUT2(6) => 
                           DATAPATH_I_RF_OUT2_6_port, OUT2(5) => 
                           DATAPATH_I_RF_OUT2_5_port, OUT2(4) => 
                           DATAPATH_I_RF_OUT2_4_port, OUT2(3) => 
                           DATAPATH_I_RF_OUT2_3_port, OUT2(2) => 
                           DATAPATH_I_RF_OUT2_2_port, OUT2(1) => 
                           DATAPATH_I_RF_OUT2_1_port, OUT2(0) => 
                           DATAPATH_I_RF_OUT2_0_port);
   DATAPATH_I_IF_ID_IR_reg_11_inst : DFF_X1 port map( D => DATAPATH_I_N45, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_11_port, QN => 
                           n_1172);
   DATAPATH_I_IF_ID_IR_reg_12_inst : DFF_X1 port map( D => DATAPATH_I_N46, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_12_port, QN => 
                           n_1173);
   DATAPATH_I_IF_ID_IR_reg_13_inst : DFF_X1 port map( D => DATAPATH_I_N47, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_13_port, QN => 
                           n_1174);
   DATAPATH_I_IF_ID_IR_reg_14_inst : DFF_X1 port map( D => DATAPATH_I_N48, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_14_port, QN => 
                           n_1175);
   DATAPATH_I_IF_ID_IR_reg_15_inst : DFF_X1 port map( D => DATAPATH_I_N49, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_15_port, QN => 
                           n_1176);
   DATAPATH_I_IF_ID_IR_reg_16_inst : DFF_X1 port map( D => DATAPATH_I_N50, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_16_port, QN => 
                           n_1177);
   DATAPATH_I_IF_ID_IR_reg_17_inst : DFF_X1 port map( D => DATAPATH_I_N51, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_17_port, QN => 
                           n_1178);
   DATAPATH_I_IF_ID_IR_reg_18_inst : DFF_X1 port map( D => DATAPATH_I_N52, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_18_port, QN => 
                           n_1179);
   DATAPATH_I_IF_ID_IR_reg_19_inst : DFF_X1 port map( D => DATAPATH_I_N53, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_19_port, QN => 
                           n_1180);
   DATAPATH_I_IF_ID_IR_reg_20_inst : DFF_X1 port map( D => DATAPATH_I_N54, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_20_port, QN => 
                           n_1181);
   DATAPATH_I_IF_ID_IR_reg_21_inst : DFF_X1 port map( D => DATAPATH_I_N55, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_21_port, QN => 
                           n_1182);
   DATAPATH_I_IF_ID_IR_reg_22_inst : DFF_X1 port map( D => DATAPATH_I_N56, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_22_port, QN => 
                           n_1183);
   DATAPATH_I_IF_ID_IR_reg_23_inst : DFF_X1 port map( D => DATAPATH_I_N57, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_23_port, QN => 
                           n_1184);
   DATAPATH_I_IF_ID_IR_reg_24_inst : DFF_X1 port map( D => DATAPATH_I_N58, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_24_port, QN => 
                           n_1185);
   DATAPATH_I_IF_ID_IR_reg_25_inst : DFF_X1 port map( D => DATAPATH_I_N59, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_25_port, QN => 
                           n_1186);
   DATAPATH_I_IF_ID_IR_reg_26_inst : DFF_X1 port map( D => DATAPATH_I_N60, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_26_port, QN => 
                           n_1187);
   DATAPATH_I_IF_ID_IR_reg_27_inst : DFF_X1 port map( D => DATAPATH_I_N61, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_27_port, QN => n441
                           );
   DATAPATH_I_IF_ID_IR_reg_28_inst : DFF_X1 port map( D => DATAPATH_I_N62, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_28_port, QN => 
                           n_1188);
   DATAPATH_I_IF_ID_IR_reg_29_inst : DFF_X1 port map( D => DATAPATH_I_N63, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_29_port, QN => 
                           n_1189);
   DATAPATH_I_IF_ID_IR_reg_30_inst : DFF_X1 port map( D => DATAPATH_I_N64, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_30_port, QN => n440
                           );
   DATAPATH_I_IF_ID_IR_reg_31_inst : DFF_X1 port map( D => DATAPATH_I_N65, CK 
                           => CLK, Q => DATAPATH_I_IF_ID_IR_31_port, QN => 
                           n_1190);
   DATAPATH_I_ID_EX_RD_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N109, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_0_port, QN => 
                           n_1191);
   DATAPATH_I_EX_MEM_RD_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N308, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_0_port, QN => 
                           n_1192);
   DATAPATH_I_MEM_WB_RD_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N410, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_0_port, QN => 
                           n_1193);
   DATAPATH_I_ID_EX_RD_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N110, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_1_port, QN => 
                           n_1194);
   DATAPATH_I_EX_MEM_RD_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N309, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_1_port, QN => 
                           n_1195);
   DATAPATH_I_MEM_WB_RD_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N411, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_1_port, QN => 
                           n_1196);
   DATAPATH_I_ID_EX_RD_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N111, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_2_port, QN => 
                           n_1197);
   DATAPATH_I_EX_MEM_RD_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N310, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_2_port, QN => 
                           n_1198);
   DATAPATH_I_MEM_WB_RD_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N412, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_2_port, QN => 
                           n_1199);
   DATAPATH_I_ID_EX_RD_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N112, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_3_port, QN => 
                           n_1200);
   DATAPATH_I_EX_MEM_RD_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N311, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_3_port, QN => 
                           n_1201);
   DATAPATH_I_MEM_WB_RD_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N413, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_3_port, QN => 
                           n_1202);
   DATAPATH_I_ID_EX_RD_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N113, CK 
                           => CLK, Q => DATAPATH_I_ID_EX_RD_4_port, QN => 
                           n_1203);
   DATAPATH_I_EX_MEM_RD_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N312, CK 
                           => CLK, Q => DATAPATH_I_EX_MEM_RD_4_port, QN => 
                           n_1204);
   DATAPATH_I_MEM_WB_RD_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N414, CK 
                           => CLK, Q => DATAPATH_I_MEM_WB_RD_4_port, QN => 
                           n_1205);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_0_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N275, CK => CLK, Q => DATA_ADDR_0_port, 
                           QN => n_1206);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_1_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N276, CK => CLK, Q => DATA_ADDR_1_port, 
                           QN => n_1207);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_2_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N277, CK => CLK, Q => DATA_ADDR_2_port, 
                           QN => n_1208);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_3_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N278, CK => CLK, Q => DATA_ADDR_3_port, 
                           QN => n_1209);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_4_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N279, CK => CLK, Q => DATA_ADDR_4_port, 
                           QN => n_1210);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_5_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N280, CK => CLK, Q => DATA_ADDR_5_port, 
                           QN => n_1211);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_6_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N281, CK => CLK, Q => DATA_ADDR_6_port, 
                           QN => n_1212);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_7_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N282, CK => CLK, Q => DATA_ADDR_7_port, 
                           QN => n_1213);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_8_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N283, CK => CLK, Q => DATA_ADDR_8_port, 
                           QN => n_1214);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_9_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N284, CK => CLK, Q => DATA_ADDR_9_port, 
                           QN => n_1215);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_10_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N285, CK => CLK, Q => DATA_ADDR_10_port, 
                           QN => n_1216);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_11_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N286, CK => CLK, Q => DATA_ADDR_11_port, 
                           QN => n_1217);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_12_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N287, CK => CLK, Q => DATA_ADDR_12_port, 
                           QN => n_1218);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_13_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N288, CK => CLK, Q => DATA_ADDR_13_port, 
                           QN => n_1219);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_14_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N289, CK => CLK, Q => DATA_ADDR_14_port, 
                           QN => n_1220);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_15_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N290, CK => CLK, Q => DATA_ADDR_15_port, 
                           QN => n_1221);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_16_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N291, CK => CLK, Q => DATA_ADDR_16_port, 
                           QN => n_1222);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_17_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N292, CK => CLK, Q => DATA_ADDR_17_port, 
                           QN => n_1223);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_18_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N293, CK => CLK, Q => DATA_ADDR_18_port, 
                           QN => n_1224);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_19_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N294, CK => CLK, Q => DATA_ADDR_19_port, 
                           QN => n_1225);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_20_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N295, CK => CLK, Q => DATA_ADDR_20_port, 
                           QN => n_1226);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_21_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N296, CK => CLK, Q => DATA_ADDR_21_port, 
                           QN => n_1227);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_22_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N297, CK => CLK, Q => DATA_ADDR_22_port, 
                           QN => n_1228);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_23_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N298, CK => CLK, Q => DATA_ADDR_23_port, 
                           QN => n_1229);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_24_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N299, CK => CLK, Q => DATA_ADDR_24_port, 
                           QN => n_1230);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_25_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N300, CK => CLK, Q => DATA_ADDR_25_port, 
                           QN => n_1231);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_26_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N301, CK => CLK, Q => DATA_ADDR_26_port, 
                           QN => n_1232);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_27_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N302, CK => CLK, Q => DATA_ADDR_27_port, 
                           QN => n_1233);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_28_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N303, CK => CLK, Q => DATA_ADDR_28_port, 
                           QN => n_1234);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_29_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N304, CK => CLK, Q => DATA_ADDR_29_port, 
                           QN => n_1235);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_30_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N305, CK => CLK, Q => DATA_ADDR_30_port, 
                           QN => n_1236);
   DATAPATH_I_EX_MEM_ALU_OUTPUT_reg_31_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N306, CK => CLK, Q => DATA_ADDR_31_port, 
                           QN => n_1237);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_0_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N378, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_0_port, QN => n_1238);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_1_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N379, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_1_port, QN => n_1239);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_2_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N380, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_2_port, QN => n_1240);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_3_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N381, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_3_port, QN => n_1241);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_4_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N382, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_4_port, QN => n_1242);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_5_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N383, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_5_port, QN => n_1243);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_6_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N384, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_6_port, QN => n_1244);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_7_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N385, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_7_port, QN => n_1245);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_8_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N386, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_8_port, QN => n_1246);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_9_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N387, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_9_port, QN => n_1247);
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_10_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N388, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_10_port, QN => n_1248)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_11_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N389, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_11_port, QN => n_1249)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_12_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N390, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_12_port, QN => n_1250)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_13_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N391, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_13_port, QN => n_1251)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_14_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N392, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_14_port, QN => n_1252)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_15_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N393, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_15_port, QN => n_1253)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_16_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N394, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_16_port, QN => n_1254)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_17_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N395, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_17_port, QN => n_1255)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_18_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N396, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_18_port, QN => n_1256)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_19_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N397, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_19_port, QN => n_1257)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_20_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N398, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_20_port, QN => n_1258)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_21_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N399, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_21_port, QN => n_1259)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_22_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N400, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_22_port, QN => n_1260)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_23_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N401, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_23_port, QN => n_1261)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_24_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N402, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_24_port, QN => n_1262)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_25_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N403, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_25_port, QN => n_1263)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_26_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N404, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_26_port, QN => n_1264)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_27_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N405, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_27_port, QN => n_1265)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_28_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N406, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_28_port, QN => n_1266)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_29_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N407, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_29_port, QN => n_1267)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_30_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N408, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_30_port, QN => n_1268)
                           ;
   DATAPATH_I_MEM_WB_DRAM_OUTPUT_reg_31_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N409, CK => CLK, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_31_port, QN => n_1269)
                           ;
   DATAPATH_I_ID_EX_RF_OUT2_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N146,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_0_port, QN 
                           => n_1270);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N243
                           , CK => CLK, Q => DATA_IN_0_port, QN => n_1271);
   DATAPATH_I_ID_EX_RF_OUT2_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N147,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_1_port, QN 
                           => n_1272);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N244
                           , CK => CLK, Q => DATA_IN_1_port, QN => n_1273);
   DATAPATH_I_ID_EX_RF_OUT2_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N148,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_2_port, QN 
                           => n_1274);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N245
                           , CK => CLK, Q => DATA_IN_2_port, QN => n_1275);
   DATAPATH_I_ID_EX_RF_OUT2_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N149,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_3_port, QN 
                           => n_1276);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N246
                           , CK => CLK, Q => DATA_IN_3_port, QN => n_1277);
   DATAPATH_I_ID_EX_RF_OUT2_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N150,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_4_port, QN 
                           => n_1278);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N247
                           , CK => CLK, Q => DATA_IN_4_port, QN => n_1279);
   DATAPATH_I_ID_EX_RF_OUT2_reg_5_inst : DFF_X1 port map( D => DATAPATH_I_N151,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_5_port, QN 
                           => n_1280);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_5_inst : DFF_X1 port map( D => DATAPATH_I_N248
                           , CK => CLK, Q => DATA_IN_5_port, QN => n_1281);
   DATAPATH_I_ID_EX_RF_OUT2_reg_6_inst : DFF_X1 port map( D => DATAPATH_I_N152,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_6_port, QN 
                           => n_1282);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_6_inst : DFF_X1 port map( D => DATAPATH_I_N249
                           , CK => CLK, Q => DATA_IN_6_port, QN => n_1283);
   DATAPATH_I_ID_EX_RF_OUT2_reg_7_inst : DFF_X1 port map( D => DATAPATH_I_N153,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_7_port, QN 
                           => n_1284);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_7_inst : DFF_X1 port map( D => DATAPATH_I_N250
                           , CK => CLK, Q => DATA_IN_7_port, QN => n_1285);
   DATAPATH_I_ID_EX_RF_OUT2_reg_8_inst : DFF_X1 port map( D => DATAPATH_I_N154,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_8_port, QN 
                           => n_1286);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_8_inst : DFF_X1 port map( D => DATAPATH_I_N251
                           , CK => CLK, Q => DATA_IN_8_port, QN => n_1287);
   DATAPATH_I_ID_EX_RF_OUT2_reg_9_inst : DFF_X1 port map( D => DATAPATH_I_N155,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_9_port, QN 
                           => n_1288);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_9_inst : DFF_X1 port map( D => DATAPATH_I_N252
                           , CK => CLK, Q => DATA_IN_9_port, QN => n_1289);
   DATAPATH_I_ID_EX_RF_OUT2_reg_10_inst : DFF_X1 port map( D => DATAPATH_I_N156
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_10_port, 
                           QN => n_1290);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_10_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N253, CK => CLK, Q => DATA_IN_10_port, QN
                           => n_1291);
   DATAPATH_I_ID_EX_RF_OUT2_reg_11_inst : DFF_X1 port map( D => DATAPATH_I_N157
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_11_port, 
                           QN => n_1292);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_11_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N254, CK => CLK, Q => DATA_IN_11_port, QN
                           => n_1293);
   DATAPATH_I_ID_EX_RF_OUT2_reg_12_inst : DFF_X1 port map( D => DATAPATH_I_N158
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_12_port, 
                           QN => n_1294);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_12_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N255, CK => CLK, Q => DATA_IN_12_port, QN
                           => n_1295);
   DATAPATH_I_ID_EX_RF_OUT2_reg_13_inst : DFF_X1 port map( D => DATAPATH_I_N159
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_13_port, 
                           QN => n_1296);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_13_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N256, CK => CLK, Q => DATA_IN_13_port, QN
                           => n_1297);
   DATAPATH_I_ID_EX_RF_OUT2_reg_14_inst : DFF_X1 port map( D => DATAPATH_I_N160
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_14_port, 
                           QN => n_1298);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_14_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N257, CK => CLK, Q => DATA_IN_14_port, QN
                           => n_1299);
   DATAPATH_I_ID_EX_RF_OUT2_reg_15_inst : DFF_X1 port map( D => DATAPATH_I_N161
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_15_port, 
                           QN => n_1300);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_15_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N258, CK => CLK, Q => DATA_IN_15_port, QN
                           => n_1301);
   DATAPATH_I_ID_EX_RF_OUT2_reg_16_inst : DFF_X1 port map( D => DATAPATH_I_N162
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_16_port, 
                           QN => n_1302);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_16_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N259, CK => CLK, Q => DATA_IN_16_port, QN
                           => n_1303);
   DATAPATH_I_ID_EX_RF_OUT2_reg_17_inst : DFF_X1 port map( D => DATAPATH_I_N163
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_17_port, 
                           QN => n_1304);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_17_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N260, CK => CLK, Q => DATA_IN_17_port, QN
                           => n_1305);
   DATAPATH_I_ID_EX_RF_OUT2_reg_18_inst : DFF_X1 port map( D => DATAPATH_I_N164
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_18_port, 
                           QN => n_1306);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_18_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N261, CK => CLK, Q => DATA_IN_18_port, QN
                           => n_1307);
   DATAPATH_I_ID_EX_RF_OUT2_reg_19_inst : DFF_X1 port map( D => DATAPATH_I_N165
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_19_port, 
                           QN => n_1308);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_19_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N262, CK => CLK, Q => DATA_IN_19_port, QN
                           => n_1309);
   DATAPATH_I_ID_EX_RF_OUT2_reg_20_inst : DFF_X1 port map( D => DATAPATH_I_N166
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_20_port, 
                           QN => n_1310);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_20_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N263, CK => CLK, Q => DATA_IN_20_port, QN
                           => n_1311);
   DATAPATH_I_ID_EX_RF_OUT2_reg_21_inst : DFF_X1 port map( D => DATAPATH_I_N167
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_21_port, 
                           QN => n_1312);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_21_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N264, CK => CLK, Q => DATA_IN_21_port, QN
                           => n_1313);
   DATAPATH_I_ID_EX_RF_OUT2_reg_22_inst : DFF_X1 port map( D => DATAPATH_I_N168
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_22_port, 
                           QN => n_1314);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_22_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N265, CK => CLK, Q => DATA_IN_22_port, QN
                           => n_1315);
   DATAPATH_I_ID_EX_RF_OUT2_reg_23_inst : DFF_X1 port map( D => DATAPATH_I_N169
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_23_port, 
                           QN => n_1316);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_23_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N266, CK => CLK, Q => DATA_IN_23_port, QN
                           => n_1317);
   DATAPATH_I_ID_EX_RF_OUT2_reg_24_inst : DFF_X1 port map( D => DATAPATH_I_N170
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_24_port, 
                           QN => n_1318);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_24_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N267, CK => CLK, Q => DATA_IN_24_port, QN
                           => n_1319);
   DATAPATH_I_ID_EX_RF_OUT2_reg_25_inst : DFF_X1 port map( D => DATAPATH_I_N171
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_25_port, 
                           QN => n_1320);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_25_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N268, CK => CLK, Q => DATA_IN_25_port, QN
                           => n_1321);
   DATAPATH_I_ID_EX_RF_OUT2_reg_26_inst : DFF_X1 port map( D => DATAPATH_I_N172
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_26_port, 
                           QN => n_1322);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_26_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N269, CK => CLK, Q => DATA_IN_26_port, QN
                           => n_1323);
   DATAPATH_I_ID_EX_RF_OUT2_reg_27_inst : DFF_X1 port map( D => DATAPATH_I_N173
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_27_port, 
                           QN => n_1324);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_27_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N270, CK => CLK, Q => DATA_IN_27_port, QN
                           => n_1325);
   DATAPATH_I_ID_EX_RF_OUT2_reg_28_inst : DFF_X1 port map( D => DATAPATH_I_N174
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_28_port, 
                           QN => n_1326);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_28_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N271, CK => CLK, Q => DATA_IN_28_port, QN
                           => n_1327);
   DATAPATH_I_ID_EX_RF_OUT2_reg_29_inst : DFF_X1 port map( D => DATAPATH_I_N175
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_29_port, 
                           QN => n_1328);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_29_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N272, CK => CLK, Q => DATA_IN_29_port, QN
                           => n_1329);
   DATAPATH_I_ID_EX_RF_OUT2_reg_30_inst : DFF_X1 port map( D => DATAPATH_I_N176
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_30_port, 
                           QN => n_1330);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_30_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N273, CK => CLK, Q => DATA_IN_30_port, QN
                           => n_1331);
   DATAPATH_I_ID_EX_RF_OUT2_reg_31_inst : DFF_X1 port map( D => DATAPATH_I_N177
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT2_31_port, 
                           QN => n_1332);
   DATAPATH_I_EX_MEM_RF_OUT2_reg_31_inst : DFF_X1 port map( D => 
                           DATAPATH_I_N274, CK => CLK, Q => DATA_IN_31_port, QN
                           => n_1333);
   DATAPATH_I_ID_EX_RF_OUT1_reg_0_inst : DFF_X1 port map( D => DATAPATH_I_N114,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_0_port, QN 
                           => n_1334);
   DATAPATH_I_ID_EX_RF_OUT1_reg_1_inst : DFF_X1 port map( D => DATAPATH_I_N115,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_1_port, QN 
                           => n_1335);
   DATAPATH_I_ID_EX_RF_OUT1_reg_2_inst : DFF_X1 port map( D => DATAPATH_I_N116,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_2_port, QN 
                           => n_1336);
   DATAPATH_I_ID_EX_RF_OUT1_reg_3_inst : DFF_X1 port map( D => DATAPATH_I_N117,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_3_port, QN 
                           => n_1337);
   DATAPATH_I_ID_EX_RF_OUT1_reg_4_inst : DFF_X1 port map( D => DATAPATH_I_N118,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_4_port, QN 
                           => n_1338);
   DATAPATH_I_ID_EX_RF_OUT1_reg_5_inst : DFF_X1 port map( D => DATAPATH_I_N119,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_5_port, QN 
                           => n_1339);
   DATAPATH_I_ID_EX_RF_OUT1_reg_6_inst : DFF_X1 port map( D => DATAPATH_I_N120,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_6_port, QN 
                           => n_1340);
   DATAPATH_I_ID_EX_RF_OUT1_reg_7_inst : DFF_X1 port map( D => DATAPATH_I_N121,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_7_port, QN 
                           => n_1341);
   DATAPATH_I_ID_EX_RF_OUT1_reg_8_inst : DFF_X1 port map( D => DATAPATH_I_N122,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_8_port, QN 
                           => n_1342);
   DATAPATH_I_ID_EX_RF_OUT1_reg_9_inst : DFF_X1 port map( D => DATAPATH_I_N123,
                           CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_9_port, QN 
                           => n_1343);
   DATAPATH_I_ID_EX_RF_OUT1_reg_10_inst : DFF_X1 port map( D => DATAPATH_I_N124
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_10_port, 
                           QN => n_1344);
   DATAPATH_I_ID_EX_RF_OUT1_reg_11_inst : DFF_X1 port map( D => DATAPATH_I_N125
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_11_port, 
                           QN => n_1345);
   DATAPATH_I_ID_EX_RF_OUT1_reg_12_inst : DFF_X1 port map( D => DATAPATH_I_N126
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_12_port, 
                           QN => n_1346);
   DATAPATH_I_ID_EX_RF_OUT1_reg_13_inst : DFF_X1 port map( D => DATAPATH_I_N127
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_13_port, 
                           QN => n_1347);
   DATAPATH_I_ID_EX_RF_OUT1_reg_14_inst : DFF_X1 port map( D => DATAPATH_I_N128
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_14_port, 
                           QN => n_1348);
   DATAPATH_I_ID_EX_RF_OUT1_reg_15_inst : DFF_X1 port map( D => DATAPATH_I_N129
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_15_port, 
                           QN => n_1349);
   DATAPATH_I_ID_EX_RF_OUT1_reg_16_inst : DFF_X1 port map( D => DATAPATH_I_N130
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_16_port, 
                           QN => n_1350);
   DATAPATH_I_ID_EX_RF_OUT1_reg_17_inst : DFF_X1 port map( D => DATAPATH_I_N131
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_17_port, 
                           QN => n_1351);
   DATAPATH_I_ID_EX_RF_OUT1_reg_18_inst : DFF_X1 port map( D => DATAPATH_I_N132
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_18_port, 
                           QN => n_1352);
   DATAPATH_I_ID_EX_RF_OUT1_reg_19_inst : DFF_X1 port map( D => DATAPATH_I_N133
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_19_port, 
                           QN => n_1353);
   DATAPATH_I_ID_EX_RF_OUT1_reg_20_inst : DFF_X1 port map( D => DATAPATH_I_N134
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_20_port, 
                           QN => n_1354);
   DATAPATH_I_ID_EX_RF_OUT1_reg_21_inst : DFF_X1 port map( D => DATAPATH_I_N135
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_21_port, 
                           QN => n_1355);
   DATAPATH_I_ID_EX_RF_OUT1_reg_22_inst : DFF_X1 port map( D => DATAPATH_I_N136
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_22_port, 
                           QN => n_1356);
   DATAPATH_I_ID_EX_RF_OUT1_reg_23_inst : DFF_X1 port map( D => DATAPATH_I_N137
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_23_port, 
                           QN => n_1357);
   DATAPATH_I_ID_EX_RF_OUT1_reg_24_inst : DFF_X1 port map( D => DATAPATH_I_N138
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_24_port, 
                           QN => n_1358);
   DATAPATH_I_ID_EX_RF_OUT1_reg_25_inst : DFF_X1 port map( D => DATAPATH_I_N139
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_25_port, 
                           QN => n_1359);
   DATAPATH_I_ID_EX_RF_OUT1_reg_26_inst : DFF_X1 port map( D => DATAPATH_I_N140
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_26_port, 
                           QN => n_1360);
   DATAPATH_I_ID_EX_RF_OUT1_reg_27_inst : DFF_X1 port map( D => DATAPATH_I_N141
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_27_port, 
                           QN => n_1361);
   DATAPATH_I_ID_EX_RF_OUT1_reg_28_inst : DFF_X1 port map( D => DATAPATH_I_N142
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_28_port, 
                           QN => n_1362);
   DATAPATH_I_ID_EX_RF_OUT1_reg_29_inst : DFF_X1 port map( D => DATAPATH_I_N143
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_29_port, 
                           QN => n_1363);
   DATAPATH_I_ID_EX_RF_OUT1_reg_30_inst : DFF_X1 port map( D => DATAPATH_I_N144
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_30_port, 
                           QN => n_1364);
   DATAPATH_I_ID_EX_RF_OUT1_reg_31_inst : DFF_X1 port map( D => DATAPATH_I_N145
                           , CK => CLK, Q => DATAPATH_I_ID_EX_RF_OUT1_31_port, 
                           QN => n_1365);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_N3, GN => RST,
                           Q => IR_0_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_N3, GN => RST,
                           Q => IR_1_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_N3, GN => RST,
                           Q => IR_2_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_N3, GN => RST,
                           Q => IR_3_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_N3, GN => RST,
                           Q => IR_4_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_N3, GN => RST,
                           Q => IR_5_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_N3, GN => RST,
                           Q => IR_6_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_N3, GN => RST,
                           Q => IR_7_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_N3, GN => RST,
                           Q => IR_8_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_N3, GN => RST,
                           Q => IR_9_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_N3, GN => RST
                           , Q => IR_10_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_N3, GN => RST
                           , Q => DATAPATH_I_n29);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_N3, GN => RST
                           , Q => DATAPATH_I_n28);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_N3, GN => RST
                           , Q => DATAPATH_I_n27);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_N3, GN => RST
                           , Q => DATAPATH_I_n26);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_N3, GN => RST
                           , Q => DATAPATH_I_n25);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_N3, GN => RST
                           , Q => DATAPATH_I_n24);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_N3, GN => RST
                           , Q => DATAPATH_I_n23);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_N3, GN => RST
                           , Q => DATAPATH_I_n22);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_N3, GN => RST
                           , Q => DATAPATH_I_n21);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_N3, GN => RST
                           , Q => DATAPATH_I_n20);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_N3, GN => RST
                           , Q => DATAPATH_I_n19);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_N3, GN => RST
                           , Q => DATAPATH_I_n18);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_N3, GN => RST
                           , Q => DATAPATH_I_n17);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_N3, GN => RST
                           , Q => DATAPATH_I_n16);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_N3, GN => RST
                           , Q => DATAPATH_I_n15);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_N3, GN => RST
                           , Q => IR_26_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_N3, GN => RST
                           , Q => IR_27_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_N3, GN => RST
                           , Q => IR_28_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_N3, GN => RST
                           , Q => IR_29_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_N3, GN => RST
                           , Q => IR_30_port);
   DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_N3, GN => RST
                           , Q => IR_31_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_0_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_0_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_1_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_1_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_2_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_2_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_3_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_3_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_4_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_4_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_5_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_5_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_6_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_6_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_7_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_7_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_8_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_8_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_9_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_9_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_10_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_10_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_11_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_11_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_12_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_12_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_13_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_13_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_14_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_14_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_15_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_15_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_16_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_16_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_17_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_17_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_18_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_18_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_19_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_19_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_20_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_20_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_21_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_21_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_22_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_22_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_23_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_23_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_24_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_24_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_25_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_25_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_26_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_26_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_27_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_27_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_28_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_28_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_29_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_29_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_30_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_30_port);
   DATAPATH_I_LATCH_ALUOUT_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_ALUOUT_LDI_31_N3, GN => RST, Q => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_31_port);
   DATAPATH_I_LATCH_LMD_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_0_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_0_port);
   DATAPATH_I_LATCH_LMD_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_1_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_1_port);
   DATAPATH_I_LATCH_LMD_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_2_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_2_port);
   DATAPATH_I_LATCH_LMD_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_3_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_3_port);
   DATAPATH_I_LATCH_LMD_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_4_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_4_port);
   DATAPATH_I_LATCH_LMD_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_5_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_5_port);
   DATAPATH_I_LATCH_LMD_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_6_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_6_port);
   DATAPATH_I_LATCH_LMD_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_7_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_7_port);
   DATAPATH_I_LATCH_LMD_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_8_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_8_port);
   DATAPATH_I_LATCH_LMD_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_9_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_9_port);
   DATAPATH_I_LATCH_LMD_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_10_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_10_port);
   DATAPATH_I_LATCH_LMD_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_11_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_11_port);
   DATAPATH_I_LATCH_LMD_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_12_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_12_port);
   DATAPATH_I_LATCH_LMD_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_13_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_13_port);
   DATAPATH_I_LATCH_LMD_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_14_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_14_port);
   DATAPATH_I_LATCH_LMD_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_15_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_15_port);
   DATAPATH_I_LATCH_LMD_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_16_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_16_port);
   DATAPATH_I_LATCH_LMD_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_17_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_17_port);
   DATAPATH_I_LATCH_LMD_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_18_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_18_port);
   DATAPATH_I_LATCH_LMD_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_19_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_19_port);
   DATAPATH_I_LATCH_LMD_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_20_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_20_port);
   DATAPATH_I_LATCH_LMD_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_21_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_21_port);
   DATAPATH_I_LATCH_LMD_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_22_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_22_port);
   DATAPATH_I_LATCH_LMD_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_23_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_23_port);
   DATAPATH_I_LATCH_LMD_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_24_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_24_port);
   DATAPATH_I_LATCH_LMD_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_25_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_25_port);
   DATAPATH_I_LATCH_LMD_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_26_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_26_port);
   DATAPATH_I_LATCH_LMD_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_27_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_27_port);
   DATAPATH_I_LATCH_LMD_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_28_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_28_port);
   DATAPATH_I_LATCH_LMD_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_29_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_29_port);
   DATAPATH_I_LATCH_LMD_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_30_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_30_port);
   DATAPATH_I_LATCH_LMD_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_LMD_LDI_31_N3, GN => RST, Q => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_31_port);
   DATAPATH_I_LATCH_RF2_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_0_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_0_port);
   DATAPATH_I_LATCH_RF2_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_1_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_1_port);
   DATAPATH_I_LATCH_RF2_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_2_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_2_port);
   DATAPATH_I_LATCH_RF2_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_3_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_3_port);
   DATAPATH_I_LATCH_RF2_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_4_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_4_port);
   DATAPATH_I_LATCH_RF2_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_5_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_5_port);
   DATAPATH_I_LATCH_RF2_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_6_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_6_port);
   DATAPATH_I_LATCH_RF2_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_7_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_7_port);
   DATAPATH_I_LATCH_RF2_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_8_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_8_port);
   DATAPATH_I_LATCH_RF2_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_9_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_9_port);
   DATAPATH_I_LATCH_RF2_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_10_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_10_port);
   DATAPATH_I_LATCH_RF2_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_11_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_11_port);
   DATAPATH_I_LATCH_RF2_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_12_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_12_port);
   DATAPATH_I_LATCH_RF2_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_13_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_13_port);
   DATAPATH_I_LATCH_RF2_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_14_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_14_port);
   DATAPATH_I_LATCH_RF2_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_15_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_15_port);
   DATAPATH_I_LATCH_RF2_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_16_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_16_port);
   DATAPATH_I_LATCH_RF2_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_17_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_17_port);
   DATAPATH_I_LATCH_RF2_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_18_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_18_port);
   DATAPATH_I_LATCH_RF2_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_19_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_19_port);
   DATAPATH_I_LATCH_RF2_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_20_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_20_port);
   DATAPATH_I_LATCH_RF2_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_21_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_21_port);
   DATAPATH_I_LATCH_RF2_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_22_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_22_port);
   DATAPATH_I_LATCH_RF2_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_23_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_23_port);
   DATAPATH_I_LATCH_RF2_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_24_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_24_port);
   DATAPATH_I_LATCH_RF2_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_25_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_25_port);
   DATAPATH_I_LATCH_RF2_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_26_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_26_port);
   DATAPATH_I_LATCH_RF2_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_27_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_27_port);
   DATAPATH_I_LATCH_RF2_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_28_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_28_port);
   DATAPATH_I_LATCH_RF2_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_29_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_29_port);
   DATAPATH_I_LATCH_RF2_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_30_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_30_port);
   DATAPATH_I_LATCH_RF2_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF2_LDI_31_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_31_port);
   DATAPATH_I_LATCH_RF1_LDI_0_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_0_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_0_port);
   DATAPATH_I_LATCH_RF1_LDI_1_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_1_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_1_port);
   DATAPATH_I_LATCH_RF1_LDI_2_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_2_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_2_port);
   DATAPATH_I_LATCH_RF1_LDI_3_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_3_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_3_port);
   DATAPATH_I_LATCH_RF1_LDI_4_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_4_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_4_port);
   DATAPATH_I_LATCH_RF1_LDI_5_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_5_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_5_port);
   DATAPATH_I_LATCH_RF1_LDI_6_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_6_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_6_port);
   DATAPATH_I_LATCH_RF1_LDI_7_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_7_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_7_port);
   DATAPATH_I_LATCH_RF1_LDI_8_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_8_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_8_port);
   DATAPATH_I_LATCH_RF1_LDI_9_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_9_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_9_port);
   DATAPATH_I_LATCH_RF1_LDI_10_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_10_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_10_port);
   DATAPATH_I_LATCH_RF1_LDI_11_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_11_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_11_port);
   DATAPATH_I_LATCH_RF1_LDI_12_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_12_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_12_port);
   DATAPATH_I_LATCH_RF1_LDI_13_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_13_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_13_port);
   DATAPATH_I_LATCH_RF1_LDI_14_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_14_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_14_port);
   DATAPATH_I_LATCH_RF1_LDI_15_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_15_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_15_port);
   DATAPATH_I_LATCH_RF1_LDI_16_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_16_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_16_port);
   DATAPATH_I_LATCH_RF1_LDI_17_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_17_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_17_port);
   DATAPATH_I_LATCH_RF1_LDI_18_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_18_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_18_port);
   DATAPATH_I_LATCH_RF1_LDI_19_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_19_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_19_port);
   DATAPATH_I_LATCH_RF1_LDI_20_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_20_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_20_port);
   DATAPATH_I_LATCH_RF1_LDI_21_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_21_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_21_port);
   DATAPATH_I_LATCH_RF1_LDI_22_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_22_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_22_port);
   DATAPATH_I_LATCH_RF1_LDI_23_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_23_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_23_port);
   DATAPATH_I_LATCH_RF1_LDI_24_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_24_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_24_port);
   DATAPATH_I_LATCH_RF1_LDI_25_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_25_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_25_port);
   DATAPATH_I_LATCH_RF1_LDI_26_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_26_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_26_port);
   DATAPATH_I_LATCH_RF1_LDI_27_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_27_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_27_port);
   DATAPATH_I_LATCH_RF1_LDI_28_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_28_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_28_port);
   DATAPATH_I_LATCH_RF1_LDI_29_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_29_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_29_port);
   DATAPATH_I_LATCH_RF1_LDI_30_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_30_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_30_port);
   DATAPATH_I_LATCH_RF1_LDI_31_Q_reg : DLL_X1 port map( D => 
                           DATAPATH_I_LATCH_RF1_LDI_31_N3, GN => RST, Q => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_31_port);
   CU_I_aluOpcode2_reg_0_inst : DFFR_X1 port map( D => CU_I_aluOpcode1_0_port, 
                           CK => CLK, RN => RST, Q => CU_I_aluOpcode2_0_port, 
                           QN => n_1366);
   CU_I_aluOpcode3_reg_0_inst : DFFR_X1 port map( D => CU_I_aluOpcode2_0_port, 
                           CK => CLK, RN => RST, Q => ALU_OPCODE_i_6_port, QN 
                           => n_1367);
   CU_I_aluOpcode2_reg_3_inst : DFFR_X1 port map( D => CU_I_aluOpcode1_3_port, 
                           CK => CLK, RN => RST, Q => CU_I_aluOpcode2_3_port, 
                           QN => n_1368);
   CU_I_aluOpcode3_reg_3_inst : DFFR_X1 port map( D => CU_I_aluOpcode2_3_port, 
                           CK => CLK, RN => RST, Q => ALU_OPCODE_i_3_port, QN 
                           => n_1369);
   CU_I_aluOpcode2_reg_4_inst : DFFR_X1 port map( D => CU_I_aluOpcode1_4_port, 
                           CK => CLK, RN => RST, Q => CU_I_aluOpcode2_4_port, 
                           QN => n_1370);
   CU_I_aluOpcode3_reg_4_inst : DFFR_X1 port map( D => CU_I_aluOpcode2_4_port, 
                           CK => CLK, RN => RST, Q => ALU_OPCODE_i_2_port, QN 
                           => n_1371);
   CU_I_aluOpcode2_reg_2_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_2_port, 
                           CK => CLK, SN => RST, Q => CU_I_aluOpcode2_2_port, 
                           QN => n_1372);
   CU_I_aluOpcode3_reg_2_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_2_port, 
                           CK => CLK, SN => RST, Q => ALU_OPCODE_i_4_port, QN 
                           => n_1373);
   CU_I_aluOpcode2_reg_1_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_1_port, 
                           CK => CLK, SN => RST, Q => CU_I_aluOpcode2_1_port, 
                           QN => n_1374);
   CU_I_aluOpcode3_reg_1_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_1_port, 
                           CK => CLK, SN => RST, Q => ALU_OPCODE_i_5_port, QN 
                           => n_1375);
   CU_I_aluOpcode2_reg_5_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_5_port, 
                           CK => CLK, SN => RST, Q => CU_I_aluOpcode2_5_port, 
                           QN => n_1376);
   CU_I_aluOpcode3_reg_5_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_5_port, 
                           CK => CLK, SN => RST, Q => ALU_OPCODE_i_1_port, QN 
                           => n_1377);
   CU_I_aluOpcode2_reg_6_inst : DFFS_X1 port map( D => CU_I_aluOpcode1_6_port, 
                           CK => CLK, SN => RST, Q => CU_I_aluOpcode2_6_port, 
                           QN => n_1378);
   CU_I_aluOpcode3_reg_6_inst : DFFS_X1 port map( D => CU_I_aluOpcode2_6_port, 
                           CK => CLK, SN => RST, Q => ALU_OPCODE_i_0_port, QN 
                           => n_1379);
   U751 : INV_X1 port map( A => RST, ZN => n317);
   U752 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_1_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_1_N3);
   U753 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_29_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_29_N3);
   U754 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_3_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_3_N3);
   U755 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_28_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_28_N3);
   U756 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_27_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_27_N3);
   U757 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_0_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_0_N3);
   U758 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_31_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_31_N3);
   U759 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_30_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_30_N3);
   U760 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_24_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_24_N3);
   U761 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_23_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_23_N3);
   U762 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_2_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_2_N3);
   U763 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_22_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_22_N3);
   U764 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_26_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_26_N3);
   U765 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_21_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_21_N3);
   U766 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_25_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_25_N3);
   U767 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_20_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_20_N3);
   U768 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_19_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_19_N3);
   U769 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_18_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_18_N3);
   U770 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_17_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_17_N3);
   U771 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_16_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_16_N3);
   U772 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_15_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_15_N3);
   U773 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_14_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_14_N3);
   U774 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_13_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_13_N3);
   U775 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_12_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_12_N3);
   U776 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_11_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_11_N3);
   U777 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_10_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_10_N3);
   U778 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_9_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_9_N3);
   U779 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_8_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_8_N3);
   U780 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_7_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_7_N3);
   U781 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_6_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_6_N3);
   U782 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_5_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_5_N3);
   U783 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_4_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_4_N3);
   U784 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_3_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_3_N3);
   U785 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_2_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_2_N3);
   U786 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_1_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_1_N3);
   U787 : AND2_X1 port map( A1 => RST, A2 => IR_BUS_0_port, ZN => 
                           DATAPATH_I_INSTRUCTION_REGISTER_LDI_0_N3);
   U788 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_4_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_4_N3);
   U789 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_26_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_26_N3);
   U790 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_27_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_27_N3);
   U791 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_28_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_28_N3);
   U792 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_29_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_29_N3);
   U793 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_30_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_30_N3);
   U794 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_31_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_31_N3);
   U795 : INV_X1 port map( A => IR_28_port, ZN => n407);
   U796 : NOR2_X1 port map( A1 => n317, A2 => n407, ZN => DATAPATH_I_N62);
   U797 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_25_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_25_N3);
   U798 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_6_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_6_N3);
   U799 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_7_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_7_N3);
   U800 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_8_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_8_N3);
   U801 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_9_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_9_N3);
   U802 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_10_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_10_N3);
   U803 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_11_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_11_N3);
   U804 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_12_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_12_N3);
   U805 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_13_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_13_N3);
   U806 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_14_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_14_N3);
   U807 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_15_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_15_N3);
   U808 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_16_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_16_N3);
   U809 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_17_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_17_N3);
   U810 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_18_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_18_N3);
   U811 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_19_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_19_N3);
   U812 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_20_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_20_N3);
   U813 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_21_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_21_N3);
   U814 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_22_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_22_N3);
   U815 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_23_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_23_N3);
   U816 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_24_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_24_N3);
   U817 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_25_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_25_N3);
   U818 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_26_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_26_N3);
   U819 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_27_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_27_N3);
   U820 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_28_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_28_N3);
   U821 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_29_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_29_N3);
   U822 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_30_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_30_N3);
   U823 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_31_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_31_N3);
   U824 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_0_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_0_N3);
   U825 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_1_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_1_N3);
   U826 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_2_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_2_N3);
   U827 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_3_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_3_N3);
   U828 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_4_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_4_N3);
   U829 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_5_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_5_N3);
   U830 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_6_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_6_N3);
   U831 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_7_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_7_N3);
   U832 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_8_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_8_N3);
   U833 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_9_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_9_N3);
   U834 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_10_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_10_N3);
   U835 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_11_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_11_N3);
   U836 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_12_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_12_N3);
   U837 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_13_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_13_N3);
   U838 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_14_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_14_N3);
   U839 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_15_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_15_N3);
   U840 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_16_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_16_N3);
   U841 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_17_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_17_N3);
   U842 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_18_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_18_N3);
   U843 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_19_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_19_N3);
   U844 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_20_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_20_N3);
   U845 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_21_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_21_N3);
   U846 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_22_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_22_N3);
   U847 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_23_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_23_N3);
   U848 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_24_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_24_N3);
   U849 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_25_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_25_N3);
   U850 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_26_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_26_N3);
   U851 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_27_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_27_N3);
   U852 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_28_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_28_N3);
   U853 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_29_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_29_N3);
   U854 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_30_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_30_N3);
   U855 : AND2_X1 port map( A1 => RST, A2 => DATA_OUT_31_port, ZN => 
                           DATAPATH_I_LATCH_LMD_LDI_31_N3);
   U856 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ALU_OUTPUT_5_port, ZN 
                           => DATAPATH_I_LATCH_ALUOUT_LDI_5_N3);
   U857 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_0_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_0_N3);
   U858 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_1_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_1_N3);
   U859 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_2_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_2_N3);
   U860 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_3_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_3_N3);
   U861 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_4_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_4_N3);
   U862 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_5_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_5_N3);
   U863 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_6_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_6_N3);
   U864 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_7_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_7_N3);
   U865 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_8_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_8_N3);
   U866 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_9_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_9_N3);
   U867 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_10_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_10_N3);
   U868 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_11_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_11_N3);
   U869 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_12_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_12_N3);
   U870 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_13_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_13_N3);
   U871 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_14_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_14_N3);
   U872 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_15_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_15_N3);
   U873 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_16_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_16_N3);
   U874 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_17_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_17_N3);
   U875 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_18_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_18_N3);
   U876 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_19_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_19_N3);
   U877 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_20_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_20_N3);
   U878 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_21_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_21_N3);
   U879 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_22_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_22_N3);
   U880 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_23_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_23_N3);
   U881 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_24_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_24_N3);
   U882 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_25_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_25_N3);
   U883 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_26_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_26_N3);
   U884 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_27_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_27_N3);
   U885 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_28_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_28_N3);
   U886 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_29_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_29_N3);
   U887 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_30_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_30_N3);
   U888 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT2_31_port, ZN => 
                           DATAPATH_I_LATCH_RF2_LDI_31_N3);
   U889 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_0_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_0_N3);
   U890 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_1_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_1_N3);
   U891 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_2_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_2_N3);
   U892 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_3_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_3_N3);
   U893 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_4_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_4_N3);
   U894 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_5_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_5_N3);
   U895 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_6_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_6_N3);
   U896 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_7_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_7_N3);
   U897 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_8_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_8_N3);
   U898 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_9_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_9_N3);
   U899 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_10_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_10_N3);
   U900 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_11_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_11_N3);
   U901 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_12_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_12_N3);
   U902 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_13_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_13_N3);
   U903 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_14_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_14_N3);
   U904 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_15_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_15_N3);
   U905 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_16_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_16_N3);
   U906 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_17_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_17_N3);
   U907 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_18_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_18_N3);
   U908 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_19_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_19_N3);
   U909 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_20_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_20_N3);
   U910 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_21_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_21_N3);
   U911 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_22_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_22_N3);
   U912 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_23_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_23_N3);
   U913 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_RF_OUT1_24_port, ZN => 
                           DATAPATH_I_LATCH_RF1_LDI_24_N3);
   U914 : NOR2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_28_port, A2 => 
                           DATAPATH_I_IF_ID_IR_30_port, ZN => n321);
   U915 : AND4_X1 port map( A1 => DATAPATH_I_IF_ID_IR_29_port, A2 => 
                           DATAPATH_I_IF_ID_IR_31_port, A3 => 
                           DATAPATH_I_IF_ID_IR_27_port, A4 => 
                           DATAPATH_I_IF_ID_IR_26_port, ZN => n320);
   U916 : OR3_X1 port map( A1 => DATAPATH_I_IF_ID_IR_28_port, A2 => 
                           DATAPATH_I_IF_ID_IR_29_port, A3 => 
                           DATAPATH_I_IF_ID_IR_31_port, ZN => n318);
   U917 : OR4_X1 port map( A1 => DATAPATH_I_IF_ID_IR_26_port, A2 => 
                           DATAPATH_I_IF_ID_IR_27_port, A3 => 
                           DATAPATH_I_IF_ID_IR_30_port, A4 => n318, ZN => n346)
                           ;
   U918 : INV_X1 port map( A => n346, ZN => n319);
   U919 : AOI21_X1 port map( B1 => n321, B2 => n320, A => n319, ZN => n322);
   U920 : INV_X1 port map( A => n322, ZN => n345);
   U921 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_20_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_4_port);
   U922 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_18_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_2_port);
   U923 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_17_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_1_port);
   U924 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_16_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_0_port);
   U925 : NOR4_X1 port map( A1 => DATAPATH_I_IF_ID_IR_28_port, A2 => 
                           DATAPATH_I_IF_ID_IR_29_port, A3 => 
                           DATAPATH_I_IF_ID_IR_31_port, A4 => n441, ZN => n347)
                           ;
   U926 : NAND2_X1 port map( A1 => n347, A2 => n440, ZN => n323);
   U927 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_25_port, A2 => n323, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_4_port);
   U928 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_23_port, A2 => n323, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_2_port);
   U929 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_22_port, A2 => n323, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_1_port);
   U930 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_21_port, A2 => n323, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_0_port);
   U931 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_0_port, ZN => 
                           DATAPATH_I_N308);
   U932 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_0_port, ZN =>
                           DATAPATH_I_N410);
   U933 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_1_port, ZN => 
                           DATAPATH_I_N309);
   U934 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_1_port, ZN =>
                           DATAPATH_I_N411);
   U935 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_2_port, ZN => 
                           DATAPATH_I_N310);
   U936 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_2_port, ZN =>
                           DATAPATH_I_N412);
   U937 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_3_port, ZN => 
                           DATAPATH_I_N311);
   U938 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_3_port, ZN =>
                           DATAPATH_I_N413);
   U939 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RD_4_port, ZN => 
                           DATAPATH_I_N312);
   U940 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_EX_MEM_RD_4_port, ZN =>
                           DATAPATH_I_N414);
   U941 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_23_port, ZN => 
                           DATAPATH_I_N169);
   U942 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_14_port, ZN => 
                           DATAPATH_I_N160);
   U943 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_21_port, ZN => 
                           DATAPATH_I_N135);
   U944 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_17_port, ZN => 
                           DATAPATH_I_N163);
   U945 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_13_port, ZN => 
                           DATAPATH_I_N159);
   U946 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_19_port, ZN => 
                           DATAPATH_I_N165);
   U947 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_15_port, ZN => 
                           DATAPATH_I_N161);
   U948 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_20_port, ZN => 
                           DATAPATH_I_N166);
   U949 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_16_port, ZN => 
                           DATAPATH_I_N162);
   U950 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_24_port, ZN => 
                           DATAPATH_I_N170);
   U951 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_22_port, ZN => 
                           DATAPATH_I_N168);
   U952 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_25_port, ZN => 
                           DATAPATH_I_N171);
   U953 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_18_port, ZN => 
                           DATAPATH_I_N164);
   U954 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_26_port, ZN => 
                           DATAPATH_I_N172);
   U955 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_27_port, ZN => 
                           DATAPATH_I_N173);
   U956 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_21_port, ZN => 
                           DATAPATH_I_N167);
   U957 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_28_port, ZN => 
                           DATAPATH_I_N174);
   U958 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_29_port, ZN => 
                           DATAPATH_I_N175);
   U959 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_30_port, ZN => 
                           DATAPATH_I_N176);
   U960 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_31_port, ZN => 
                           DATAPATH_I_N177);
   U961 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_0_port, ZN => 
                           DATAPATH_I_N114);
   U962 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_1_port, ZN => 
                           DATAPATH_I_N115);
   U963 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_2_port, ZN => 
                           DATAPATH_I_N116);
   U964 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_3_port, ZN => 
                           DATAPATH_I_N117);
   U965 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_4_port, ZN => 
                           DATAPATH_I_N118);
   U966 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_5_port, ZN => 
                           DATAPATH_I_N119);
   U967 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_6_port, ZN => 
                           DATAPATH_I_N120);
   U968 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_7_port, ZN => 
                           DATAPATH_I_N121);
   U969 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_8_port, ZN => 
                           DATAPATH_I_N122);
   U970 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_12_port, ZN => 
                           DATAPATH_I_N158);
   U971 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_9_port, ZN => 
                           DATAPATH_I_N123);
   U972 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_10_port, ZN => 
                           DATAPATH_I_N124);
   U973 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_11_port, ZN => 
                           DATAPATH_I_N125);
   U974 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_31_port, ZN => 
                           DATAPATH_I_N145);
   U975 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_12_port, ZN => 
                           DATAPATH_I_N126);
   U976 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_30_port, ZN => 
                           DATAPATH_I_N144);
   U977 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_29_port, ZN => 
                           DATAPATH_I_N143);
   U978 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_28_port, ZN => 
                           DATAPATH_I_N142);
   U979 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_13_port, ZN => 
                           DATAPATH_I_N127);
   U980 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_14_port, ZN => 
                           DATAPATH_I_N128);
   U981 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_27_port, ZN => 
                           DATAPATH_I_N141);
   U982 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_26_port, ZN => 
                           DATAPATH_I_N140);
   U983 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_15_port, ZN => 
                           DATAPATH_I_N129);
   U984 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_25_port, ZN => 
                           DATAPATH_I_N139);
   U985 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_16_port, ZN => 
                           DATAPATH_I_N130);
   U986 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_17_port, ZN => 
                           DATAPATH_I_N131);
   U987 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_24_port, ZN => 
                           DATAPATH_I_N138);
   U988 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_18_port, ZN => 
                           DATAPATH_I_N132);
   U989 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_23_port, ZN => 
                           DATAPATH_I_N137);
   U990 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_19_port, ZN => 
                           DATAPATH_I_N133);
   U991 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_22_port, ZN => 
                           DATAPATH_I_N136);
   U992 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT1_NEXT_20_port, ZN => 
                           DATAPATH_I_N134);
   U993 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n28, ZN => 
                           DATAPATH_I_N46);
   U994 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n27, ZN => 
                           DATAPATH_I_N47);
   U995 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n26, ZN => 
                           DATAPATH_I_N48);
   U996 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n25, ZN => 
                           DATAPATH_I_N49);
   U997 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n24, ZN => 
                           DATAPATH_I_N50);
   U998 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n23, ZN => 
                           DATAPATH_I_N51);
   U999 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n22, ZN => 
                           DATAPATH_I_N52);
   U1000 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n21, ZN => 
                           DATAPATH_I_N53);
   U1001 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n20, ZN => 
                           DATAPATH_I_N54);
   U1002 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n19, ZN => 
                           DATAPATH_I_N55);
   U1003 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n18, ZN => 
                           DATAPATH_I_N56);
   U1004 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n17, ZN => 
                           DATAPATH_I_N57);
   U1005 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n16, ZN => 
                           DATAPATH_I_N58);
   U1006 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n15, ZN => 
                           DATAPATH_I_N59);
   U1007 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_0_port, ZN => 
                           DATAPATH_I_N275);
   U1008 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_1_port, ZN => 
                           DATAPATH_I_N276);
   U1009 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_2_port, ZN => 
                           DATAPATH_I_N277);
   U1010 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_3_port, ZN => 
                           DATAPATH_I_N278);
   U1011 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_4_port, ZN => 
                           DATAPATH_I_N279);
   U1012 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_5_port, ZN => 
                           DATAPATH_I_N280);
   U1013 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_6_port, ZN => 
                           DATAPATH_I_N281);
   U1014 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_7_port, ZN => 
                           DATAPATH_I_N282);
   U1015 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_8_port, ZN => 
                           DATAPATH_I_N283);
   U1016 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_9_port, ZN => 
                           DATAPATH_I_N284);
   U1017 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_10_port, ZN => 
                           DATAPATH_I_N285);
   U1018 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_11_port, ZN => 
                           DATAPATH_I_N286);
   U1019 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_12_port, ZN => 
                           DATAPATH_I_N287);
   U1020 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_13_port, ZN => 
                           DATAPATH_I_N288);
   U1021 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_14_port, ZN => 
                           DATAPATH_I_N289);
   U1022 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_15_port, ZN => 
                           DATAPATH_I_N290);
   U1023 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_16_port, ZN => 
                           DATAPATH_I_N291);
   U1024 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_17_port, ZN => 
                           DATAPATH_I_N292);
   U1025 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_18_port, ZN => 
                           DATAPATH_I_N293);
   U1026 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_19_port, ZN => 
                           DATAPATH_I_N294);
   U1027 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_20_port, ZN => 
                           DATAPATH_I_N295);
   U1028 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_21_port, ZN => 
                           DATAPATH_I_N296);
   U1029 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_22_port, ZN => 
                           DATAPATH_I_N297);
   U1030 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_23_port, ZN => 
                           DATAPATH_I_N298);
   U1031 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_24_port, ZN => 
                           DATAPATH_I_N299);
   U1032 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_25_port, ZN => 
                           DATAPATH_I_N300);
   U1033 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_26_port, ZN => 
                           DATAPATH_I_N301);
   U1034 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_n29, ZN => 
                           DATAPATH_I_N45);
   U1035 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_27_port, ZN => 
                           DATAPATH_I_N302);
   U1036 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_28_port, ZN => 
                           DATAPATH_I_N303);
   U1037 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_29_port, ZN => 
                           DATAPATH_I_N304);
   U1038 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_30_port, ZN => 
                           DATAPATH_I_N305);
   U1039 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_EX_MEM_ALU_OUTPUT_NEXT_31_port, ZN => 
                           DATAPATH_I_N306);
   U1040 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_0_port, ZN => 
                           DATAPATH_I_N378);
   U1041 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_1_port, ZN => 
                           DATAPATH_I_N379);
   U1042 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_2_port, ZN => 
                           DATAPATH_I_N380);
   U1043 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_3_port, ZN => 
                           DATAPATH_I_N381);
   U1044 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_4_port, ZN => 
                           DATAPATH_I_N382);
   U1045 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_5_port, ZN => 
                           DATAPATH_I_N383);
   U1046 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_6_port, ZN => 
                           DATAPATH_I_N384);
   U1047 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_7_port, ZN => 
                           DATAPATH_I_N385);
   U1048 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_8_port, ZN => 
                           DATAPATH_I_N386);
   U1049 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_9_port, ZN => 
                           DATAPATH_I_N387);
   U1050 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_10_port, ZN => 
                           DATAPATH_I_N388);
   U1051 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_11_port, ZN => 
                           DATAPATH_I_N389);
   U1052 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_12_port, ZN => 
                           DATAPATH_I_N390);
   U1053 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_13_port, ZN => 
                           DATAPATH_I_N391);
   U1054 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_14_port, ZN => 
                           DATAPATH_I_N392);
   U1055 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_15_port, ZN => 
                           DATAPATH_I_N393);
   U1056 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_16_port, ZN => 
                           DATAPATH_I_N394);
   U1057 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_17_port, ZN => 
                           DATAPATH_I_N395);
   U1058 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_18_port, ZN => 
                           DATAPATH_I_N396);
   U1059 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_19_port, ZN => 
                           DATAPATH_I_N397);
   U1060 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_20_port, ZN => 
                           DATAPATH_I_N398);
   U1061 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_21_port, ZN => 
                           DATAPATH_I_N399);
   U1062 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_22_port, ZN => 
                           DATAPATH_I_N400);
   U1063 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_23_port, ZN => 
                           DATAPATH_I_N401);
   U1064 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_24_port, ZN => 
                           DATAPATH_I_N402);
   U1065 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_25_port, ZN => 
                           DATAPATH_I_N403);
   U1066 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_26_port, ZN => 
                           DATAPATH_I_N404);
   U1067 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_27_port, ZN => 
                           DATAPATH_I_N405);
   U1068 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_28_port, ZN => 
                           DATAPATH_I_N406);
   U1069 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_29_port, ZN => 
                           DATAPATH_I_N407);
   U1070 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_30_port, ZN => 
                           DATAPATH_I_N408);
   U1071 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_MEM_WB_DRAM_OUTPUT_NEXT_31_port, ZN => 
                           DATAPATH_I_N409);
   U1072 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_0_port, ZN => 
                           DATAPATH_I_N146);
   U1073 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_1_port, ZN => 
                           DATAPATH_I_N147);
   U1074 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_2_port, ZN => 
                           DATAPATH_I_N148);
   U1075 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_3_port, ZN => 
                           DATAPATH_I_N149);
   U1076 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_4_port, ZN => 
                           DATAPATH_I_N150);
   U1077 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_5_port, ZN => 
                           DATAPATH_I_N151);
   U1078 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_6_port, ZN => 
                           DATAPATH_I_N152);
   U1079 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_7_port, ZN => 
                           DATAPATH_I_N153);
   U1080 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_8_port, ZN => 
                           DATAPATH_I_N154);
   U1081 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_9_port, ZN => 
                           DATAPATH_I_N155);
   U1082 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_10_port, ZN => 
                           DATAPATH_I_N156);
   U1083 : AND2_X1 port map( A1 => RST, A2 => 
                           DATAPATH_I_ID_EX_RF_OUT2_NEXT_11_port, ZN => 
                           DATAPATH_I_N157);
   U1084 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_23_port,
                           ZN => DATAPATH_I_N266);
   U1085 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_13_port,
                           ZN => DATAPATH_I_N256);
   U1086 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_15_port,
                           ZN => DATAPATH_I_N258);
   U1087 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_20_port,
                           ZN => DATAPATH_I_N263);
   U1088 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_14_port,
                           ZN => DATAPATH_I_N257);
   U1089 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_22_port,
                           ZN => DATAPATH_I_N265);
   U1090 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_16_port,
                           ZN => DATAPATH_I_N259);
   U1091 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_17_port,
                           ZN => DATAPATH_I_N260);
   U1092 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_12_port,
                           ZN => DATAPATH_I_N255);
   U1093 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_21_port,
                           ZN => DATAPATH_I_N264);
   U1094 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_24_port,
                           ZN => DATAPATH_I_N267);
   U1095 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_25_port,
                           ZN => DATAPATH_I_N268);
   U1096 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_18_port,
                           ZN => DATAPATH_I_N261);
   U1097 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_19_port,
                           ZN => DATAPATH_I_N262);
   U1098 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_27_port,
                           ZN => DATAPATH_I_N270);
   U1099 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_28_port,
                           ZN => DATAPATH_I_N271);
   U1100 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_29_port,
                           ZN => DATAPATH_I_N272);
   U1101 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_30_port,
                           ZN => DATAPATH_I_N273);
   U1102 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_31_port,
                           ZN => DATAPATH_I_N274);
   U1103 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_11_port,
                           ZN => DATAPATH_I_N254);
   U1104 : AND2_X1 port map( A1 => RST, A2 => IR_30_port, ZN => DATAPATH_I_N64)
                           ;
   U1105 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_0_port, 
                           ZN => DATAPATH_I_N243);
   U1106 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_1_port, 
                           ZN => DATAPATH_I_N244);
   U1107 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_2_port, 
                           ZN => DATAPATH_I_N245);
   U1108 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_3_port, 
                           ZN => DATAPATH_I_N246);
   U1109 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_4_port, 
                           ZN => DATAPATH_I_N247);
   U1110 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_5_port, 
                           ZN => DATAPATH_I_N248);
   U1111 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_6_port, 
                           ZN => DATAPATH_I_N249);
   U1112 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_7_port, 
                           ZN => DATAPATH_I_N250);
   U1113 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_8_port, 
                           ZN => DATAPATH_I_N251);
   U1114 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_9_port, 
                           ZN => DATAPATH_I_N252);
   U1115 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_10_port,
                           ZN => DATAPATH_I_N253);
   U1116 : AND2_X1 port map( A1 => RST, A2 => DATAPATH_I_ID_EX_RF_OUT2_26_port,
                           ZN => DATAPATH_I_N269);
   U1117 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_19_port, A2 => n345, ZN 
                           => DATAPATH_I_ID_EX_RS2_NEXT_3_port);
   U1118 : AND2_X1 port map( A1 => DATAPATH_I_IF_ID_IR_24_port, A2 => n323, ZN 
                           => DATAPATH_I_ID_EX_RS1_NEXT_3_port);
   U1119 : INV_X1 port map( A => IR_26_port, ZN => n387);
   U1120 : NOR2_X1 port map( A1 => n317, A2 => n387, ZN => DATAPATH_I_N60);
   U1121 : INV_X1 port map( A => IR_5_port, ZN => n384);
   U1122 : OR4_X1 port map( A1 => IR_6_port, A2 => IR_9_port, A3 => IR_7_port, 
                           A4 => IR_8_port, ZN => n324);
   U1123 : NOR2_X1 port map( A1 => IR_10_port, A2 => n324, ZN => n325);
   U1124 : INV_X1 port map( A => IR_4_port, ZN => n327);
   U1125 : NAND2_X1 port map( A1 => n325, A2 => n327, ZN => n329);
   U1126 : NOR2_X1 port map( A1 => n384, A2 => n329, ZN => n332);
   U1127 : INV_X1 port map( A => n332, ZN => n328);
   U1128 : NOR2_X1 port map( A1 => IR_1_port, A2 => n328, ZN => n367);
   U1129 : INV_X1 port map( A => IR_1_port, ZN => n370);
   U1130 : INV_X1 port map( A => IR_2_port, ZN => n330);
   U1131 : NAND2_X1 port map( A1 => n325, A2 => IR_3_port, ZN => n326);
   U1132 : NOR2_X1 port map( A1 => n327, A2 => n326, ZN => n385);
   U1133 : NAND2_X1 port map( A1 => IR_5_port, A2 => n385, ZN => n375);
   U1134 : AOI221_X1 port map( B1 => IR_1_port, B2 => IR_2_port, C1 => n370, C2
                           => n330, A => n375, ZN => n383);
   U1135 : AOI21_X1 port map( B1 => IR_3_port, B2 => n367, A => n383, ZN => 
                           n405);
   U1136 : NOR2_X1 port map( A1 => IR_31_port, A2 => IR_30_port, ZN => n362);
   U1137 : INV_X1 port map( A => IR_29_port, ZN => n357);
   U1138 : NAND2_X1 port map( A1 => n362, A2 => n357, ZN => n408);
   U1139 : NOR4_X1 port map( A1 => IR_28_port, A2 => IR_27_port, A3 => 
                           IR_26_port, A4 => n408, ZN => n439);
   U1140 : INV_X1 port map( A => IR_3_port, ZN => n366);
   U1141 : NAND2_X1 port map( A1 => n330, A2 => IR_1_port, ZN => n376);
   U1142 : NOR2_X1 port map( A1 => n376, A2 => n328, ZN => n371);
   U1143 : OR4_X1 port map( A1 => IR_5_port, A2 => IR_3_port, A3 => n330, A4 =>
                           n329, ZN => n372);
   U1144 : NOR2_X1 port map( A1 => n370, A2 => n372, ZN => n380);
   U1145 : AOI21_X1 port map( B1 => n366, B2 => n371, A => n380, ZN => n331);
   U1146 : INV_X1 port map( A => n331, ZN => n404);
   U1147 : INV_X1 port map( A => n367, ZN => n418);
   U1148 : NOR2_X1 port map( A1 => IR_2_port, A2 => n418, ZN => n382);
   U1149 : INV_X1 port map( A => IR_0_port, ZN => n421);
   U1150 : OAI211_X1 port map( C1 => n404, C2 => n382, A => n366, B => n421, ZN
                           => n334);
   U1151 : NAND3_X1 port map( A1 => IR_3_port, A2 => n371, A3 => IR_0_port, ZN 
                           => n333);
   U1152 : NAND4_X1 port map( A1 => IR_2_port, A2 => n332, A3 => n366, A4 => 
                           n421, ZN => n369);
   U1153 : AND4_X1 port map( A1 => n439, A2 => n334, A3 => n333, A4 => n369, ZN
                           => n344);
   U1154 : NAND2_X1 port map( A1 => IR_29_port, A2 => n362, ZN => n406);
   U1155 : INV_X1 port map( A => n406, ZN => n430);
   U1156 : INV_X1 port map( A => DATAPATH_I_N62, ZN => n398);
   U1157 : NOR4_X1 port map( A1 => IR_27_port, A2 => n408, A3 => n387, A4 => 
                           n398, ZN => n342);
   U1158 : INV_X1 port map( A => IR_27_port, ZN => n356);
   U1159 : NAND2_X1 port map( A1 => IR_28_port, A2 => n356, ZN => n427);
   U1160 : NAND3_X1 port map( A1 => IR_29_port, A2 => IR_31_port, A3 => 
                           IR_30_port, ZN => n389);
   U1161 : NOR2_X1 port map( A1 => n427, A2 => n389, ZN => n336);
   U1162 : INV_X1 port map( A => IR_31_port, ZN => n358);
   U1163 : NAND3_X1 port map( A1 => IR_29_port, A2 => IR_30_port, A3 => n358, 
                           ZN => n400);
   U1164 : NAND2_X1 port map( A1 => IR_27_port, A2 => n407, ZN => n411);
   U1165 : NOR2_X1 port map( A1 => n400, A2 => n411, ZN => n359);
   U1166 : NAND2_X1 port map( A1 => n356, A2 => n387, ZN => n399);
   U1167 : INV_X1 port map( A => n439, ZN => n335);
   U1168 : OAI21_X1 port map( B1 => n399, B2 => n400, A => n335, ZN => n379);
   U1169 : AOI221_X1 port map( B1 => n336, B2 => IR_26_port, C1 => n359, C2 => 
                           n387, A => n379, ZN => n340);
   U1170 : INV_X1 port map( A => n411, ZN => n360);
   U1171 : NAND2_X1 port map( A1 => IR_26_port, A2 => n360, ZN => n390);
   U1172 : NOR3_X1 port map( A1 => IR_30_port, A2 => n358, A3 => n390, ZN => 
                           n417);
   U1173 : AOI21_X1 port map( B1 => n408, B2 => n389, A => n390, ZN => n338);
   U1174 : NAND3_X1 port map( A1 => IR_30_port, A2 => n357, A3 => n358, ZN => 
                           n412);
   U1175 : NOR3_X1 port map( A1 => n407, A2 => n356, A3 => n412, ZN => n402);
   U1176 : INV_X1 port map( A => n402, ZN => n337);
   U1177 : OAI22_X1 port map( A1 => IR_26_port, A2 => n337, B1 => n412, B2 => 
                           n390, ZN => n391);
   U1178 : AOI211_X1 port map( C1 => n417, C2 => n357, A => n338, B => n391, ZN
                           => n339);
   U1179 : AOI21_X1 port map( B1 => n340, B2 => n339, A => n317, ZN => n341);
   U1180 : AOI211_X1 port map( C1 => n430, C2 => DATAPATH_I_N60, A => n342, B 
                           => n341, ZN => n343);
   U1181 : AOI221_X1 port map( B1 => n405, B2 => n344, C1 => n421, C2 => n344, 
                           A => n343, ZN => CU_I_aluOpcode1_0_port);
   DATAPATH_I_MEM_WB_RF_WE <= '0';
   U1183 : NOR3_X1 port map( A1 => n347, A2 => n317, A3 => n345, ZN => n353);
   U1184 : NOR2_X1 port map( A1 => n317, A2 => n346, ZN => n352);
   U1185 : AOI22_X1 port map( A1 => DATAPATH_I_IF_ID_IR_16_port, A2 => n353, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_11_port, ZN => 
                           n348);
   U1186 : NAND3_X1 port map( A1 => RST, A2 => n347, A3 => 
                           DATAPATH_I_IF_ID_IR_26_port, ZN => n354);
   U1187 : NAND2_X1 port map( A1 => n348, A2 => n354, ZN => DATAPATH_I_N109);
   U1188 : AOI22_X1 port map( A1 => n353, A2 => DATAPATH_I_IF_ID_IR_17_port, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_12_port, ZN => 
                           n349);
   U1189 : NAND2_X1 port map( A1 => n349, A2 => n354, ZN => DATAPATH_I_N110);
   U1190 : AOI22_X1 port map( A1 => n353, A2 => DATAPATH_I_IF_ID_IR_18_port, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_13_port, ZN => 
                           n350);
   U1191 : NAND2_X1 port map( A1 => n350, A2 => n354, ZN => DATAPATH_I_N111);
   U1192 : AOI22_X1 port map( A1 => n353, A2 => DATAPATH_I_IF_ID_IR_19_port, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_14_port, ZN => 
                           n351);
   U1193 : NAND2_X1 port map( A1 => n351, A2 => n354, ZN => DATAPATH_I_N112);
   U1194 : AOI22_X1 port map( A1 => n353, A2 => DATAPATH_I_IF_ID_IR_20_port, B1
                           => n352, B2 => DATAPATH_I_IF_ID_IR_15_port, ZN => 
                           n355);
   U1195 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => DATAPATH_I_N113);
   U1196 : NOR2_X1 port map( A1 => n317, A2 => n356, ZN => DATAPATH_I_N61);
   U1197 : NOR2_X1 port map( A1 => n317, A2 => n357, ZN => DATAPATH_I_N63);
   U1198 : NOR2_X1 port map( A1 => n317, A2 => n358, ZN => DATAPATH_I_N65);
   U1199 : INV_X1 port map( A => n417, ZN => n365);
   U1200 : INV_X1 port map( A => n412, ZN => n388);
   U1201 : OAI221_X1 port map( B1 => IR_28_port, B2 => n388, C1 => n407, C2 => 
                           n430, A => IR_27_port, ZN => n424);
   U1202 : OAI21_X1 port map( B1 => n402, B2 => n359, A => IR_26_port, ZN => 
                           n364);
   U1203 : INV_X1 port map( A => n389, ZN => n361);
   U1204 : OAI21_X1 port map( B1 => n362, B2 => n361, A => n360, ZN => n363);
   U1205 : NAND4_X1 port map( A1 => n365, A2 => n424, A3 => n364, A4 => n363, 
                           ZN => n378);
   U1206 : NAND2_X1 port map( A1 => IR_0_port, A2 => n366, ZN => n381);
   U1207 : INV_X1 port map( A => n381, ZN => n373);
   U1208 : NAND3_X1 port map( A1 => IR_2_port, A2 => n373, A3 => n367, ZN => 
                           n368);
   U1209 : OAI21_X1 port map( B1 => n370, B2 => n369, A => n368, ZN => n397);
   U1210 : AOI21_X1 port map( B1 => n371, B2 => n381, A => n397, ZN => n419);
   U1211 : OAI21_X1 port map( B1 => IR_0_port, B2 => n372, A => n439, ZN => 
                           n403);
   U1212 : AOI21_X1 port map( B1 => n373, B2 => n382, A => n403, ZN => n374);
   U1213 : OAI211_X1 port map( C1 => n376, C2 => n375, A => n419, B => n374, ZN
                           => n377);
   U1214 : OAI211_X1 port map( C1 => n379, C2 => n378, A => RST, B => n377, ZN 
                           => CU_I_aluOpcode1_1_port);
   U1215 : AOI211_X1 port map( C1 => n382, C2 => n381, A => n380, B => n403, ZN
                           => n386);
   U1216 : INV_X1 port map( A => n383, ZN => n435);
   U1217 : NAND4_X1 port map( A1 => IR_1_port, A2 => IR_2_port, A3 => n385, A4 
                           => n384, ZN => n434);
   U1218 : NAND3_X1 port map( A1 => n386, A2 => n435, A3 => n434, ZN => n396);
   U1219 : OR2_X1 port map( A1 => n408, A2 => IR_27_port, ZN => n394);
   U1220 : NAND2_X1 port map( A1 => n427, A2 => n411, ZN => n429);
   U1221 : NAND2_X1 port map( A1 => n388, A2 => n387, ZN => n426);
   U1222 : NAND3_X1 port map( A1 => n406, A2 => n426, A3 => n389, ZN => n392);
   U1223 : AOI21_X1 port map( B1 => n427, B2 => n390, A => n400, ZN => n416);
   U1224 : AOI211_X1 port map( C1 => n429, C2 => n392, A => n416, B => n391, ZN
                           => n393);
   U1225 : OAI221_X1 port map( B1 => n394, B2 => IR_26_port, C1 => n394, C2 => 
                           n407, A => n393, ZN => n395);
   U1226 : OAI211_X1 port map( C1 => n397, C2 => n396, A => RST, B => n395, ZN 
                           => CU_I_aluOpcode1_2_port);
   U1227 : OR3_X1 port map( A1 => n399, A2 => n398, A3 => n412, ZN => n415);
   U1228 : AOI211_X1 port map( C1 => IR_27_port, C2 => IR_26_port, A => 
                           IR_28_port, B => n400, ZN => n401);
   U1229 : NOR2_X1 port map( A1 => n402, A2 => n401, ZN => n425);
   U1230 : NOR2_X1 port map( A1 => n404, A2 => n403, ZN => n420);
   U1231 : OAI211_X1 port map( C1 => IR_0_port, C2 => n434, A => n419, B => 
                           n405, ZN => n409);
   U1232 : AOI221_X1 port map( B1 => IR_28_port, B2 => n408, C1 => n407, C2 => 
                           n406, A => IR_27_port, ZN => n438);
   U1233 : AOI21_X1 port map( B1 => n420, B2 => n409, A => n438, ZN => n410);
   U1234 : OAI211_X1 port map( C1 => n412, C2 => n411, A => n425, B => n410, ZN
                           => n413);
   U1235 : AOI22_X1 port map( A1 => RST, A2 => n413, B1 => n417, B2 => 
                           DATAPATH_I_N63, ZN => n414);
   U1236 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => 
                           CU_I_aluOpcode1_3_port);
   U1237 : NOR2_X1 port map( A1 => n417, A2 => n416, ZN => n431);
   U1238 : AND3_X1 port map( A1 => n420, A2 => n419, A3 => n418, ZN => n436);
   U1239 : OAI21_X1 port map( B1 => n421, B2 => n434, A => n435, ZN => n422);
   U1240 : AOI21_X1 port map( B1 => n436, B2 => n422, A => n438, ZN => n423);
   U1241 : AOI21_X1 port map( B1 => n431, B2 => n423, A => n317, ZN => 
                           CU_I_aluOpcode1_4_port);
   U1242 : OAI211_X1 port map( C1 => n427, C2 => n426, A => n425, B => n424, ZN
                           => n428);
   U1243 : AOI211_X1 port map( C1 => n430, C2 => n429, A => n439, B => n428, ZN
                           => n432);
   U1244 : AOI22_X1 port map( A1 => n432, A2 => n431, B1 => n436, B2 => n435, 
                           ZN => n433);
   U1245 : NAND2_X1 port map( A1 => RST, A2 => n433, ZN => 
                           CU_I_aluOpcode1_5_port);
   U1246 : NAND3_X1 port map( A1 => n436, A2 => n435, A3 => n434, ZN => n437);
   U1247 : OAI211_X1 port map( C1 => n439, C2 => n438, A => RST, B => n437, ZN 
                           => CU_I_aluOpcode1_6_port);
   n285 <= '1';

end SYN_DLX_RTL;

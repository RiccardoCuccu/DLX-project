
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (OP_SLL, OP_SRL, OP_SRA, OP_ADD, OP_ADDU, OP_SUB, OP_SUBU, 
   OP_AND, OP_OR, OP_XOR, OP_SEQ, OP_SNE, OP_SLT, OP_SGT, OP_SLE, OP_SGE, 
   OP_MOVI2S, OP_MOVS2I, OP_MOVF, OP_MOVD, OP_MOVFP2I, OP_MOVI2FP, OP_MOVI2T, 
   OP_MOVT2I, OP_SLTU, OP_SGTU, OP_SLEU, OP_SGEU, OP_ADDF, OP_SUBF, OP_MULTF, 
   OP_DIVF, OP_ADDD, OP_SUBD, OP_MULTD, OP_DIVD, OP_CVTF2D, OP_CVTF2I, 
   OP_CVTD2F, OP_CVTD2I, OP_CVTI2F, OP_CVTI2D, OP_MULT, OP_DIV, OP_EQF, OP_NEF,
   OP_LTF, OP_GTF, OP_LEF, OP_GEF, OP_MULTU, OP_DIVU, OP_EQD, OP_NED, OP_LTD, 
   OP_GTD, OP_LED, OP_GED, OP_BEQZ, OP_BNEZ, OP_BFPT, OP_BFPF, OP_ADDI, 
   OP_ADDUI, OP_SUBI, OP_SUBUI, OP_ANDI, OP_ORI, OP_XORI, OP_LHI, OP_RFE, 
   OP_TRAP, OP_JR, OP_JALR, OP_SLLI, OP_SRLI, OP_SRAI, OP_SEQI, OP_SNEI, 
   OP_SLTI, OP_SGTI, OP_SLEI, OP_SGEI, OP_LB, OP_LH, OP_LW, OP_LBU, OP_LHU, 
   OP_LF, OP_LD, OP_SB, OP_SH, OP_SW, OP_SF, OP_SD, OP_ITLB, OP_SLTUI, 
   OP_SGTUI, OP_SLEUI, OP_SGEUI, OP_J, OP_JAL, OP_NOP);
attribute ENUM_ENCODING of aluOp : type is 
   "0000000 0000001 0000010 0000011 0000100 0000101 0000110 0000111 0001000 0001001 0001010 0001011 0001100 0001101 0001110 0001111 0010000 0010001 0010010 0010011 0010100 0010101 0010110 0010111 0011000 0011001 0011010 0011011 0011100 0011101 0011110 0011111 0100000 0100001 0100010 0100011 0100100 0100101 0100110 0100111 0101000 0101001 0101010 0101011 0101100 0101101 0101110 0101111 0110000 0110001 0110010 0110011 0110100 0110101 0110110 0110111 0111000 0111001 0111010 0111011 0111100 0111101 0111110 0111111 1000000 1000001 1000010 1000011 1000100 1000101 1000110 1000111 1001000 1001001 1001010 1001011 1001100 1001101 1001110 1001111 1010000 1010001 1010010 1010011 1010100 1010101 1010110 1010111 1011000 1011001 1011010 1011011 1011100 1011101 1011110 1011111 1100000 1100001 1100010 1100011 1100100 1100101 1100110";
   
   -- Declarations for conversion functions.
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when OP_SLL => return "0000000";
         when OP_SRL => return "0000001";
         when OP_SRA => return "0000010";
         when OP_ADD => return "0000011";
         when OP_ADDU => return "0000100";
         when OP_SUB => return "0000101";
         when OP_SUBU => return "0000110";
         when OP_AND => return "0000111";
         when OP_OR => return "0001000";
         when OP_XOR => return "0001001";
         when OP_SEQ => return "0001010";
         when OP_SNE => return "0001011";
         when OP_SLT => return "0001100";
         when OP_SGT => return "0001101";
         when OP_SLE => return "0001110";
         when OP_SGE => return "0001111";
         when OP_MOVI2S => return "0010000";
         when OP_MOVS2I => return "0010001";
         when OP_MOVF => return "0010010";
         when OP_MOVD => return "0010011";
         when OP_MOVFP2I => return "0010100";
         when OP_MOVI2FP => return "0010101";
         when OP_MOVI2T => return "0010110";
         when OP_MOVT2I => return "0010111";
         when OP_SLTU => return "0011000";
         when OP_SGTU => return "0011001";
         when OP_SLEU => return "0011010";
         when OP_SGEU => return "0011011";
         when OP_ADDF => return "0011100";
         when OP_SUBF => return "0011101";
         when OP_MULTF => return "0011110";
         when OP_DIVF => return "0011111";
         when OP_ADDD => return "0100000";
         when OP_SUBD => return "0100001";
         when OP_MULTD => return "0100010";
         when OP_DIVD => return "0100011";
         when OP_CVTF2D => return "0100100";
         when OP_CVTF2I => return "0100101";
         when OP_CVTD2F => return "0100110";
         when OP_CVTD2I => return "0100111";
         when OP_CVTI2F => return "0101000";
         when OP_CVTI2D => return "0101001";
         when OP_MULT => return "0101010";
         when OP_DIV => return "0101011";
         when OP_EQF => return "0101100";
         when OP_NEF => return "0101101";
         when OP_LTF => return "0101110";
         when OP_GTF => return "0101111";
         when OP_LEF => return "0110000";
         when OP_GEF => return "0110001";
         when OP_MULTU => return "0110010";
         when OP_DIVU => return "0110011";
         when OP_EQD => return "0110100";
         when OP_NED => return "0110101";
         when OP_LTD => return "0110110";
         when OP_GTD => return "0110111";
         when OP_LED => return "0111000";
         when OP_GED => return "0111001";
         when OP_BEQZ => return "0111010";
         when OP_BNEZ => return "0111011";
         when OP_BFPT => return "0111100";
         when OP_BFPF => return "0111101";
         when OP_ADDI => return "0111110";
         when OP_ADDUI => return "0111111";
         when OP_SUBI => return "1000000";
         when OP_SUBUI => return "1000001";
         when OP_ANDI => return "1000010";
         when OP_ORI => return "1000011";
         when OP_XORI => return "1000100";
         when OP_LHI => return "1000101";
         when OP_RFE => return "1000110";
         when OP_TRAP => return "1000111";
         when OP_JR => return "1001000";
         when OP_JALR => return "1001001";
         when OP_SLLI => return "1001010";
         when OP_SRLI => return "1001011";
         when OP_SRAI => return "1001100";
         when OP_SEQI => return "1001101";
         when OP_SNEI => return "1001110";
         when OP_SLTI => return "1001111";
         when OP_SGTI => return "1010000";
         when OP_SLEI => return "1010001";
         when OP_SGEI => return "1010010";
         when OP_LB => return "1010011";
         when OP_LH => return "1010100";
         when OP_LW => return "1010101";
         when OP_LBU => return "1010110";
         when OP_LHU => return "1010111";
         when OP_LF => return "1011000";
         when OP_LD => return "1011001";
         when OP_SB => return "1011010";
         when OP_SH => return "1011011";
         when OP_SW => return "1011100";
         when OP_SF => return "1011101";
         when OP_SD => return "1011110";
         when OP_ITLB => return "1011111";
         when OP_SLTUI => return "1100000";
         when OP_SGTUI => return "1100001";
         when OP_SLEUI => return "1100010";
         when OP_SGEUI => return "1100011";
         when OP_J => return "1100100";
         when OP_JAL => return "1100101";
         when OP_NOP => return "1100110";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

   port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  DOUT :
         out std_logic_vector (31 downto 0));

end DLX_IRAM_RAM_DEPTH256_I_SIZE32;

architecture SYN_BEHAVIORAL of DLX_IRAM_RAM_DEPTH256_I_SIZE32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_DRAM_N256_NW32 is

   port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector (31 
         downto 0);  DOUT : out std_logic_vector (31 downto 0));

end DLX_DRAM_N256_NW32;

architecture SYN_BEHAVIORAL of DLX_DRAM_N256_NW32 is

begin

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5;

architecture SYN_rpl of COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal GT_port, n203, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202 : std_logic;

begin
   GT <= GT_port;
   
   U1 : AND2_X1 port map( A1 => n2, A2 => n203, ZN => EQ);
   U2 : INV_X1 port map( A => n142, ZN => n51);
   U3 : INV_X1 port map( A => n130, ZN => n43);
   U4 : INV_X1 port map( A => n118, ZN => n35);
   U5 : INV_X1 port map( A => n106, ZN => n27);
   U6 : INV_X1 port map( A => n94, ZN => n19);
   U7 : INV_X1 port map( A => n82, ZN => n11);
   U8 : INV_X1 port map( A => n139, ZN => n49);
   U9 : INV_X1 port map( A => n127, ZN => n41);
   U10 : INV_X1 port map( A => n115, ZN => n33);
   U11 : INV_X1 port map( A => n103, ZN => n25);
   U12 : INV_X1 port map( A => n91, ZN => n17);
   U13 : INV_X1 port map( A => n79, ZN => n9);
   U14 : INV_X1 port map( A => n154, ZN => n59);
   U15 : INV_X1 port map( A => n144, ZN => n54);
   U16 : INV_X1 port map( A => n132, ZN => n46);
   U17 : INV_X1 port map( A => n120, ZN => n38);
   U18 : INV_X1 port map( A => n141, ZN => n52);
   U19 : INV_X1 port map( A => n129, ZN => n44);
   U20 : INV_X1 port map( A => n117, ZN => n36);
   U21 : INV_X1 port map( A => n108, ZN => n30);
   U22 : INV_X1 port map( A => n96, ZN => n22);
   U23 : INV_X1 port map( A => n84, ZN => n14);
   U24 : INV_X1 port map( A => n105, ZN => n28);
   U25 : INV_X1 port map( A => n93, ZN => n20);
   U26 : INV_X1 port map( A => n81, ZN => n12);
   U27 : INV_X1 port map( A => A(15), ZN => n34);
   U28 : INV_X1 port map( A => B(1), ZN => n65);
   U29 : INV_X1 port map( A => n68, ZN => n4);
   U30 : INV_X1 port map( A => A(30), ZN => n5);
   U31 : INV_X1 port map( A => n72, ZN => n6);
   U32 : INV_X1 port map( A => A(0), ZN => n62);
   U33 : INV_X1 port map( A => A(7), ZN => n50);
   U34 : INV_X1 port map( A => n151, ZN => n57);
   U35 : INV_X1 port map( A => A(3), ZN => n58);
   U36 : INV_X1 port map( A => A(11), ZN => n42);
   U37 : INV_X1 port map( A => A(14), ZN => n37);
   U38 : INV_X1 port map( A => A(6), ZN => n53);
   U39 : INV_X1 port map( A => A(10), ZN => n45);
   U40 : INV_X1 port map( A => A(2), ZN => n60);
   U41 : INV_X1 port map( A => A(8), ZN => n48);
   U42 : INV_X1 port map( A => A(4), ZN => n56);
   U43 : INV_X1 port map( A => A(12), ZN => n40);
   U44 : INV_X1 port map( A => A(13), ZN => n39);
   U45 : INV_X1 port map( A => A(5), ZN => n55);
   U46 : INV_X1 port map( A => A(9), ZN => n47);
   U47 : INV_X1 port map( A => GT_port, ZN => n2);
   U48 : INV_X1 port map( A => B(30), ZN => n64);
   U49 : INV_X1 port map( A => A(19), ZN => n26);
   U50 : INV_X1 port map( A => A(23), ZN => n18);
   U51 : INV_X1 port map( A => A(27), ZN => n10);
   U52 : INV_X1 port map( A => A(18), ZN => n29);
   U53 : INV_X1 port map( A => A(22), ZN => n21);
   U54 : INV_X1 port map( A => A(26), ZN => n13);
   U55 : INV_X1 port map( A => A(16), ZN => n32);
   U56 : INV_X1 port map( A => A(20), ZN => n24);
   U57 : INV_X1 port map( A => A(24), ZN => n16);
   U58 : INV_X1 port map( A => A(28), ZN => n8);
   U59 : INV_X1 port map( A => A(17), ZN => n31);
   U60 : INV_X1 port map( A => A(21), ZN => n23);
   U61 : INV_X1 port map( A => A(25), ZN => n15);
   U62 : INV_X1 port map( A => A(29), ZN => n7);
   U63 : INV_X1 port map( A => B(31), ZN => n63);
   U64 : INV_X1 port map( A => n203, ZN => LT);
   U65 : INV_X1 port map( A => n202, ZN => n61);
   U66 : AOI21_X1 port map( B1 => n66, B2 => n4, A => n67, ZN => n203);
   U67 : AOI22_X1 port map( A1 => B(30), A2 => n5, B1 => n69, B2 => n70, ZN => 
                           n68);
   U68 : AOI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n69);
   U69 : AOI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n71);
   U70 : AOI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n74);
   U71 : AOI21_X1 port map( B1 => n80, B2 => n11, A => n12, ZN => n77);
   U72 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n80);
   U73 : AOI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n83);
   U74 : AOI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n86);
   U75 : AOI21_X1 port map( B1 => n92, B2 => n19, A => n20, ZN => n89);
   U76 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n92);
   U77 : AOI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n95);
   U78 : AOI21_X1 port map( B1 => n101, B2 => n102, A => n103, ZN => n98);
   U79 : AOI21_X1 port map( B1 => n104, B2 => n27, A => n28, ZN => n101);
   U80 : AOI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n104);
   U81 : AOI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n107);
   U82 : AOI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n110);
   U83 : AOI21_X1 port map( B1 => n116, B2 => n35, A => n36, ZN => n113);
   U84 : AOI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n116);
   U85 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n119);
   U86 : AOI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n122);
   U87 : AOI21_X1 port map( B1 => n128, B2 => n43, A => n44, ZN => n125);
   U88 : AOI21_X1 port map( B1 => n131, B2 => n132, A => n133, ZN => n128);
   U89 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n131);
   U90 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n134);
   U91 : AOI21_X1 port map( B1 => n140, B2 => n51, A => n52, ZN => n137);
   U92 : AOI21_X1 port map( B1 => n143, B2 => n144, A => n145, ZN => n140);
   U93 : AOI21_X1 port map( B1 => n146, B2 => n147, A => n148, ZN => n143);
   U94 : AOI21_X1 port map( B1 => n149, B2 => n150, A => n151, ZN => n146);
   U95 : AOI21_X1 port map( B1 => n152, B2 => n153, A => n59, ZN => n149);
   U96 : AOI22_X1 port map( A1 => n155, A2 => n65, B1 => A(1), B2 => n156, ZN 
                           => n152);
   U97 : OR2_X1 port map( A1 => n156, A2 => A(1), ZN => n155);
   U98 : NAND2_X1 port map( A1 => B(0), A2 => n62, ZN => n156);
   U99 : OAI21_X1 port map( B1 => n67, B2 => n157, A => n66, ZN => GT_port);
   U100 : NAND2_X1 port map( A1 => A(31), A2 => n63, ZN => n66);
   U101 : AOI22_X1 port map( A1 => A(30), A2 => n64, B1 => n158, B2 => n70, ZN 
                           => n157);
   U102 : XOR2_X1 port map( A => A(30), B => n64, Z => n70);
   U103 : AOI21_X1 port map( B1 => n159, B2 => n160, A => n6, ZN => n158);
   U104 : NAND2_X1 port map( A1 => B(29), A2 => n7, ZN => n72);
   U105 : OAI211_X1 port map( C1 => n161, C2 => n162, A => n78, B => n75, ZN =>
                           n160);
   U106 : NOR2_X1 port map( A1 => n163, A2 => n76, ZN => n75);
   U107 : AND2_X1 port map( A1 => B(28), A2 => n8, ZN => n76);
   U108 : NAND2_X1 port map( A1 => B(27), A2 => n10, ZN => n78);
   U109 : NAND2_X1 port map( A1 => n9, A2 => n164, ZN => n162);
   U110 : NOR2_X1 port map( A1 => n10, A2 => B(27), ZN => n79);
   U111 : AOI211_X1 port map( C1 => n165, C2 => n166, A => n82, B => n14, ZN =>
                           n161);
   U112 : NAND2_X1 port map( A1 => B(25), A2 => n15, ZN => n84);
   U113 : NAND2_X1 port map( A1 => n164, A2 => n81, ZN => n82);
   U114 : NAND2_X1 port map( A1 => B(26), A2 => n13, ZN => n81);
   U115 : OR2_X1 port map( A1 => n13, A2 => B(26), ZN => n164);
   U116 : OAI211_X1 port map( C1 => n167, C2 => n168, A => n90, B => n87, ZN =>
                           n166);
   U117 : NOR2_X1 port map( A1 => n169, A2 => n88, ZN => n87);
   U118 : AND2_X1 port map( A1 => B(24), A2 => n16, ZN => n88);
   U119 : NAND2_X1 port map( A1 => B(23), A2 => n18, ZN => n90);
   U120 : NAND2_X1 port map( A1 => n17, A2 => n170, ZN => n168);
   U121 : NOR2_X1 port map( A1 => n18, A2 => B(23), ZN => n91);
   U122 : AOI211_X1 port map( C1 => n171, C2 => n172, A => n94, B => n22, ZN =>
                           n167);
   U123 : NAND2_X1 port map( A1 => B(21), A2 => n23, ZN => n96);
   U124 : NAND2_X1 port map( A1 => n170, A2 => n93, ZN => n94);
   U125 : NAND2_X1 port map( A1 => B(22), A2 => n21, ZN => n93);
   U126 : OR2_X1 port map( A1 => n21, A2 => B(22), ZN => n170);
   U127 : OAI211_X1 port map( C1 => n173, C2 => n174, A => n102, B => n99, ZN 
                           => n172);
   U128 : NOR2_X1 port map( A1 => n175, A2 => n100, ZN => n99);
   U129 : AND2_X1 port map( A1 => B(20), A2 => n24, ZN => n100);
   U130 : NAND2_X1 port map( A1 => B(19), A2 => n26, ZN => n102);
   U131 : NAND2_X1 port map( A1 => n25, A2 => n176, ZN => n174);
   U132 : NOR2_X1 port map( A1 => n26, A2 => B(19), ZN => n103);
   U133 : AOI211_X1 port map( C1 => n177, C2 => n178, A => n106, B => n30, ZN 
                           => n173);
   U134 : NAND2_X1 port map( A1 => B(17), A2 => n31, ZN => n108);
   U135 : NAND2_X1 port map( A1 => n176, A2 => n105, ZN => n106);
   U136 : NAND2_X1 port map( A1 => B(18), A2 => n29, ZN => n105);
   U137 : OR2_X1 port map( A1 => n29, A2 => B(18), ZN => n176);
   U138 : OAI211_X1 port map( C1 => n179, C2 => n180, A => n114, B => n111, ZN 
                           => n178);
   U139 : NOR2_X1 port map( A1 => n181, A2 => n112, ZN => n111);
   U140 : AND2_X1 port map( A1 => B(16), A2 => n32, ZN => n112);
   U141 : NAND2_X1 port map( A1 => B(15), A2 => n34, ZN => n114);
   U142 : NAND2_X1 port map( A1 => n33, A2 => n182, ZN => n180);
   U143 : NOR2_X1 port map( A1 => n34, A2 => B(15), ZN => n115);
   U144 : AOI211_X1 port map( C1 => n183, C2 => n184, A => n118, B => n38, ZN 
                           => n179);
   U145 : NAND2_X1 port map( A1 => B(13), A2 => n39, ZN => n120);
   U146 : NAND2_X1 port map( A1 => n182, A2 => n117, ZN => n118);
   U147 : NAND2_X1 port map( A1 => B(14), A2 => n37, ZN => n117);
   U148 : OR2_X1 port map( A1 => n37, A2 => B(14), ZN => n182);
   U149 : OAI211_X1 port map( C1 => n185, C2 => n186, A => n126, B => n123, ZN 
                           => n184);
   U150 : NOR2_X1 port map( A1 => n187, A2 => n124, ZN => n123);
   U151 : AND2_X1 port map( A1 => B(12), A2 => n40, ZN => n124);
   U152 : NAND2_X1 port map( A1 => B(11), A2 => n42, ZN => n126);
   U153 : NAND2_X1 port map( A1 => n41, A2 => n188, ZN => n186);
   U154 : NOR2_X1 port map( A1 => n42, A2 => B(11), ZN => n127);
   U155 : AOI211_X1 port map( C1 => n189, C2 => n190, A => n130, B => n46, ZN 
                           => n185);
   U156 : NAND2_X1 port map( A1 => B(9), A2 => n47, ZN => n132);
   U157 : NAND2_X1 port map( A1 => n188, A2 => n129, ZN => n130);
   U158 : NAND2_X1 port map( A1 => B(10), A2 => n45, ZN => n129);
   U159 : OR2_X1 port map( A1 => n45, A2 => B(10), ZN => n188);
   U160 : OAI211_X1 port map( C1 => n191, C2 => n192, A => n138, B => n135, ZN 
                           => n190);
   U161 : NOR2_X1 port map( A1 => n193, A2 => n136, ZN => n135);
   U162 : AND2_X1 port map( A1 => B(8), A2 => n48, ZN => n136);
   U163 : NAND2_X1 port map( A1 => B(7), A2 => n50, ZN => n138);
   U164 : NAND2_X1 port map( A1 => n49, A2 => n194, ZN => n192);
   U165 : NOR2_X1 port map( A1 => n50, A2 => B(7), ZN => n139);
   U166 : AOI211_X1 port map( C1 => n195, C2 => n196, A => n142, B => n54, ZN 
                           => n191);
   U167 : NAND2_X1 port map( A1 => B(5), A2 => n55, ZN => n144);
   U168 : NAND2_X1 port map( A1 => n194, A2 => n141, ZN => n142);
   U169 : NAND2_X1 port map( A1 => B(6), A2 => n53, ZN => n141);
   U170 : OR2_X1 port map( A1 => n53, A2 => B(6), ZN => n194);
   U171 : NAND3_X1 port map( A1 => n197, A2 => n150, A3 => n147, ZN => n196);
   U172 : NOR2_X1 port map( A1 => n198, A2 => n148, ZN => n147);
   U173 : AND2_X1 port map( A1 => B(4), A2 => n56, ZN => n148);
   U174 : NAND2_X1 port map( A1 => B(3), A2 => n58, ZN => n150);
   U175 : NAND3_X1 port map( A1 => n57, A2 => n199, A3 => n200, ZN => n197);
   U176 : OAI211_X1 port map( C1 => A(1), C2 => n201, A => n61, B => n153, ZN 
                           => n200);
   U177 : AND2_X1 port map( A1 => n199, A2 => n154, ZN => n153);
   U178 : NAND2_X1 port map( A1 => B(2), A2 => n60, ZN => n154);
   U179 : AOI21_X1 port map( B1 => A(1), B2 => n201, A => n65, ZN => n202);
   U180 : NOR2_X1 port map( A1 => n62, A2 => B(0), ZN => n201);
   U181 : OR2_X1 port map( A1 => n60, A2 => B(2), ZN => n199);
   U182 : NOR2_X1 port map( A1 => n58, A2 => B(3), ZN => n151);
   U183 : NOR2_X1 port map( A1 => n198, A2 => n145, ZN => n195);
   U184 : NOR2_X1 port map( A1 => n55, A2 => B(5), ZN => n145);
   U185 : NOR2_X1 port map( A1 => n56, A2 => B(4), ZN => n198);
   U186 : NOR2_X1 port map( A1 => n193, A2 => n133, ZN => n189);
   U187 : NOR2_X1 port map( A1 => n47, A2 => B(9), ZN => n133);
   U188 : NOR2_X1 port map( A1 => n48, A2 => B(8), ZN => n193);
   U189 : NOR2_X1 port map( A1 => n187, A2 => n121, ZN => n183);
   U190 : NOR2_X1 port map( A1 => n39, A2 => B(13), ZN => n121);
   U191 : NOR2_X1 port map( A1 => n40, A2 => B(12), ZN => n187);
   U192 : NOR2_X1 port map( A1 => n181, A2 => n109, ZN => n177);
   U193 : NOR2_X1 port map( A1 => n31, A2 => B(17), ZN => n109);
   U194 : NOR2_X1 port map( A1 => n32, A2 => B(16), ZN => n181);
   U195 : NOR2_X1 port map( A1 => n175, A2 => n97, ZN => n171);
   U196 : NOR2_X1 port map( A1 => n23, A2 => B(21), ZN => n97);
   U197 : NOR2_X1 port map( A1 => n24, A2 => B(20), ZN => n175);
   U198 : NOR2_X1 port map( A1 => n169, A2 => n85, ZN => n165);
   U199 : NOR2_X1 port map( A1 => n15, A2 => B(25), ZN => n85);
   U200 : NOR2_X1 port map( A1 => n16, A2 => B(24), ZN => n169);
   U201 : NOR2_X1 port map( A1 => n163, A2 => n73, ZN => n159);
   U202 : NOR2_X1 port map( A1 => n7, A2 => B(29), ZN => n73);
   U203 : NOR2_X1 port map( A1 => n8, A2 => B(28), ZN => n163);
   U204 : NOR2_X1 port map( A1 => n63, A2 => A(31), ZN => n67);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4;

architecture SYN_rpl of COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n202, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30
      , n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88
      , n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102
      , n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n131, ZN => n26);
   U2 : INV_X1 port map( A => n111, ZN => n18);
   U3 : INV_X1 port map( A => n91, ZN => n10);
   U4 : INV_X1 port map( A => n137, ZN => n30);
   U5 : INV_X1 port map( A => n121, ZN => n22);
   U6 : INV_X1 port map( A => n122, ZN => n24);
   U7 : INV_X1 port map( A => n127, ZN => n25);
   U8 : INV_X1 port map( A => n101, ZN => n14);
   U9 : INV_X1 port map( A => n102, ZN => n16);
   U10 : INV_X1 port map( A => n81, ZN => n6);
   U11 : INV_X1 port map( A => n82, ZN => n8);
   U12 : INV_X1 port map( A => n107, ZN => n17);
   U13 : INV_X1 port map( A => n87, ZN => n9);
   U14 : INV_X1 port map( A => n132, ZN => n28);
   U15 : INV_X1 port map( A => n112, ZN => n20);
   U16 : INV_X1 port map( A => n92, ZN => n12);
   U17 : INV_X1 port map( A => n72, ZN => n4);
   U18 : INV_X1 port map( A => n181, ZN => n19);
   U19 : INV_X1 port map( A => n193, ZN => n27);
   U20 : INV_X1 port map( A => n187, ZN => n23);
   U21 : INV_X1 port map( A => n175, ZN => n15);
   U22 : INV_X1 port map( A => n169, ZN => n11);
   U23 : INV_X1 port map( A => n163, ZN => n7);
   U24 : INV_X1 port map( A => n136, ZN => n29);
   U25 : INV_X1 port map( A => n117, ZN => n21);
   U26 : INV_X1 port map( A => n97, ZN => n13);
   U27 : INV_X1 port map( A => n77, ZN => n5);
   U28 : INV_X1 port map( A => B(0), ZN => n64);
   U29 : INV_X1 port map( A => B(3), ZN => n62);
   U30 : INV_X1 port map( A => B(4), ZN => n61);
   U31 : INV_X1 port map( A => B(2), ZN => n63);
   U32 : INV_X1 port map( A => A(1), ZN => n32);
   U33 : INV_X1 port map( A => n199, ZN => n31);
   U34 : INV_X1 port map( A => A(30), ZN => n3);
   U35 : INV_X1 port map( A => n202, ZN => GT);
   U36 : INV_X1 port map( A => B(7), ZN => n58);
   U37 : INV_X1 port map( A => B(11), ZN => n54);
   U38 : INV_X1 port map( A => B(5), ZN => n60);
   U39 : INV_X1 port map( A => B(9), ZN => n56);
   U40 : INV_X1 port map( A => B(13), ZN => n52);
   U41 : INV_X1 port map( A => B(8), ZN => n57);
   U42 : INV_X1 port map( A => B(12), ZN => n53);
   U43 : INV_X1 port map( A => n141, ZN => n33);
   U44 : INV_X1 port map( A => B(15), ZN => n50);
   U45 : INV_X1 port map( A => B(6), ZN => n59);
   U46 : INV_X1 port map( A => B(10), ZN => n55);
   U47 : INV_X1 port map( A => B(14), ZN => n51);
   U48 : INV_X1 port map( A => B(16), ZN => n49);
   U49 : INV_X1 port map( A => B(20), ZN => n45);
   U50 : INV_X1 port map( A => B(24), ZN => n41);
   U51 : INV_X1 port map( A => B(28), ZN => n37);
   U52 : INV_X1 port map( A => B(31), ZN => n34);
   U53 : INV_X1 port map( A => B(18), ZN => n47);
   U54 : INV_X1 port map( A => B(22), ZN => n43);
   U55 : INV_X1 port map( A => B(26), ZN => n39);
   U56 : INV_X1 port map( A => B(19), ZN => n46);
   U57 : INV_X1 port map( A => B(23), ZN => n42);
   U58 : INV_X1 port map( A => B(27), ZN => n38);
   U59 : INV_X1 port map( A => B(17), ZN => n48);
   U60 : INV_X1 port map( A => B(21), ZN => n44);
   U61 : INV_X1 port map( A => B(25), ZN => n40);
   U62 : INV_X1 port map( A => B(29), ZN => n36);
   U63 : INV_X1 port map( A => n67, ZN => n2);
   U64 : INV_X1 port map( A => B(30), ZN => n35);
   U65 : AOI21_X1 port map( B1 => n65, B2 => n2, A => n66, ZN => n202);
   U66 : AOI22_X1 port map( A1 => A(30), A2 => n35, B1 => n68, B2 => n69, ZN =>
                           n67);
   U67 : AOI21_X1 port map( B1 => n70, B2 => n71, A => n72, ZN => n68);
   U68 : OAI211_X1 port map( C1 => n73, C2 => n74, A => n75, B => n76, ZN => 
                           n71);
   U69 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => n74);
   U70 : AOI211_X1 port map( C1 => n79, C2 => n80, A => n81, B => n82, ZN => 
                           n73);
   U71 : OAI211_X1 port map( C1 => n83, C2 => n84, A => n85, B => n86, ZN => 
                           n80);
   U72 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => n84);
   U73 : AOI211_X1 port map( C1 => n89, C2 => n90, A => n91, B => n92, ZN => 
                           n83);
   U74 : OAI211_X1 port map( C1 => n93, C2 => n94, A => n95, B => n96, ZN => 
                           n90);
   U75 : NAND2_X1 port map( A1 => n97, A2 => n98, ZN => n94);
   U76 : AOI211_X1 port map( C1 => n99, C2 => n100, A => n101, B => n102, ZN =>
                           n93);
   U77 : OAI211_X1 port map( C1 => n103, C2 => n104, A => n105, B => n106, ZN 
                           => n100);
   U78 : NAND2_X1 port map( A1 => n107, A2 => n108, ZN => n104);
   U79 : AOI211_X1 port map( C1 => n109, C2 => n110, A => n111, B => n112, ZN 
                           => n103);
   U80 : OAI211_X1 port map( C1 => n113, C2 => n114, A => n115, B => n116, ZN 
                           => n110);
   U81 : NAND2_X1 port map( A1 => n117, A2 => n118, ZN => n114);
   U82 : AOI211_X1 port map( C1 => n119, C2 => n120, A => n121, B => n122, ZN 
                           => n113);
   U83 : OAI211_X1 port map( C1 => n123, C2 => n124, A => n125, B => n126, ZN 
                           => n120);
   U84 : NAND2_X1 port map( A1 => n127, A2 => n128, ZN => n124);
   U85 : AOI211_X1 port map( C1 => n129, C2 => n130, A => n131, B => n132, ZN 
                           => n123);
   U86 : NAND3_X1 port map( A1 => n133, A2 => n134, A3 => n135, ZN => n130);
   U87 : NAND3_X1 port map( A1 => n136, A2 => n137, A3 => n138, ZN => n133);
   U88 : OAI211_X1 port map( C1 => A(1), C2 => n33, A => n139, B => n140, ZN =>
                           n138);
   U89 : OAI21_X1 port map( B1 => n32, B2 => n141, A => B(1), ZN => n139);
   U90 : NAND2_X1 port map( A1 => A(0), A2 => n64, ZN => n141);
   U91 : NOR2_X1 port map( A1 => n142, A2 => n143, ZN => n129);
   U92 : NOR2_X1 port map( A1 => n144, A2 => n145, ZN => n119);
   U93 : NOR2_X1 port map( A1 => n146, A2 => n147, ZN => n109);
   U94 : NOR2_X1 port map( A1 => n148, A2 => n149, ZN => n99);
   U95 : NOR2_X1 port map( A1 => n150, A2 => n151, ZN => n89);
   U96 : NOR2_X1 port map( A1 => n152, A2 => n153, ZN => n79);
   U97 : NOR2_X1 port map( A1 => n154, A2 => n155, ZN => n70);
   U98 : OAI21_X1 port map( B1 => n66, B2 => n156, A => n65, ZN => LT);
   U99 : NAND2_X1 port map( A1 => A(31), A2 => n34, ZN => n65);
   U100 : AOI22_X1 port map( A1 => B(30), A2 => n3, B1 => n157, B2 => n69, ZN 
                           => n156);
   U101 : XOR2_X1 port map( A => n3, B => B(30), Z => n69);
   U102 : AOI21_X1 port map( B1 => n158, B2 => n4, A => n155, ZN => n157);
   U103 : AND2_X1 port map( A1 => A(29), A2 => n36, ZN => n155);
   U104 : NOR2_X1 port map( A1 => n36, A2 => A(29), ZN => n72);
   U105 : AOI21_X1 port map( B1 => n159, B2 => n76, A => n160, ZN => n158);
   U106 : NOR2_X1 port map( A1 => n160, A2 => n154, ZN => n76);
   U107 : AND2_X1 port map( A1 => A(28), A2 => n37, ZN => n154);
   U108 : NOR2_X1 port map( A1 => n37, A2 => A(28), ZN => n160);
   U109 : AOI21_X1 port map( B1 => n161, B2 => n75, A => n5, ZN => n159);
   U110 : NAND2_X1 port map( A1 => A(27), A2 => n38, ZN => n77);
   U111 : OR2_X1 port map( A1 => n38, A2 => A(27), ZN => n75);
   U112 : AOI21_X1 port map( B1 => n162, B2 => n6, A => n163, ZN => n161);
   U113 : NAND2_X1 port map( A1 => n7, A2 => n78, ZN => n81);
   U114 : NAND2_X1 port map( A1 => A(26), A2 => n39, ZN => n78);
   U115 : NOR2_X1 port map( A1 => n39, A2 => A(26), ZN => n163);
   U116 : AOI21_X1 port map( B1 => n164, B2 => n8, A => n153, ZN => n162);
   U117 : AND2_X1 port map( A1 => A(25), A2 => n40, ZN => n153);
   U118 : NOR2_X1 port map( A1 => n40, A2 => A(25), ZN => n82);
   U119 : AOI21_X1 port map( B1 => n165, B2 => n86, A => n166, ZN => n164);
   U120 : NOR2_X1 port map( A1 => n166, A2 => n152, ZN => n86);
   U121 : AND2_X1 port map( A1 => A(24), A2 => n41, ZN => n152);
   U122 : NOR2_X1 port map( A1 => n41, A2 => A(24), ZN => n166);
   U123 : AOI21_X1 port map( B1 => n167, B2 => n85, A => n9, ZN => n165);
   U124 : NAND2_X1 port map( A1 => A(23), A2 => n42, ZN => n87);
   U125 : OR2_X1 port map( A1 => n42, A2 => A(23), ZN => n85);
   U126 : AOI21_X1 port map( B1 => n168, B2 => n10, A => n169, ZN => n167);
   U127 : NAND2_X1 port map( A1 => n11, A2 => n88, ZN => n91);
   U128 : NAND2_X1 port map( A1 => A(22), A2 => n43, ZN => n88);
   U129 : NOR2_X1 port map( A1 => n43, A2 => A(22), ZN => n169);
   U130 : AOI21_X1 port map( B1 => n170, B2 => n12, A => n151, ZN => n168);
   U131 : AND2_X1 port map( A1 => A(21), A2 => n44, ZN => n151);
   U132 : NOR2_X1 port map( A1 => n44, A2 => A(21), ZN => n92);
   U133 : AOI21_X1 port map( B1 => n171, B2 => n96, A => n172, ZN => n170);
   U134 : NOR2_X1 port map( A1 => n172, A2 => n150, ZN => n96);
   U135 : AND2_X1 port map( A1 => A(20), A2 => n45, ZN => n150);
   U136 : NOR2_X1 port map( A1 => n45, A2 => A(20), ZN => n172);
   U137 : AOI21_X1 port map( B1 => n173, B2 => n95, A => n13, ZN => n171);
   U138 : NAND2_X1 port map( A1 => A(19), A2 => n46, ZN => n97);
   U139 : OR2_X1 port map( A1 => n46, A2 => A(19), ZN => n95);
   U140 : AOI21_X1 port map( B1 => n174, B2 => n14, A => n175, ZN => n173);
   U141 : NAND2_X1 port map( A1 => n15, A2 => n98, ZN => n101);
   U142 : NAND2_X1 port map( A1 => A(18), A2 => n47, ZN => n98);
   U143 : NOR2_X1 port map( A1 => n47, A2 => A(18), ZN => n175);
   U144 : AOI21_X1 port map( B1 => n176, B2 => n16, A => n149, ZN => n174);
   U145 : AND2_X1 port map( A1 => A(17), A2 => n48, ZN => n149);
   U146 : NOR2_X1 port map( A1 => n48, A2 => A(17), ZN => n102);
   U147 : AOI21_X1 port map( B1 => n177, B2 => n106, A => n178, ZN => n176);
   U148 : NOR2_X1 port map( A1 => n178, A2 => n148, ZN => n106);
   U149 : AND2_X1 port map( A1 => A(16), A2 => n49, ZN => n148);
   U150 : NOR2_X1 port map( A1 => n49, A2 => A(16), ZN => n178);
   U151 : AOI21_X1 port map( B1 => n179, B2 => n105, A => n17, ZN => n177);
   U152 : NAND2_X1 port map( A1 => A(15), A2 => n50, ZN => n107);
   U153 : OR2_X1 port map( A1 => n50, A2 => A(15), ZN => n105);
   U154 : AOI21_X1 port map( B1 => n180, B2 => n18, A => n181, ZN => n179);
   U155 : NAND2_X1 port map( A1 => n19, A2 => n108, ZN => n111);
   U156 : NAND2_X1 port map( A1 => A(14), A2 => n51, ZN => n108);
   U157 : NOR2_X1 port map( A1 => n51, A2 => A(14), ZN => n181);
   U158 : AOI21_X1 port map( B1 => n182, B2 => n20, A => n147, ZN => n180);
   U159 : AND2_X1 port map( A1 => A(13), A2 => n52, ZN => n147);
   U160 : NOR2_X1 port map( A1 => n52, A2 => A(13), ZN => n112);
   U161 : AOI21_X1 port map( B1 => n183, B2 => n116, A => n184, ZN => n182);
   U162 : NOR2_X1 port map( A1 => n184, A2 => n146, ZN => n116);
   U163 : AND2_X1 port map( A1 => A(12), A2 => n53, ZN => n146);
   U164 : NOR2_X1 port map( A1 => n53, A2 => A(12), ZN => n184);
   U165 : AOI21_X1 port map( B1 => n185, B2 => n115, A => n21, ZN => n183);
   U166 : NAND2_X1 port map( A1 => A(11), A2 => n54, ZN => n117);
   U167 : OR2_X1 port map( A1 => n54, A2 => A(11), ZN => n115);
   U168 : AOI21_X1 port map( B1 => n186, B2 => n22, A => n187, ZN => n185);
   U169 : NAND2_X1 port map( A1 => n23, A2 => n118, ZN => n121);
   U170 : NAND2_X1 port map( A1 => A(10), A2 => n55, ZN => n118);
   U171 : NOR2_X1 port map( A1 => n55, A2 => A(10), ZN => n187);
   U172 : AOI21_X1 port map( B1 => n188, B2 => n24, A => n145, ZN => n186);
   U173 : AND2_X1 port map( A1 => A(9), A2 => n56, ZN => n145);
   U174 : NOR2_X1 port map( A1 => n56, A2 => A(9), ZN => n122);
   U175 : AOI21_X1 port map( B1 => n189, B2 => n126, A => n190, ZN => n188);
   U176 : NOR2_X1 port map( A1 => n190, A2 => n144, ZN => n126);
   U177 : AND2_X1 port map( A1 => A(8), A2 => n57, ZN => n144);
   U178 : NOR2_X1 port map( A1 => n57, A2 => A(8), ZN => n190);
   U179 : AOI21_X1 port map( B1 => n191, B2 => n125, A => n25, ZN => n189);
   U180 : NAND2_X1 port map( A1 => A(7), A2 => n58, ZN => n127);
   U181 : OR2_X1 port map( A1 => n58, A2 => A(7), ZN => n125);
   U182 : AOI21_X1 port map( B1 => n192, B2 => n26, A => n193, ZN => n191);
   U183 : NAND2_X1 port map( A1 => n27, A2 => n128, ZN => n131);
   U184 : NAND2_X1 port map( A1 => A(6), A2 => n59, ZN => n128);
   U185 : NOR2_X1 port map( A1 => n59, A2 => A(6), ZN => n193);
   U186 : AOI21_X1 port map( B1 => n194, B2 => n28, A => n143, ZN => n192);
   U187 : AND2_X1 port map( A1 => A(5), A2 => n60, ZN => n143);
   U188 : NOR2_X1 port map( A1 => n60, A2 => A(5), ZN => n132);
   U189 : AOI21_X1 port map( B1 => n195, B2 => n135, A => n196, ZN => n194);
   U190 : NOR2_X1 port map( A1 => n196, A2 => n142, ZN => n135);
   U191 : AND2_X1 port map( A1 => A(4), A2 => n61, ZN => n142);
   U192 : NOR2_X1 port map( A1 => n61, A2 => A(4), ZN => n196);
   U193 : AOI21_X1 port map( B1 => n197, B2 => n134, A => n29, ZN => n195);
   U194 : NAND2_X1 port map( A1 => A(3), A2 => n62, ZN => n136);
   U195 : OR2_X1 port map( A1 => n62, A2 => A(3), ZN => n134);
   U196 : AOI21_X1 port map( B1 => n31, B2 => n140, A => n198, ZN => n197);
   U197 : NOR2_X1 port map( A1 => n198, A2 => n30, ZN => n140);
   U198 : NAND2_X1 port map( A1 => A(2), A2 => n63, ZN => n137);
   U199 : NOR2_X1 port map( A1 => n63, A2 => A(2), ZN => n198);
   U200 : OAI22_X1 port map( A1 => n200, A2 => B(1), B1 => n32, B2 => n201, ZN 
                           => n199);
   U201 : AND2_X1 port map( A1 => n201, A2 => n32, ZN => n200);
   U202 : NOR2_X1 port map( A1 => n64, A2 => A(0), ZN => n201);
   U203 : NOR2_X1 port map( A1 => n34, A2 => A(31), ZN => n66);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity 
   DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0 
   is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0
   ;

architecture SYN_rpl of 
   DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0 
   is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, SUM_30_port, 
      SUM_29_port, SUM_28_port, SUM_27_port, SUM_26_port, SUM_25_port, 
      SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, 
      SUM_19_port, SUM_18_port, SUM_17_port, SUM_16_port, SUM_15_port, 
      SUM_14_port, SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, 
      SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port, SUM_5_port, SUM_4_port, 
      SUM_3_port, SUM_31_port, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n1);
   U2 : AND2_X1 port map( A1 => A(4), A2 => n1, ZN => n2);
   U3 : AND2_X1 port map( A1 => A(5), A2 => n2, ZN => n3);
   U4 : AND2_X1 port map( A1 => A(6), A2 => n3, ZN => n4);
   U5 : AND2_X1 port map( A1 => A(7), A2 => n4, ZN => n5);
   U6 : AND2_X1 port map( A1 => A(8), A2 => n5, ZN => n6);
   U7 : AND2_X1 port map( A1 => A(9), A2 => n6, ZN => n7);
   U8 : AND2_X1 port map( A1 => A(10), A2 => n7, ZN => n8);
   U9 : AND2_X1 port map( A1 => A(11), A2 => n8, ZN => n9);
   U10 : AND2_X1 port map( A1 => A(12), A2 => n9, ZN => n10);
   U11 : AND2_X1 port map( A1 => A(13), A2 => n10, ZN => n11);
   U12 : AND2_X1 port map( A1 => A(14), A2 => n11, ZN => n12);
   U13 : AND2_X1 port map( A1 => A(15), A2 => n12, ZN => n13);
   U14 : AND2_X1 port map( A1 => A(16), A2 => n13, ZN => n14);
   U15 : AND2_X1 port map( A1 => A(17), A2 => n14, ZN => n15);
   U16 : AND2_X1 port map( A1 => A(18), A2 => n15, ZN => n16);
   U17 : AND2_X1 port map( A1 => A(19), A2 => n16, ZN => n17);
   U18 : AND2_X1 port map( A1 => A(20), A2 => n17, ZN => n18);
   U19 : AND2_X1 port map( A1 => A(21), A2 => n18, ZN => n19);
   U20 : AND2_X1 port map( A1 => A(22), A2 => n19, ZN => n20);
   U21 : AND2_X1 port map( A1 => A(23), A2 => n20, ZN => n21);
   U22 : AND2_X1 port map( A1 => A(24), A2 => n21, ZN => n22);
   U23 : AND2_X1 port map( A1 => A(25), A2 => n22, ZN => n23);
   U24 : AND2_X1 port map( A1 => A(26), A2 => n23, ZN => n24);
   U25 : AND2_X1 port map( A1 => A(27), A2 => n24, ZN => n25);
   U26 : AND2_X1 port map( A1 => A(28), A2 => n25, ZN => n26);
   U27 : AND2_X1 port map( A1 => A(29), A2 => n26, ZN => n27);
   U28 : XOR2_X1 port map( A => A(30), B => n27, Z => SUM_30_port);
   U29 : XOR2_X1 port map( A => A(29), B => n26, Z => SUM_29_port);
   U30 : XOR2_X1 port map( A => A(28), B => n25, Z => SUM_28_port);
   U31 : XOR2_X1 port map( A => A(27), B => n24, Z => SUM_27_port);
   U32 : XOR2_X1 port map( A => A(26), B => n23, Z => SUM_26_port);
   U33 : XOR2_X1 port map( A => A(25), B => n22, Z => SUM_25_port);
   U34 : XOR2_X1 port map( A => A(24), B => n21, Z => SUM_24_port);
   U35 : XOR2_X1 port map( A => A(23), B => n20, Z => SUM_23_port);
   U36 : XOR2_X1 port map( A => A(22), B => n19, Z => SUM_22_port);
   U37 : XOR2_X1 port map( A => A(21), B => n18, Z => SUM_21_port);
   U38 : XOR2_X1 port map( A => A(20), B => n17, Z => SUM_20_port);
   U39 : XOR2_X1 port map( A => A(19), B => n16, Z => SUM_19_port);
   U40 : XOR2_X1 port map( A => A(18), B => n15, Z => SUM_18_port);
   U41 : XOR2_X1 port map( A => A(17), B => n14, Z => SUM_17_port);
   U42 : XOR2_X1 port map( A => A(16), B => n13, Z => SUM_16_port);
   U43 : XOR2_X1 port map( A => A(15), B => n12, Z => SUM_15_port);
   U44 : XOR2_X1 port map( A => A(14), B => n11, Z => SUM_14_port);
   U45 : XOR2_X1 port map( A => A(13), B => n10, Z => SUM_13_port);
   U46 : XOR2_X1 port map( A => A(12), B => n9, Z => SUM_12_port);
   U47 : XOR2_X1 port map( A => A(11), B => n8, Z => SUM_11_port);
   U48 : XOR2_X1 port map( A => A(10), B => n7, Z => SUM_10_port);
   U49 : XOR2_X1 port map( A => A(9), B => n6, Z => SUM_9_port);
   U50 : XOR2_X1 port map( A => A(8), B => n5, Z => SUM_8_port);
   U51 : XOR2_X1 port map( A => A(7), B => n4, Z => SUM_7_port);
   U52 : XOR2_X1 port map( A => A(6), B => n3, Z => SUM_6_port);
   U53 : XOR2_X1 port map( A => A(5), B => n2, Z => SUM_5_port);
   U54 : XOR2_X1 port map( A => A(4), B => n1, Z => SUM_4_port);
   U55 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U56 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U57 : XNOR2_X1 port map( A => A(31), B => n57, ZN => SUM_31_port);
   U58 : NAND2_X1 port map( A1 => A(30), A2 => n27, ZN => n57);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_6;

architecture SYN_BEHAVIORAL of MUX21_N4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_5;

architecture SYN_BEHAVIORAL of MUX21_N4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_4;

architecture SYN_BEHAVIORAL of MUX21_N4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_3;

architecture SYN_BEHAVIORAL of MUX21_N4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_2;

architecture SYN_BEHAVIORAL of MUX21_N4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_1;

architecture SYN_BEHAVIORAL of MUX21_N4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_0;

architecture SYN_BEHAVIORAL of MUX21_N4_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_BEHAVIORAL of RCA_N4_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_BEHAVIORAL of RCA_N4_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_BEHAVIORAL of RCA_N4_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_BEHAVIORAL of RCA_N4_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_BEHAVIORAL of RCA_N4_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_BEHAVIORAL of RCA_N4_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_BEHAVIORAL of RCA_N4_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_BEHAVIORAL of RCA_N4_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_BEHAVIORAL of RCA_N4_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_BEHAVIORAL of RCA_N4_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_BEHAVIORAL of RCA_N4_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_BEHAVIORAL of RCA_N4_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_BEHAVIORAL of RCA_N4_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_BEHAVIORAL of RCA_N4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_BEHAVIORAL of RCA_N4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_6 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_6;

architecture SYN_BEHAVIORAL of ENCODER_6 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : AND3_X1 port map( A1 => B(2), A2 => n1, A3 => n2, ZN => Y(2));
   U4 : INV_X1 port map( A => n3, ZN => Y(1));
   U5 : MUX2_X1 port map( A => n1, B => n2, S => B(2), Z => n3);
   U6 : AOI21_X1 port map( B1 => n2, B2 => n1, A => B(2), ZN => Y(0));
   U7 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n1);
   U8 : XNOR2_X1 port map( A => B(0), B => B(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_5 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_5;

architecture SYN_BEHAVIORAL of ENCODER_5 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : AND3_X1 port map( A1 => B(2), A2 => n1, A3 => n2, ZN => Y(2));
   U4 : INV_X1 port map( A => n3, ZN => Y(1));
   U5 : MUX2_X1 port map( A => n1, B => n2, S => B(2), Z => n3);
   U6 : AOI21_X1 port map( B1 => n2, B2 => n1, A => B(2), ZN => Y(0));
   U7 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n1);
   U8 : XNOR2_X1 port map( A => B(0), B => B(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_4 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_4;

architecture SYN_BEHAVIORAL of ENCODER_4 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : AND3_X1 port map( A1 => B(2), A2 => n1, A3 => n2, ZN => Y(2));
   U4 : INV_X1 port map( A => n3, ZN => Y(1));
   U5 : MUX2_X1 port map( A => n1, B => n2, S => B(2), Z => n3);
   U6 : AOI21_X1 port map( B1 => n2, B2 => n1, A => B(2), ZN => Y(0));
   U7 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n1);
   U8 : XNOR2_X1 port map( A => B(0), B => B(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_3 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_3;

architecture SYN_BEHAVIORAL of ENCODER_3 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : AND3_X1 port map( A1 => B(2), A2 => n1, A3 => n2, ZN => Y(2));
   U4 : INV_X1 port map( A => n3, ZN => Y(1));
   U5 : MUX2_X1 port map( A => n1, B => n2, S => B(2), Z => n3);
   U6 : AOI21_X1 port map( B1 => n2, B2 => n1, A => B(2), ZN => Y(0));
   U7 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n1);
   U8 : XNOR2_X1 port map( A => B(0), B => B(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_2 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_2;

architecture SYN_BEHAVIORAL of ENCODER_2 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : AND3_X1 port map( A1 => B(2), A2 => n1, A3 => n2, ZN => Y(2));
   U4 : INV_X1 port map( A => n3, ZN => Y(1));
   U5 : MUX2_X1 port map( A => n1, B => n2, S => B(2), Z => n3);
   U6 : AOI21_X1 port map( B1 => n2, B2 => n1, A => B(2), ZN => Y(0));
   U7 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n1);
   U8 : XNOR2_X1 port map( A => B(0), B => B(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_1 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_1;

architecture SYN_BEHAVIORAL of ENCODER_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : AND3_X1 port map( A1 => B(2), A2 => n1, A3 => n2, ZN => Y(2));
   U4 : INV_X1 port map( A => n3, ZN => Y(1));
   U5 : MUX2_X1 port map( A => n1, B => n2, S => B(2), Z => n3);
   U6 : AOI21_X1 port map( B1 => n2, B2 => n1, A => B(2), ZN => Y(0));
   U7 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n1);
   U8 : XNOR2_X1 port map( A => B(0), B => B(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_0 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_0;

architecture SYN_BEHAVIORAL of ENCODER_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : AND3_X1 port map( A1 => B(2), A2 => n1, A3 => n2, ZN => Y(2));
   U4 : INV_X1 port map( A => n3, ZN => Y(1));
   U5 : MUX2_X1 port map( A => n1, B => n2, S => B(2), Z => n3);
   U6 : AOI21_X1 port map( B1 => n2, B2 => n1, A => B(2), ZN => Y(0));
   U7 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n1);
   U8 : XNOR2_X1 port map( A => B(0), B => B(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_5;

architecture SYN_STRUCTURAL of CSB_N4_5 is

   component MUX21_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1208, 
      n_1209 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1208);
   RCA1 : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1209);
   MUX : MUX21_N4_5 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_4;

architecture SYN_STRUCTURAL of CSB_N4_4 is

   component MUX21_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1210, 
      n_1211 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1210);
   RCA1 : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1211);
   MUX : MUX21_N4_4 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_3;

architecture SYN_STRUCTURAL of CSB_N4_3 is

   component MUX21_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1212, 
      n_1213 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1212);
   RCA1 : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1213);
   MUX : MUX21_N4_3 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_2;

architecture SYN_STRUCTURAL of CSB_N4_2 is

   component MUX21_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1214, 
      n_1215 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1214);
   RCA1 : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1215);
   MUX : MUX21_N4_2 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_1;

architecture SYN_STRUCTURAL of CSB_N4_1 is

   component MUX21_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1216, 
      n_1217 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1216);
   RCA1 : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1217);
   MUX : MUX21_N4_1 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_0;

architecture SYN_STRUCTURAL of CSB_N4_0 is

   component MUX21_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1218, 
      n_1219 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1218);
   RCA1 : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1219);
   MUX : MUX21_N4_0 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_32 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_32;

architecture SYN_BEHAVIORAL of PG_BLOCK_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_31 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_31;

architecture SYN_BEHAVIORAL of PG_BLOCK_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_30 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_30;

architecture SYN_BEHAVIORAL of PG_BLOCK_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_29 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_29;

architecture SYN_BEHAVIORAL of PG_BLOCK_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_28 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_28;

architecture SYN_BEHAVIORAL of PG_BLOCK_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_27 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_27;

architecture SYN_BEHAVIORAL of PG_BLOCK_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_26 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_26;

architecture SYN_BEHAVIORAL of PG_BLOCK_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_25 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_25;

architecture SYN_BEHAVIORAL of PG_BLOCK_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_24 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_24;

architecture SYN_BEHAVIORAL of PG_BLOCK_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_23 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_23;

architecture SYN_BEHAVIORAL of PG_BLOCK_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_22 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_22;

architecture SYN_BEHAVIORAL of PG_BLOCK_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_21 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_21;

architecture SYN_BEHAVIORAL of PG_BLOCK_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_20 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_20;

architecture SYN_BEHAVIORAL of PG_BLOCK_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_19 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_19;

architecture SYN_BEHAVIORAL of PG_BLOCK_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_18 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_18;

architecture SYN_BEHAVIORAL of PG_BLOCK_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_17 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_17;

architecture SYN_BEHAVIORAL of PG_BLOCK_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_16 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_16;

architecture SYN_BEHAVIORAL of PG_BLOCK_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_15 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_15;

architecture SYN_BEHAVIORAL of PG_BLOCK_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_14 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_14;

architecture SYN_BEHAVIORAL of PG_BLOCK_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_13 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_13;

architecture SYN_BEHAVIORAL of PG_BLOCK_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_12 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_12;

architecture SYN_BEHAVIORAL of PG_BLOCK_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_11 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_11;

architecture SYN_BEHAVIORAL of PG_BLOCK_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_10 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_10;

architecture SYN_BEHAVIORAL of PG_BLOCK_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_9 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_9;

architecture SYN_BEHAVIORAL of PG_BLOCK_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_8 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_8;

architecture SYN_BEHAVIORAL of PG_BLOCK_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_7 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_7;

architecture SYN_BEHAVIORAL of PG_BLOCK_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_6 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_6;

architecture SYN_BEHAVIORAL of PG_BLOCK_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_5 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_5;

architecture SYN_BEHAVIORAL of PG_BLOCK_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_4 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_4;

architecture SYN_BEHAVIORAL of PG_BLOCK_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_3 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_3;

architecture SYN_BEHAVIORAL of PG_BLOCK_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_2 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_2;

architecture SYN_BEHAVIORAL of PG_BLOCK_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_1 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_1;

architecture SYN_BEHAVIORAL of PG_BLOCK_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_0 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_0;

architecture SYN_BEHAVIORAL of PG_BLOCK_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_7 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_7;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_6 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_6;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_5 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_5;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_4 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_4;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_3 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_3;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_2 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_2;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_1 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_1;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_0 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_0;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_N32_1;

architecture SYN_BEHAVIORAL of RCA_N32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(9));
   U2 : XOR2_X1 port map( A => B(9), B => A(9), Z => n2);
   U3 : XNOR2_X1 port map( A => n3, B => n4, ZN => S(8));
   U4 : XNOR2_X1 port map( A => A(8), B => B(8), ZN => n4);
   U5 : XOR2_X1 port map( A => n5, B => n6, Z => S(7));
   U6 : XNOR2_X1 port map( A => B(7), B => n7, ZN => n6);
   U7 : XNOR2_X1 port map( A => n8, B => n9, ZN => S(6));
   U8 : XNOR2_X1 port map( A => A(6), B => B(6), ZN => n9);
   U9 : XOR2_X1 port map( A => n10, B => n11, Z => S(5));
   U10 : XOR2_X1 port map( A => B(5), B => A(5), Z => n11);
   U11 : XNOR2_X1 port map( A => n12, B => n13, ZN => S(4));
   U12 : XNOR2_X1 port map( A => A(4), B => B(4), ZN => n13);
   U13 : XNOR2_X1 port map( A => n14, B => n15, ZN => S(3));
   U14 : XNOR2_X1 port map( A => B(3), B => n16, ZN => n15);
   U15 : XOR2_X1 port map( A => n17, B => n18, Z => S(31));
   U16 : XOR2_X1 port map( A => B(31), B => A(31), Z => n18);
   U17 : XNOR2_X1 port map( A => n19, B => n20, ZN => S(30));
   U18 : XNOR2_X1 port map( A => B(30), B => n21, ZN => n20);
   U19 : XNOR2_X1 port map( A => n22, B => n23, ZN => S(2));
   U20 : XOR2_X1 port map( A => B(2), B => A(2), Z => n23);
   U21 : XOR2_X1 port map( A => n24, B => n25, Z => S(29));
   U22 : XOR2_X1 port map( A => B(29), B => A(29), Z => n25);
   U23 : XNOR2_X1 port map( A => n26, B => n27, ZN => S(28));
   U24 : XNOR2_X1 port map( A => B(28), B => n28, ZN => n27);
   U25 : XNOR2_X1 port map( A => n29, B => n30, ZN => S(27));
   U26 : XOR2_X1 port map( A => B(27), B => A(27), Z => n30);
   U27 : XOR2_X1 port map( A => n31, B => n32, Z => S(26));
   U28 : XOR2_X1 port map( A => B(26), B => A(26), Z => n32);
   U29 : XNOR2_X1 port map( A => n33, B => n34, ZN => S(25));
   U30 : XNOR2_X1 port map( A => B(25), B => n35, ZN => n34);
   U31 : XOR2_X1 port map( A => n36, B => n37, Z => S(24));
   U32 : XOR2_X1 port map( A => B(24), B => A(24), Z => n37);
   U33 : XNOR2_X1 port map( A => n38, B => n39, ZN => S(23));
   U34 : XNOR2_X1 port map( A => B(23), B => n40, ZN => n39);
   U35 : XOR2_X1 port map( A => n41, B => n42, Z => S(22));
   U36 : XOR2_X1 port map( A => B(22), B => A(22), Z => n42);
   U37 : XNOR2_X1 port map( A => n43, B => n44, ZN => S(21));
   U38 : XNOR2_X1 port map( A => B(21), B => n45, ZN => n44);
   U39 : XOR2_X1 port map( A => n46, B => n47, Z => S(20));
   U40 : XOR2_X1 port map( A => B(20), B => A(20), Z => n47);
   U41 : XNOR2_X1 port map( A => n48, B => n49, ZN => S(1));
   U42 : XOR2_X1 port map( A => B(1), B => A(1), Z => n49);
   U43 : XNOR2_X1 port map( A => n50, B => n51, ZN => S(19));
   U44 : XNOR2_X1 port map( A => B(19), B => n52, ZN => n51);
   U45 : XNOR2_X1 port map( A => n53, B => n54, ZN => S(18));
   U46 : XNOR2_X1 port map( A => B(18), B => n55, ZN => n54);
   U47 : XOR2_X1 port map( A => n56, B => n57, Z => S(17));
   U48 : XOR2_X1 port map( A => B(17), B => A(17), Z => n57);
   U49 : XNOR2_X1 port map( A => n58, B => n59, ZN => S(16));
   U50 : XNOR2_X1 port map( A => B(16), B => n60, ZN => n59);
   U51 : XOR2_X1 port map( A => n61, B => n62, Z => S(15));
   U52 : XOR2_X1 port map( A => B(15), B => A(15), Z => n62);
   U53 : XNOR2_X1 port map( A => n63, B => n64, ZN => S(14));
   U54 : XOR2_X1 port map( A => B(14), B => A(14), Z => n64);
   U55 : XOR2_X1 port map( A => n65, B => n66, Z => S(13));
   U56 : XOR2_X1 port map( A => B(13), B => A(13), Z => n66);
   U57 : XNOR2_X1 port map( A => n67, B => n68, ZN => S(12));
   U58 : XNOR2_X1 port map( A => A(12), B => B(12), ZN => n68);
   U59 : XOR2_X1 port map( A => n69, B => n70, Z => S(11));
   U60 : XOR2_X1 port map( A => B(11), B => A(11), Z => n70);
   U61 : XNOR2_X1 port map( A => n71, B => n72, ZN => S(10));
   U62 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => n72);
   U63 : XOR2_X1 port map( A => A(0), B => n73, Z => S(0));
   U64 : XOR2_X1 port map( A => Ci, B => B(0), Z => n73);
   U65 : INV_X1 port map( A => n74, ZN => Co);
   U66 : AOI22_X1 port map( A1 => A(31), A2 => n17, B1 => n75, B2 => B(31), ZN 
                           => n74);
   U67 : OR2_X1 port map( A1 => n17, A2 => A(31), ZN => n75);
   U68 : AOI21_X1 port map( B1 => n21, B2 => n19, A => n76, ZN => n17);
   U69 : AOI21_X1 port map( B1 => n77, B2 => A(30), A => B(30), ZN => n76);
   U70 : INV_X1 port map( A => n19, ZN => n77);
   U71 : AOI22_X1 port map( A1 => n24, A2 => A(29), B1 => n78, B2 => B(29), ZN 
                           => n19);
   U72 : OR2_X1 port map( A1 => A(29), A2 => n24, ZN => n78);
   U73 : OAI21_X1 port map( B1 => n26, B2 => n28, A => n79, ZN => n24);
   U74 : OAI21_X1 port map( B1 => n80, B2 => A(28), A => B(28), ZN => n79);
   U75 : INV_X1 port map( A => n26, ZN => n80);
   U76 : INV_X1 port map( A => A(28), ZN => n28);
   U77 : OAI21_X1 port map( B1 => A(27), B2 => n81, A => n82, ZN => n26);
   U78 : INV_X1 port map( A => n83, ZN => n82);
   U79 : AOI21_X1 port map( B1 => n81, B2 => A(27), A => B(27), ZN => n83);
   U80 : INV_X1 port map( A => n29, ZN => n81);
   U81 : AOI22_X1 port map( A1 => n31, A2 => A(26), B1 => n84, B2 => B(26), ZN 
                           => n29);
   U82 : OR2_X1 port map( A1 => n31, A2 => A(26), ZN => n84);
   U83 : AOI21_X1 port map( B1 => n35, B2 => n33, A => n85, ZN => n31);
   U84 : AOI21_X1 port map( B1 => n86, B2 => A(25), A => B(25), ZN => n85);
   U85 : INV_X1 port map( A => n33, ZN => n86);
   U86 : AOI21_X1 port map( B1 => n36, B2 => A(24), A => n87, ZN => n33);
   U87 : INV_X1 port map( A => n88, ZN => n87);
   U88 : OAI21_X1 port map( B1 => n36, B2 => A(24), A => B(24), ZN => n88);
   U89 : AOI21_X1 port map( B1 => n40, B2 => n38, A => n89, ZN => n36);
   U90 : AOI21_X1 port map( B1 => n90, B2 => A(23), A => B(23), ZN => n89);
   U91 : INV_X1 port map( A => n38, ZN => n90);
   U92 : AOI21_X1 port map( B1 => n41, B2 => A(22), A => n91, ZN => n38);
   U93 : INV_X1 port map( A => n92, ZN => n91);
   U94 : OAI21_X1 port map( B1 => n41, B2 => A(22), A => B(22), ZN => n92);
   U95 : AOI21_X1 port map( B1 => n45, B2 => n43, A => n93, ZN => n41);
   U96 : AOI21_X1 port map( B1 => n94, B2 => A(21), A => B(21), ZN => n93);
   U97 : INV_X1 port map( A => n43, ZN => n94);
   U98 : AOI22_X1 port map( A1 => n46, A2 => A(20), B1 => n95, B2 => B(20), ZN 
                           => n43);
   U99 : OR2_X1 port map( A1 => n46, A2 => A(20), ZN => n95);
   U100 : AOI21_X1 port map( B1 => n52, B2 => n50, A => n96, ZN => n46);
   U101 : AOI21_X1 port map( B1 => n97, B2 => A(19), A => B(19), ZN => n96);
   U102 : INV_X1 port map( A => n97, ZN => n50);
   U103 : OAI21_X1 port map( B1 => n53, B2 => n55, A => n98, ZN => n97);
   U104 : OAI21_X1 port map( B1 => n99, B2 => A(18), A => B(18), ZN => n98);
   U105 : INV_X1 port map( A => n53, ZN => n99);
   U106 : INV_X1 port map( A => A(18), ZN => n55);
   U107 : OAI21_X1 port map( B1 => A(17), B2 => n56, A => n100, ZN => n53);
   U108 : INV_X1 port map( A => n101, ZN => n100);
   U109 : AOI21_X1 port map( B1 => n56, B2 => A(17), A => B(17), ZN => n101);
   U110 : OAI21_X1 port map( B1 => n58, B2 => n60, A => n102, ZN => n56);
   U111 : OAI21_X1 port map( B1 => n103, B2 => A(16), A => B(16), ZN => n102);
   U112 : INV_X1 port map( A => n58, ZN => n103);
   U113 : INV_X1 port map( A => A(16), ZN => n60);
   U114 : OAI21_X1 port map( B1 => A(15), B2 => n61, A => n104, ZN => n58);
   U115 : INV_X1 port map( A => n105, ZN => n104);
   U116 : AOI21_X1 port map( B1 => n61, B2 => A(15), A => B(15), ZN => n105);
   U117 : OAI21_X1 port map( B1 => n63, B2 => n106, A => n107, ZN => n61);
   U118 : OAI21_X1 port map( B1 => n108, B2 => A(14), A => B(14), ZN => n107);
   U119 : INV_X1 port map( A => n63, ZN => n108);
   U120 : INV_X1 port map( A => A(14), ZN => n106);
   U121 : OAI21_X1 port map( B1 => A(13), B2 => n65, A => n109, ZN => n63);
   U122 : INV_X1 port map( A => n110, ZN => n109);
   U123 : AOI21_X1 port map( B1 => n65, B2 => A(13), A => B(13), ZN => n110);
   U124 : OAI21_X1 port map( B1 => n111, B2 => n112, A => n113, ZN => n65);
   U125 : OAI21_X1 port map( B1 => n67, B2 => A(12), A => B(12), ZN => n113);
   U126 : INV_X1 port map( A => n111, ZN => n67);
   U127 : INV_X1 port map( A => A(12), ZN => n112);
   U128 : OAI21_X1 port map( B1 => A(11), B2 => n69, A => n114, ZN => n111);
   U129 : INV_X1 port map( A => n115, ZN => n114);
   U130 : AOI21_X1 port map( B1 => n69, B2 => A(11), A => B(11), ZN => n115);
   U131 : OAI21_X1 port map( B1 => n116, B2 => n117, A => n118, ZN => n69);
   U132 : OAI21_X1 port map( B1 => n71, B2 => A(10), A => B(10), ZN => n118);
   U133 : INV_X1 port map( A => A(10), ZN => n117);
   U134 : INV_X1 port map( A => n71, ZN => n116);
   U135 : AOI21_X1 port map( B1 => n119, B2 => n1, A => n120, ZN => n71);
   U136 : AOI21_X1 port map( B1 => n121, B2 => A(9), A => B(9), ZN => n120);
   U137 : INV_X1 port map( A => n1, ZN => n121);
   U138 : AOI21_X1 port map( B1 => n3, B2 => A(8), A => n122, ZN => n1);
   U139 : INV_X1 port map( A => n123, ZN => n122);
   U140 : OAI21_X1 port map( B1 => n3, B2 => A(8), A => B(8), ZN => n123);
   U141 : AOI21_X1 port map( B1 => n7, B2 => n124, A => n125, ZN => n3);
   U142 : AOI21_X1 port map( B1 => n5, B2 => A(7), A => B(7), ZN => n125);
   U143 : INV_X1 port map( A => n124, ZN => n5);
   U144 : AOI21_X1 port map( B1 => n8, B2 => A(6), A => n126, ZN => n124);
   U145 : INV_X1 port map( A => n127, ZN => n126);
   U146 : OAI21_X1 port map( B1 => n8, B2 => A(6), A => B(6), ZN => n127);
   U147 : AOI21_X1 port map( B1 => n128, B2 => n129, A => n130, ZN => n8);
   U148 : AOI21_X1 port map( B1 => n10, B2 => A(5), A => B(5), ZN => n130);
   U149 : INV_X1 port map( A => n129, ZN => n10);
   U150 : AOI21_X1 port map( B1 => n12, B2 => A(4), A => n131, ZN => n129);
   U151 : INV_X1 port map( A => n132, ZN => n131);
   U152 : OAI21_X1 port map( B1 => n12, B2 => A(4), A => B(4), ZN => n132);
   U153 : AOI21_X1 port map( B1 => n16, B2 => n14, A => n133, ZN => n12);
   U154 : AOI21_X1 port map( B1 => n134, B2 => A(3), A => B(3), ZN => n133);
   U155 : INV_X1 port map( A => n14, ZN => n134);
   U156 : OAI22_X1 port map( A1 => A(2), A2 => n135, B1 => B(2), B2 => n136, ZN
                           => n14);
   U157 : AND2_X1 port map( A1 => n135, A2 => A(2), ZN => n136);
   U158 : INV_X1 port map( A => n22, ZN => n135);
   U159 : OAI22_X1 port map( A1 => A(1), A2 => n137, B1 => B(1), B2 => n138, ZN
                           => n22);
   U160 : AND2_X1 port map( A1 => n137, A2 => A(1), ZN => n138);
   U161 : INV_X1 port map( A => n48, ZN => n137);
   U162 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n139, ZN => n48);
   U163 : INV_X1 port map( A => n140, ZN => n139);
   U164 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n140);
   U165 : INV_X1 port map( A => A(3), ZN => n16);
   U166 : INV_X1 port map( A => A(5), ZN => n128);
   U167 : INV_X1 port map( A => A(7), ZN => n7);
   U168 : INV_X1 port map( A => A(9), ZN => n119);
   U169 : INV_X1 port map( A => A(19), ZN => n52);
   U170 : INV_X1 port map( A => A(21), ZN => n45);
   U171 : INV_X1 port map( A => A(23), ZN => n40);
   U172 : INV_X1 port map( A => A(25), ZN => n35);
   U173 : INV_X1 port map( A => A(30), ZN => n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_N32_0;

architecture SYN_BEHAVIORAL of RCA_N32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(9));
   U2 : XOR2_X1 port map( A => B(9), B => A(9), Z => n2);
   U3 : XNOR2_X1 port map( A => n3, B => n4, ZN => S(8));
   U4 : XNOR2_X1 port map( A => A(8), B => B(8), ZN => n4);
   U5 : XOR2_X1 port map( A => n5, B => n6, Z => S(7));
   U6 : XNOR2_X1 port map( A => B(7), B => n7, ZN => n6);
   U7 : XNOR2_X1 port map( A => n8, B => n9, ZN => S(6));
   U8 : XNOR2_X1 port map( A => A(6), B => B(6), ZN => n9);
   U9 : XOR2_X1 port map( A => n10, B => n11, Z => S(5));
   U10 : XOR2_X1 port map( A => B(5), B => A(5), Z => n11);
   U11 : XNOR2_X1 port map( A => n12, B => n13, ZN => S(4));
   U12 : XNOR2_X1 port map( A => A(4), B => B(4), ZN => n13);
   U13 : XNOR2_X1 port map( A => n14, B => n15, ZN => S(3));
   U14 : XNOR2_X1 port map( A => B(3), B => n16, ZN => n15);
   U15 : XOR2_X1 port map( A => n17, B => n18, Z => S(31));
   U16 : XOR2_X1 port map( A => B(31), B => A(31), Z => n18);
   U17 : XNOR2_X1 port map( A => n19, B => n20, ZN => S(30));
   U18 : XNOR2_X1 port map( A => B(30), B => n21, ZN => n20);
   U19 : XNOR2_X1 port map( A => n22, B => n23, ZN => S(2));
   U20 : XOR2_X1 port map( A => B(2), B => A(2), Z => n23);
   U21 : XOR2_X1 port map( A => n24, B => n25, Z => S(29));
   U22 : XOR2_X1 port map( A => B(29), B => A(29), Z => n25);
   U23 : XNOR2_X1 port map( A => n26, B => n27, ZN => S(28));
   U24 : XNOR2_X1 port map( A => B(28), B => n28, ZN => n27);
   U25 : XNOR2_X1 port map( A => n29, B => n30, ZN => S(27));
   U26 : XOR2_X1 port map( A => B(27), B => A(27), Z => n30);
   U27 : XOR2_X1 port map( A => n31, B => n32, Z => S(26));
   U28 : XOR2_X1 port map( A => B(26), B => A(26), Z => n32);
   U29 : XNOR2_X1 port map( A => n33, B => n34, ZN => S(25));
   U30 : XNOR2_X1 port map( A => B(25), B => n35, ZN => n34);
   U31 : XOR2_X1 port map( A => n36, B => n37, Z => S(24));
   U32 : XOR2_X1 port map( A => B(24), B => A(24), Z => n37);
   U33 : XNOR2_X1 port map( A => n38, B => n39, ZN => S(23));
   U34 : XNOR2_X1 port map( A => B(23), B => n40, ZN => n39);
   U35 : XOR2_X1 port map( A => n41, B => n42, Z => S(22));
   U36 : XOR2_X1 port map( A => B(22), B => A(22), Z => n42);
   U37 : XNOR2_X1 port map( A => n43, B => n44, ZN => S(21));
   U38 : XNOR2_X1 port map( A => B(21), B => n45, ZN => n44);
   U39 : XOR2_X1 port map( A => n46, B => n47, Z => S(20));
   U40 : XOR2_X1 port map( A => B(20), B => A(20), Z => n47);
   U41 : XNOR2_X1 port map( A => n48, B => n49, ZN => S(1));
   U42 : XOR2_X1 port map( A => B(1), B => A(1), Z => n49);
   U43 : XNOR2_X1 port map( A => n50, B => n51, ZN => S(19));
   U44 : XNOR2_X1 port map( A => B(19), B => n52, ZN => n51);
   U45 : XNOR2_X1 port map( A => n53, B => n54, ZN => S(18));
   U46 : XNOR2_X1 port map( A => B(18), B => n55, ZN => n54);
   U47 : XOR2_X1 port map( A => n56, B => n57, Z => S(17));
   U48 : XOR2_X1 port map( A => B(17), B => A(17), Z => n57);
   U49 : XNOR2_X1 port map( A => n58, B => n59, ZN => S(16));
   U50 : XNOR2_X1 port map( A => B(16), B => n60, ZN => n59);
   U51 : XOR2_X1 port map( A => n61, B => n62, Z => S(15));
   U52 : XOR2_X1 port map( A => B(15), B => A(15), Z => n62);
   U53 : XNOR2_X1 port map( A => n63, B => n64, ZN => S(14));
   U54 : XOR2_X1 port map( A => B(14), B => A(14), Z => n64);
   U55 : XOR2_X1 port map( A => n65, B => n66, Z => S(13));
   U56 : XOR2_X1 port map( A => B(13), B => A(13), Z => n66);
   U57 : XNOR2_X1 port map( A => n67, B => n68, ZN => S(12));
   U58 : XNOR2_X1 port map( A => A(12), B => B(12), ZN => n68);
   U59 : XOR2_X1 port map( A => n69, B => n70, Z => S(11));
   U60 : XOR2_X1 port map( A => B(11), B => A(11), Z => n70);
   U61 : XNOR2_X1 port map( A => n71, B => n72, ZN => S(10));
   U62 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => n72);
   U63 : XOR2_X1 port map( A => A(0), B => n73, Z => S(0));
   U64 : XOR2_X1 port map( A => Ci, B => B(0), Z => n73);
   U65 : INV_X1 port map( A => n74, ZN => Co);
   U66 : AOI22_X1 port map( A1 => A(31), A2 => n17, B1 => n75, B2 => B(31), ZN 
                           => n74);
   U67 : OR2_X1 port map( A1 => n17, A2 => A(31), ZN => n75);
   U68 : AOI21_X1 port map( B1 => n21, B2 => n19, A => n76, ZN => n17);
   U69 : AOI21_X1 port map( B1 => n77, B2 => A(30), A => B(30), ZN => n76);
   U70 : INV_X1 port map( A => n19, ZN => n77);
   U71 : AOI22_X1 port map( A1 => n24, A2 => A(29), B1 => n78, B2 => B(29), ZN 
                           => n19);
   U72 : OR2_X1 port map( A1 => A(29), A2 => n24, ZN => n78);
   U73 : OAI21_X1 port map( B1 => n26, B2 => n28, A => n79, ZN => n24);
   U74 : OAI21_X1 port map( B1 => n80, B2 => A(28), A => B(28), ZN => n79);
   U75 : INV_X1 port map( A => n26, ZN => n80);
   U76 : INV_X1 port map( A => A(28), ZN => n28);
   U77 : OAI21_X1 port map( B1 => A(27), B2 => n81, A => n82, ZN => n26);
   U78 : INV_X1 port map( A => n83, ZN => n82);
   U79 : AOI21_X1 port map( B1 => n81, B2 => A(27), A => B(27), ZN => n83);
   U80 : INV_X1 port map( A => n29, ZN => n81);
   U81 : AOI22_X1 port map( A1 => n31, A2 => A(26), B1 => n84, B2 => B(26), ZN 
                           => n29);
   U82 : OR2_X1 port map( A1 => n31, A2 => A(26), ZN => n84);
   U83 : AOI21_X1 port map( B1 => n35, B2 => n33, A => n85, ZN => n31);
   U84 : AOI21_X1 port map( B1 => n86, B2 => A(25), A => B(25), ZN => n85);
   U85 : INV_X1 port map( A => n33, ZN => n86);
   U86 : AOI21_X1 port map( B1 => n36, B2 => A(24), A => n87, ZN => n33);
   U87 : INV_X1 port map( A => n88, ZN => n87);
   U88 : OAI21_X1 port map( B1 => n36, B2 => A(24), A => B(24), ZN => n88);
   U89 : AOI21_X1 port map( B1 => n40, B2 => n38, A => n89, ZN => n36);
   U90 : AOI21_X1 port map( B1 => n90, B2 => A(23), A => B(23), ZN => n89);
   U91 : INV_X1 port map( A => n38, ZN => n90);
   U92 : AOI21_X1 port map( B1 => n41, B2 => A(22), A => n91, ZN => n38);
   U93 : INV_X1 port map( A => n92, ZN => n91);
   U94 : OAI21_X1 port map( B1 => n41, B2 => A(22), A => B(22), ZN => n92);
   U95 : AOI21_X1 port map( B1 => n45, B2 => n43, A => n93, ZN => n41);
   U96 : AOI21_X1 port map( B1 => n94, B2 => A(21), A => B(21), ZN => n93);
   U97 : INV_X1 port map( A => n43, ZN => n94);
   U98 : AOI22_X1 port map( A1 => n46, A2 => A(20), B1 => n95, B2 => B(20), ZN 
                           => n43);
   U99 : OR2_X1 port map( A1 => n46, A2 => A(20), ZN => n95);
   U100 : AOI21_X1 port map( B1 => n52, B2 => n50, A => n96, ZN => n46);
   U101 : AOI21_X1 port map( B1 => n97, B2 => A(19), A => B(19), ZN => n96);
   U102 : INV_X1 port map( A => n97, ZN => n50);
   U103 : OAI21_X1 port map( B1 => n53, B2 => n55, A => n98, ZN => n97);
   U104 : OAI21_X1 port map( B1 => n99, B2 => A(18), A => B(18), ZN => n98);
   U105 : INV_X1 port map( A => n53, ZN => n99);
   U106 : INV_X1 port map( A => A(18), ZN => n55);
   U107 : OAI21_X1 port map( B1 => A(17), B2 => n56, A => n100, ZN => n53);
   U108 : INV_X1 port map( A => n101, ZN => n100);
   U109 : AOI21_X1 port map( B1 => n56, B2 => A(17), A => B(17), ZN => n101);
   U110 : OAI21_X1 port map( B1 => n58, B2 => n60, A => n102, ZN => n56);
   U111 : OAI21_X1 port map( B1 => n103, B2 => A(16), A => B(16), ZN => n102);
   U112 : INV_X1 port map( A => n58, ZN => n103);
   U113 : INV_X1 port map( A => A(16), ZN => n60);
   U114 : OAI21_X1 port map( B1 => A(15), B2 => n61, A => n104, ZN => n58);
   U115 : INV_X1 port map( A => n105, ZN => n104);
   U116 : AOI21_X1 port map( B1 => n61, B2 => A(15), A => B(15), ZN => n105);
   U117 : OAI21_X1 port map( B1 => n63, B2 => n106, A => n107, ZN => n61);
   U118 : OAI21_X1 port map( B1 => n108, B2 => A(14), A => B(14), ZN => n107);
   U119 : INV_X1 port map( A => n63, ZN => n108);
   U120 : INV_X1 port map( A => A(14), ZN => n106);
   U121 : OAI21_X1 port map( B1 => A(13), B2 => n65, A => n109, ZN => n63);
   U122 : INV_X1 port map( A => n110, ZN => n109);
   U123 : AOI21_X1 port map( B1 => n65, B2 => A(13), A => B(13), ZN => n110);
   U124 : OAI21_X1 port map( B1 => n111, B2 => n112, A => n113, ZN => n65);
   U125 : OAI21_X1 port map( B1 => n67, B2 => A(12), A => B(12), ZN => n113);
   U126 : INV_X1 port map( A => n111, ZN => n67);
   U127 : INV_X1 port map( A => A(12), ZN => n112);
   U128 : OAI21_X1 port map( B1 => A(11), B2 => n69, A => n114, ZN => n111);
   U129 : INV_X1 port map( A => n115, ZN => n114);
   U130 : AOI21_X1 port map( B1 => n69, B2 => A(11), A => B(11), ZN => n115);
   U131 : OAI21_X1 port map( B1 => n116, B2 => n117, A => n118, ZN => n69);
   U132 : OAI21_X1 port map( B1 => n71, B2 => A(10), A => B(10), ZN => n118);
   U133 : INV_X1 port map( A => A(10), ZN => n117);
   U134 : INV_X1 port map( A => n71, ZN => n116);
   U135 : AOI21_X1 port map( B1 => n119, B2 => n1, A => n120, ZN => n71);
   U136 : AOI21_X1 port map( B1 => n121, B2 => A(9), A => B(9), ZN => n120);
   U137 : INV_X1 port map( A => n1, ZN => n121);
   U138 : AOI21_X1 port map( B1 => n3, B2 => A(8), A => n122, ZN => n1);
   U139 : INV_X1 port map( A => n123, ZN => n122);
   U140 : OAI21_X1 port map( B1 => n3, B2 => A(8), A => B(8), ZN => n123);
   U141 : AOI21_X1 port map( B1 => n7, B2 => n124, A => n125, ZN => n3);
   U142 : AOI21_X1 port map( B1 => n5, B2 => A(7), A => B(7), ZN => n125);
   U143 : INV_X1 port map( A => n124, ZN => n5);
   U144 : AOI21_X1 port map( B1 => n8, B2 => A(6), A => n126, ZN => n124);
   U145 : INV_X1 port map( A => n127, ZN => n126);
   U146 : OAI21_X1 port map( B1 => n8, B2 => A(6), A => B(6), ZN => n127);
   U147 : AOI21_X1 port map( B1 => n128, B2 => n129, A => n130, ZN => n8);
   U148 : AOI21_X1 port map( B1 => n10, B2 => A(5), A => B(5), ZN => n130);
   U149 : INV_X1 port map( A => n129, ZN => n10);
   U150 : AOI21_X1 port map( B1 => n12, B2 => A(4), A => n131, ZN => n129);
   U151 : INV_X1 port map( A => n132, ZN => n131);
   U152 : OAI21_X1 port map( B1 => n12, B2 => A(4), A => B(4), ZN => n132);
   U153 : AOI21_X1 port map( B1 => n16, B2 => n14, A => n133, ZN => n12);
   U154 : AOI21_X1 port map( B1 => n134, B2 => A(3), A => B(3), ZN => n133);
   U155 : INV_X1 port map( A => n14, ZN => n134);
   U156 : OAI22_X1 port map( A1 => A(2), A2 => n135, B1 => B(2), B2 => n136, ZN
                           => n14);
   U157 : AND2_X1 port map( A1 => n135, A2 => A(2), ZN => n136);
   U158 : INV_X1 port map( A => n22, ZN => n135);
   U159 : OAI22_X1 port map( A1 => A(1), A2 => n137, B1 => B(1), B2 => n138, ZN
                           => n22);
   U160 : AND2_X1 port map( A1 => n137, A2 => A(1), ZN => n138);
   U161 : INV_X1 port map( A => n48, ZN => n137);
   U162 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n139, ZN => n48);
   U163 : INV_X1 port map( A => n140, ZN => n139);
   U164 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n140);
   U165 : INV_X1 port map( A => A(3), ZN => n16);
   U166 : INV_X1 port map( A => A(5), ZN => n128);
   U167 : INV_X1 port map( A => A(7), ZN => n7);
   U168 : INV_X1 port map( A => A(9), ZN => n119);
   U169 : INV_X1 port map( A => A(19), ZN => n52);
   U170 : INV_X1 port map( A => A(21), ZN => n45);
   U171 : INV_X1 port map( A => A(23), ZN => n40);
   U172 : INV_X1 port map( A => A(25), ZN => n35);
   U173 : INV_X1 port map( A => A(30), ZN => n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX81_N32_2 is

   port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX81_N32_2;

architecture SYN_BEHAVIORAL of MUX81_N32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142 : std_logic;

begin
   
   U1 : OR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n142, ZN => n1);
   U2 : OR3_X1 port map( A1 => S(1), A2 => S(2), A3 => S(0), ZN => n2);
   U3 : OR3_X1 port map( A1 => n142, A2 => S(2), A3 => n141, ZN => n3);
   U4 : OR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n141, ZN => n4);
   U5 : AND3_X2 port map( A1 => S(2), A2 => S(1), A3 => S(0), ZN => n14);
   U6 : AND3_X2 port map( A1 => S(2), A2 => n142, A3 => S(0), ZN => n16);
   U7 : AND3_X2 port map( A1 => S(1), A2 => n141, A3 => S(2), ZN => n13);
   U8 : AND3_X2 port map( A1 => n141, A2 => n142, A3 => S(2), ZN => n15);
   U9 : INV_X2 port map( A => n3, ZN => n5);
   U10 : INV_X2 port map( A => n4, ZN => n6);
   U11 : INV_X2 port map( A => n1, ZN => n7);
   U12 : INV_X2 port map( A => n2, ZN => n8);
   U13 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => 
                           Y(9));
   U14 : AOI22_X1 port map( A1 => G(9), A2 => n13, B1 => H(9), B2 => n14, ZN =>
                           n12);
   U15 : AOI22_X1 port map( A1 => E(9), A2 => n15, B1 => F(9), B2 => n16, ZN =>
                           n11);
   U16 : AOI22_X1 port map( A1 => C(9), A2 => n7, B1 => D(9), B2 => n5, ZN => 
                           n10);
   U17 : AOI22_X1 port map( A1 => A(9), A2 => n8, B1 => B(9), B2 => n6, ZN => 
                           n9);
   U18 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           Y(8));
   U19 : AOI22_X1 port map( A1 => G(8), A2 => n13, B1 => H(8), B2 => n14, ZN =>
                           n20);
   U20 : AOI22_X1 port map( A1 => E(8), A2 => n15, B1 => F(8), B2 => n16, ZN =>
                           n19);
   U21 : AOI22_X1 port map( A1 => C(8), A2 => n7, B1 => D(8), B2 => n5, ZN => 
                           n18);
   U22 : AOI22_X1 port map( A1 => A(8), A2 => n8, B1 => B(8), B2 => n6, ZN => 
                           n17);
   U23 : NAND4_X1 port map( A1 => n21, A2 => n22, A3 => n23, A4 => n24, ZN => 
                           Y(7));
   U24 : AOI22_X1 port map( A1 => G(7), A2 => n13, B1 => H(7), B2 => n14, ZN =>
                           n24);
   U25 : AOI22_X1 port map( A1 => E(7), A2 => n15, B1 => F(7), B2 => n16, ZN =>
                           n23);
   U26 : AOI22_X1 port map( A1 => C(7), A2 => n7, B1 => D(7), B2 => n5, ZN => 
                           n22);
   U27 : AOI22_X1 port map( A1 => A(7), A2 => n8, B1 => B(7), B2 => n6, ZN => 
                           n21);
   U28 : NAND4_X1 port map( A1 => n25, A2 => n26, A3 => n27, A4 => n28, ZN => 
                           Y(6));
   U29 : AOI22_X1 port map( A1 => G(6), A2 => n13, B1 => H(6), B2 => n14, ZN =>
                           n28);
   U30 : AOI22_X1 port map( A1 => E(6), A2 => n15, B1 => F(6), B2 => n16, ZN =>
                           n27);
   U31 : AOI22_X1 port map( A1 => C(6), A2 => n7, B1 => D(6), B2 => n5, ZN => 
                           n26);
   U32 : AOI22_X1 port map( A1 => A(6), A2 => n8, B1 => B(6), B2 => n6, ZN => 
                           n25);
   U33 : NAND4_X1 port map( A1 => n29, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           Y(5));
   U34 : AOI22_X1 port map( A1 => G(5), A2 => n13, B1 => H(5), B2 => n14, ZN =>
                           n32);
   U35 : AOI22_X1 port map( A1 => E(5), A2 => n15, B1 => F(5), B2 => n16, ZN =>
                           n31);
   U36 : AOI22_X1 port map( A1 => C(5), A2 => n7, B1 => D(5), B2 => n5, ZN => 
                           n30);
   U37 : AOI22_X1 port map( A1 => A(5), A2 => n8, B1 => B(5), B2 => n6, ZN => 
                           n29);
   U38 : NAND4_X1 port map( A1 => n33, A2 => n34, A3 => n35, A4 => n36, ZN => 
                           Y(4));
   U39 : AOI22_X1 port map( A1 => G(4), A2 => n13, B1 => H(4), B2 => n14, ZN =>
                           n36);
   U40 : AOI22_X1 port map( A1 => E(4), A2 => n15, B1 => F(4), B2 => n16, ZN =>
                           n35);
   U41 : AOI22_X1 port map( A1 => C(4), A2 => n7, B1 => D(4), B2 => n5, ZN => 
                           n34);
   U42 : AOI22_X1 port map( A1 => A(4), A2 => n8, B1 => B(4), B2 => n6, ZN => 
                           n33);
   U43 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           Y(3));
   U44 : AOI22_X1 port map( A1 => G(3), A2 => n13, B1 => H(3), B2 => n14, ZN =>
                           n40);
   U45 : AOI22_X1 port map( A1 => E(3), A2 => n15, B1 => F(3), B2 => n16, ZN =>
                           n39);
   U46 : AOI22_X1 port map( A1 => C(3), A2 => n7, B1 => D(3), B2 => n5, ZN => 
                           n38);
   U47 : AOI22_X1 port map( A1 => A(3), A2 => n8, B1 => B(3), B2 => n6, ZN => 
                           n37);
   U48 : NAND4_X1 port map( A1 => n41, A2 => n42, A3 => n43, A4 => n44, ZN => 
                           Y(31));
   U49 : AOI22_X1 port map( A1 => G(31), A2 => n13, B1 => H(31), B2 => n14, ZN 
                           => n44);
   U50 : AOI22_X1 port map( A1 => E(31), A2 => n15, B1 => F(31), B2 => n16, ZN 
                           => n43);
   U51 : AOI22_X1 port map( A1 => C(31), A2 => n7, B1 => D(31), B2 => n5, ZN =>
                           n42);
   U52 : AOI22_X1 port map( A1 => A(31), A2 => n8, B1 => B(31), B2 => n6, ZN =>
                           n41);
   U53 : NAND4_X1 port map( A1 => n45, A2 => n46, A3 => n47, A4 => n48, ZN => 
                           Y(30));
   U54 : AOI22_X1 port map( A1 => G(30), A2 => n13, B1 => H(30), B2 => n14, ZN 
                           => n48);
   U55 : AOI22_X1 port map( A1 => E(30), A2 => n15, B1 => F(30), B2 => n16, ZN 
                           => n47);
   U56 : AOI22_X1 port map( A1 => C(30), A2 => n7, B1 => D(30), B2 => n5, ZN =>
                           n46);
   U57 : AOI22_X1 port map( A1 => A(30), A2 => n8, B1 => B(30), B2 => n6, ZN =>
                           n45);
   U58 : NAND4_X1 port map( A1 => n49, A2 => n50, A3 => n51, A4 => n52, ZN => 
                           Y(2));
   U59 : AOI22_X1 port map( A1 => G(2), A2 => n13, B1 => H(2), B2 => n14, ZN =>
                           n52);
   U60 : AOI22_X1 port map( A1 => E(2), A2 => n15, B1 => F(2), B2 => n16, ZN =>
                           n51);
   U61 : AOI22_X1 port map( A1 => C(2), A2 => n7, B1 => D(2), B2 => n5, ZN => 
                           n50);
   U62 : AOI22_X1 port map( A1 => A(2), A2 => n8, B1 => B(2), B2 => n6, ZN => 
                           n49);
   U63 : NAND4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           Y(29));
   U64 : AOI22_X1 port map( A1 => G(29), A2 => n13, B1 => H(29), B2 => n14, ZN 
                           => n56);
   U65 : AOI22_X1 port map( A1 => E(29), A2 => n15, B1 => F(29), B2 => n16, ZN 
                           => n55);
   U66 : AOI22_X1 port map( A1 => C(29), A2 => n7, B1 => D(29), B2 => n5, ZN =>
                           n54);
   U67 : AOI22_X1 port map( A1 => A(29), A2 => n8, B1 => B(29), B2 => n6, ZN =>
                           n53);
   U68 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           Y(28));
   U69 : AOI22_X1 port map( A1 => G(28), A2 => n13, B1 => H(28), B2 => n14, ZN 
                           => n60);
   U70 : AOI22_X1 port map( A1 => E(28), A2 => n15, B1 => F(28), B2 => n16, ZN 
                           => n59);
   U71 : AOI22_X1 port map( A1 => C(28), A2 => n7, B1 => D(28), B2 => n5, ZN =>
                           n58);
   U72 : AOI22_X1 port map( A1 => A(28), A2 => n8, B1 => B(28), B2 => n6, ZN =>
                           n57);
   U73 : NAND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           Y(27));
   U74 : AOI22_X1 port map( A1 => G(27), A2 => n13, B1 => H(27), B2 => n14, ZN 
                           => n64);
   U75 : AOI22_X1 port map( A1 => E(27), A2 => n15, B1 => F(27), B2 => n16, ZN 
                           => n63);
   U76 : AOI22_X1 port map( A1 => C(27), A2 => n7, B1 => D(27), B2 => n5, ZN =>
                           n62);
   U77 : AOI22_X1 port map( A1 => A(27), A2 => n8, B1 => B(27), B2 => n6, ZN =>
                           n61);
   U78 : NAND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n68, ZN => 
                           Y(26));
   U79 : AOI22_X1 port map( A1 => G(26), A2 => n13, B1 => H(26), B2 => n14, ZN 
                           => n68);
   U80 : AOI22_X1 port map( A1 => E(26), A2 => n15, B1 => F(26), B2 => n16, ZN 
                           => n67);
   U81 : AOI22_X1 port map( A1 => C(26), A2 => n7, B1 => D(26), B2 => n5, ZN =>
                           n66);
   U82 : AOI22_X1 port map( A1 => A(26), A2 => n8, B1 => B(26), B2 => n6, ZN =>
                           n65);
   U83 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           Y(25));
   U84 : AOI22_X1 port map( A1 => G(25), A2 => n13, B1 => H(25), B2 => n14, ZN 
                           => n72);
   U85 : AOI22_X1 port map( A1 => E(25), A2 => n15, B1 => F(25), B2 => n16, ZN 
                           => n71);
   U86 : AOI22_X1 port map( A1 => C(25), A2 => n7, B1 => D(25), B2 => n5, ZN =>
                           n70);
   U87 : AOI22_X1 port map( A1 => A(25), A2 => n8, B1 => B(25), B2 => n6, ZN =>
                           n69);
   U88 : NAND4_X1 port map( A1 => n73, A2 => n74, A3 => n75, A4 => n76, ZN => 
                           Y(24));
   U89 : AOI22_X1 port map( A1 => G(24), A2 => n13, B1 => H(24), B2 => n14, ZN 
                           => n76);
   U90 : AOI22_X1 port map( A1 => E(24), A2 => n15, B1 => F(24), B2 => n16, ZN 
                           => n75);
   U91 : AOI22_X1 port map( A1 => C(24), A2 => n7, B1 => D(24), B2 => n5, ZN =>
                           n74);
   U92 : AOI22_X1 port map( A1 => A(24), A2 => n8, B1 => B(24), B2 => n6, ZN =>
                           n73);
   U93 : NAND4_X1 port map( A1 => n77, A2 => n78, A3 => n79, A4 => n80, ZN => 
                           Y(23));
   U94 : AOI22_X1 port map( A1 => G(23), A2 => n13, B1 => H(23), B2 => n14, ZN 
                           => n80);
   U95 : AOI22_X1 port map( A1 => E(23), A2 => n15, B1 => F(23), B2 => n16, ZN 
                           => n79);
   U96 : AOI22_X1 port map( A1 => C(23), A2 => n7, B1 => D(23), B2 => n5, ZN =>
                           n78);
   U97 : AOI22_X1 port map( A1 => A(23), A2 => n8, B1 => B(23), B2 => n6, ZN =>
                           n77);
   U98 : NAND4_X1 port map( A1 => n81, A2 => n82, A3 => n83, A4 => n84, ZN => 
                           Y(22));
   U99 : AOI22_X1 port map( A1 => G(22), A2 => n13, B1 => H(22), B2 => n14, ZN 
                           => n84);
   U100 : AOI22_X1 port map( A1 => E(22), A2 => n15, B1 => F(22), B2 => n16, ZN
                           => n83);
   U101 : AOI22_X1 port map( A1 => C(22), A2 => n7, B1 => D(22), B2 => n5, ZN 
                           => n82);
   U102 : AOI22_X1 port map( A1 => A(22), A2 => n8, B1 => B(22), B2 => n6, ZN 
                           => n81);
   U103 : NAND4_X1 port map( A1 => n85, A2 => n86, A3 => n87, A4 => n88, ZN => 
                           Y(21));
   U104 : AOI22_X1 port map( A1 => G(21), A2 => n13, B1 => H(21), B2 => n14, ZN
                           => n88);
   U105 : AOI22_X1 port map( A1 => E(21), A2 => n15, B1 => F(21), B2 => n16, ZN
                           => n87);
   U106 : AOI22_X1 port map( A1 => C(21), A2 => n7, B1 => D(21), B2 => n5, ZN 
                           => n86);
   U107 : AOI22_X1 port map( A1 => A(21), A2 => n8, B1 => B(21), B2 => n6, ZN 
                           => n85);
   U108 : NAND4_X1 port map( A1 => n89, A2 => n90, A3 => n91, A4 => n92, ZN => 
                           Y(20));
   U109 : AOI22_X1 port map( A1 => G(20), A2 => n13, B1 => H(20), B2 => n14, ZN
                           => n92);
   U110 : AOI22_X1 port map( A1 => E(20), A2 => n15, B1 => F(20), B2 => n16, ZN
                           => n91);
   U111 : AOI22_X1 port map( A1 => C(20), A2 => n7, B1 => D(20), B2 => n5, ZN 
                           => n90);
   U112 : AOI22_X1 port map( A1 => A(20), A2 => n8, B1 => B(20), B2 => n6, ZN 
                           => n89);
   U113 : NAND4_X1 port map( A1 => n93, A2 => n94, A3 => n95, A4 => n96, ZN => 
                           Y(1));
   U114 : AOI22_X1 port map( A1 => G(1), A2 => n13, B1 => H(1), B2 => n14, ZN 
                           => n96);
   U115 : AOI22_X1 port map( A1 => E(1), A2 => n15, B1 => F(1), B2 => n16, ZN 
                           => n95);
   U116 : AOI22_X1 port map( A1 => C(1), A2 => n7, B1 => D(1), B2 => n5, ZN => 
                           n94);
   U117 : AOI22_X1 port map( A1 => A(1), A2 => n8, B1 => B(1), B2 => n6, ZN => 
                           n93);
   U118 : NAND4_X1 port map( A1 => n97, A2 => n98, A3 => n99, A4 => n100, ZN =>
                           Y(19));
   U119 : AOI22_X1 port map( A1 => G(19), A2 => n13, B1 => H(19), B2 => n14, ZN
                           => n100);
   U120 : AOI22_X1 port map( A1 => E(19), A2 => n15, B1 => F(19), B2 => n16, ZN
                           => n99);
   U121 : AOI22_X1 port map( A1 => C(19), A2 => n7, B1 => D(19), B2 => n5, ZN 
                           => n98);
   U122 : AOI22_X1 port map( A1 => A(19), A2 => n8, B1 => B(19), B2 => n6, ZN 
                           => n97);
   U123 : NAND4_X1 port map( A1 => n101, A2 => n102, A3 => n103, A4 => n104, ZN
                           => Y(18));
   U124 : AOI22_X1 port map( A1 => G(18), A2 => n13, B1 => H(18), B2 => n14, ZN
                           => n104);
   U125 : AOI22_X1 port map( A1 => E(18), A2 => n15, B1 => F(18), B2 => n16, ZN
                           => n103);
   U126 : AOI22_X1 port map( A1 => C(18), A2 => n7, B1 => D(18), B2 => n5, ZN 
                           => n102);
   U127 : AOI22_X1 port map( A1 => A(18), A2 => n8, B1 => B(18), B2 => n6, ZN 
                           => n101);
   U128 : NAND4_X1 port map( A1 => n105, A2 => n106, A3 => n107, A4 => n108, ZN
                           => Y(17));
   U129 : AOI22_X1 port map( A1 => G(17), A2 => n13, B1 => H(17), B2 => n14, ZN
                           => n108);
   U130 : AOI22_X1 port map( A1 => E(17), A2 => n15, B1 => F(17), B2 => n16, ZN
                           => n107);
   U131 : AOI22_X1 port map( A1 => C(17), A2 => n7, B1 => D(17), B2 => n5, ZN 
                           => n106);
   U132 : AOI22_X1 port map( A1 => A(17), A2 => n8, B1 => B(17), B2 => n6, ZN 
                           => n105);
   U133 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n111, A4 => n112, ZN
                           => Y(16));
   U134 : AOI22_X1 port map( A1 => G(16), A2 => n13, B1 => H(16), B2 => n14, ZN
                           => n112);
   U135 : AOI22_X1 port map( A1 => E(16), A2 => n15, B1 => F(16), B2 => n16, ZN
                           => n111);
   U136 : AOI22_X1 port map( A1 => C(16), A2 => n7, B1 => D(16), B2 => n5, ZN 
                           => n110);
   U137 : AOI22_X1 port map( A1 => A(16), A2 => n8, B1 => B(16), B2 => n6, ZN 
                           => n109);
   U138 : NAND4_X1 port map( A1 => n113, A2 => n114, A3 => n115, A4 => n116, ZN
                           => Y(15));
   U139 : AOI22_X1 port map( A1 => G(15), A2 => n13, B1 => H(15), B2 => n14, ZN
                           => n116);
   U140 : AOI22_X1 port map( A1 => E(15), A2 => n15, B1 => F(15), B2 => n16, ZN
                           => n115);
   U141 : AOI22_X1 port map( A1 => C(15), A2 => n7, B1 => D(15), B2 => n5, ZN 
                           => n114);
   U142 : AOI22_X1 port map( A1 => A(15), A2 => n8, B1 => B(15), B2 => n6, ZN 
                           => n113);
   U143 : NAND4_X1 port map( A1 => n117, A2 => n118, A3 => n119, A4 => n120, ZN
                           => Y(14));
   U144 : AOI22_X1 port map( A1 => G(14), A2 => n13, B1 => H(14), B2 => n14, ZN
                           => n120);
   U145 : AOI22_X1 port map( A1 => E(14), A2 => n15, B1 => F(14), B2 => n16, ZN
                           => n119);
   U146 : AOI22_X1 port map( A1 => C(14), A2 => n7, B1 => D(14), B2 => n5, ZN 
                           => n118);
   U147 : AOI22_X1 port map( A1 => A(14), A2 => n8, B1 => B(14), B2 => n6, ZN 
                           => n117);
   U148 : NAND4_X1 port map( A1 => n121, A2 => n122, A3 => n123, A4 => n124, ZN
                           => Y(13));
   U149 : AOI22_X1 port map( A1 => G(13), A2 => n13, B1 => H(13), B2 => n14, ZN
                           => n124);
   U150 : AOI22_X1 port map( A1 => E(13), A2 => n15, B1 => F(13), B2 => n16, ZN
                           => n123);
   U151 : AOI22_X1 port map( A1 => C(13), A2 => n7, B1 => D(13), B2 => n5, ZN 
                           => n122);
   U152 : AOI22_X1 port map( A1 => A(13), A2 => n8, B1 => B(13), B2 => n6, ZN 
                           => n121);
   U153 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => Y(12));
   U154 : AOI22_X1 port map( A1 => G(12), A2 => n13, B1 => H(12), B2 => n14, ZN
                           => n128);
   U155 : AOI22_X1 port map( A1 => E(12), A2 => n15, B1 => F(12), B2 => n16, ZN
                           => n127);
   U156 : AOI22_X1 port map( A1 => C(12), A2 => n7, B1 => D(12), B2 => n5, ZN 
                           => n126);
   U157 : AOI22_X1 port map( A1 => A(12), A2 => n8, B1 => B(12), B2 => n6, ZN 
                           => n125);
   U158 : NAND4_X1 port map( A1 => n129, A2 => n130, A3 => n131, A4 => n132, ZN
                           => Y(11));
   U159 : AOI22_X1 port map( A1 => G(11), A2 => n13, B1 => H(11), B2 => n14, ZN
                           => n132);
   U160 : AOI22_X1 port map( A1 => E(11), A2 => n15, B1 => F(11), B2 => n16, ZN
                           => n131);
   U161 : AOI22_X1 port map( A1 => C(11), A2 => n7, B1 => D(11), B2 => n5, ZN 
                           => n130);
   U162 : AOI22_X1 port map( A1 => A(11), A2 => n8, B1 => B(11), B2 => n6, ZN 
                           => n129);
   U163 : NAND4_X1 port map( A1 => n133, A2 => n134, A3 => n135, A4 => n136, ZN
                           => Y(10));
   U164 : AOI22_X1 port map( A1 => G(10), A2 => n13, B1 => H(10), B2 => n14, ZN
                           => n136);
   U165 : AOI22_X1 port map( A1 => E(10), A2 => n15, B1 => F(10), B2 => n16, ZN
                           => n135);
   U166 : AOI22_X1 port map( A1 => C(10), A2 => n7, B1 => D(10), B2 => n5, ZN 
                           => n134);
   U167 : AOI22_X1 port map( A1 => A(10), A2 => n8, B1 => B(10), B2 => n6, ZN 
                           => n133);
   U168 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => Y(0));
   U169 : AOI22_X1 port map( A1 => G(0), A2 => n13, B1 => H(0), B2 => n14, ZN 
                           => n140);
   U170 : AOI22_X1 port map( A1 => E(0), A2 => n15, B1 => F(0), B2 => n16, ZN 
                           => n139);
   U171 : AOI22_X1 port map( A1 => C(0), A2 => n7, B1 => D(0), B2 => n5, ZN => 
                           n138);
   U172 : INV_X1 port map( A => S(1), ZN => n142);
   U173 : AOI22_X1 port map( A1 => A(0), A2 => n8, B1 => B(0), B2 => n6, ZN => 
                           n137);
   U174 : INV_X1 port map( A => S(0), ZN => n141);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX81_N32_1 is

   port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX81_N32_1;

architecture SYN_BEHAVIORAL of MUX81_N32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142 : std_logic;

begin
   
   U1 : AND3_X2 port map( A1 => S(2), A2 => S(1), A3 => S(0), ZN => n10);
   U2 : AND3_X2 port map( A1 => S(2), A2 => n142, A3 => S(0), ZN => n12);
   U3 : AND3_X2 port map( A1 => S(1), A2 => n141, A3 => S(2), ZN => n9);
   U4 : AND3_X2 port map( A1 => n141, A2 => n142, A3 => S(2), ZN => n11);
   U5 : OR3_X1 port map( A1 => n142, A2 => S(2), A3 => n141, ZN => n14);
   U6 : INV_X2 port map( A => n14, ZN => n1);
   U7 : OR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n141, ZN => n16);
   U8 : INV_X2 port map( A => n16, ZN => n2);
   U9 : OR3_X1 port map( A1 => S(1), A2 => S(2), A3 => S(0), ZN => n15);
   U10 : INV_X2 port map( A => n15, ZN => n3);
   U11 : OR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n142, ZN => n13);
   U12 : INV_X2 port map( A => n13, ZN => n4);
   U13 : NAND4_X1 port map( A1 => n5, A2 => n6, A3 => n7, A4 => n8, ZN => Y(9))
                           ;
   U14 : AOI22_X1 port map( A1 => G(9), A2 => n9, B1 => H(9), B2 => n10, ZN => 
                           n8);
   U15 : AOI22_X1 port map( A1 => E(9), A2 => n11, B1 => F(9), B2 => n12, ZN =>
                           n7);
   U16 : AOI22_X1 port map( A1 => C(9), A2 => n4, B1 => D(9), B2 => n1, ZN => 
                           n6);
   U17 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => B(9), B2 => n2, ZN => 
                           n5);
   U18 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           Y(8));
   U19 : AOI22_X1 port map( A1 => G(8), A2 => n9, B1 => H(8), B2 => n10, ZN => 
                           n20);
   U20 : AOI22_X1 port map( A1 => E(8), A2 => n11, B1 => F(8), B2 => n12, ZN =>
                           n19);
   U21 : AOI22_X1 port map( A1 => C(8), A2 => n4, B1 => D(8), B2 => n1, ZN => 
                           n18);
   U22 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => n2, ZN => 
                           n17);
   U23 : NAND4_X1 port map( A1 => n21, A2 => n22, A3 => n23, A4 => n24, ZN => 
                           Y(7));
   U24 : AOI22_X1 port map( A1 => G(7), A2 => n9, B1 => H(7), B2 => n10, ZN => 
                           n24);
   U25 : AOI22_X1 port map( A1 => E(7), A2 => n11, B1 => F(7), B2 => n12, ZN =>
                           n23);
   U26 : AOI22_X1 port map( A1 => C(7), A2 => n4, B1 => D(7), B2 => n1, ZN => 
                           n22);
   U27 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => n2, ZN => 
                           n21);
   U28 : NAND4_X1 port map( A1 => n25, A2 => n26, A3 => n27, A4 => n28, ZN => 
                           Y(6));
   U29 : AOI22_X1 port map( A1 => G(6), A2 => n9, B1 => H(6), B2 => n10, ZN => 
                           n28);
   U30 : AOI22_X1 port map( A1 => E(6), A2 => n11, B1 => F(6), B2 => n12, ZN =>
                           n27);
   U31 : AOI22_X1 port map( A1 => C(6), A2 => n4, B1 => D(6), B2 => n1, ZN => 
                           n26);
   U32 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => n2, ZN => 
                           n25);
   U33 : NAND4_X1 port map( A1 => n29, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           Y(5));
   U34 : AOI22_X1 port map( A1 => G(5), A2 => n9, B1 => H(5), B2 => n10, ZN => 
                           n32);
   U35 : AOI22_X1 port map( A1 => E(5), A2 => n11, B1 => F(5), B2 => n12, ZN =>
                           n31);
   U36 : AOI22_X1 port map( A1 => C(5), A2 => n4, B1 => D(5), B2 => n1, ZN => 
                           n30);
   U37 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => n2, ZN => 
                           n29);
   U38 : NAND4_X1 port map( A1 => n33, A2 => n34, A3 => n35, A4 => n36, ZN => 
                           Y(4));
   U39 : AOI22_X1 port map( A1 => G(4), A2 => n9, B1 => H(4), B2 => n10, ZN => 
                           n36);
   U40 : AOI22_X1 port map( A1 => E(4), A2 => n11, B1 => F(4), B2 => n12, ZN =>
                           n35);
   U41 : AOI22_X1 port map( A1 => C(4), A2 => n4, B1 => D(4), B2 => n1, ZN => 
                           n34);
   U42 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => n2, ZN => 
                           n33);
   U43 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           Y(3));
   U44 : AOI22_X1 port map( A1 => G(3), A2 => n9, B1 => H(3), B2 => n10, ZN => 
                           n40);
   U45 : AOI22_X1 port map( A1 => E(3), A2 => n11, B1 => F(3), B2 => n12, ZN =>
                           n39);
   U46 : AOI22_X1 port map( A1 => C(3), A2 => n4, B1 => D(3), B2 => n1, ZN => 
                           n38);
   U47 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => n2, ZN => 
                           n37);
   U48 : NAND4_X1 port map( A1 => n41, A2 => n42, A3 => n43, A4 => n44, ZN => 
                           Y(31));
   U49 : AOI22_X1 port map( A1 => G(31), A2 => n9, B1 => H(31), B2 => n10, ZN 
                           => n44);
   U50 : AOI22_X1 port map( A1 => E(31), A2 => n11, B1 => F(31), B2 => n12, ZN 
                           => n43);
   U51 : AOI22_X1 port map( A1 => C(31), A2 => n4, B1 => D(31), B2 => n1, ZN =>
                           n42);
   U52 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => n2, ZN =>
                           n41);
   U53 : NAND4_X1 port map( A1 => n45, A2 => n46, A3 => n47, A4 => n48, ZN => 
                           Y(30));
   U54 : AOI22_X1 port map( A1 => G(30), A2 => n9, B1 => H(30), B2 => n10, ZN 
                           => n48);
   U55 : AOI22_X1 port map( A1 => E(30), A2 => n11, B1 => F(30), B2 => n12, ZN 
                           => n47);
   U56 : AOI22_X1 port map( A1 => C(30), A2 => n4, B1 => D(30), B2 => n1, ZN =>
                           n46);
   U57 : AOI22_X1 port map( A1 => A(30), A2 => n3, B1 => B(30), B2 => n2, ZN =>
                           n45);
   U58 : NAND4_X1 port map( A1 => n49, A2 => n50, A3 => n51, A4 => n52, ZN => 
                           Y(2));
   U59 : AOI22_X1 port map( A1 => G(2), A2 => n9, B1 => H(2), B2 => n10, ZN => 
                           n52);
   U60 : AOI22_X1 port map( A1 => E(2), A2 => n11, B1 => F(2), B2 => n12, ZN =>
                           n51);
   U61 : AOI22_X1 port map( A1 => C(2), A2 => n4, B1 => D(2), B2 => n1, ZN => 
                           n50);
   U62 : AOI22_X1 port map( A1 => A(2), A2 => n3, B1 => B(2), B2 => n2, ZN => 
                           n49);
   U63 : NAND4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           Y(29));
   U64 : AOI22_X1 port map( A1 => G(29), A2 => n9, B1 => H(29), B2 => n10, ZN 
                           => n56);
   U65 : AOI22_X1 port map( A1 => E(29), A2 => n11, B1 => F(29), B2 => n12, ZN 
                           => n55);
   U66 : AOI22_X1 port map( A1 => C(29), A2 => n4, B1 => D(29), B2 => n1, ZN =>
                           n54);
   U67 : AOI22_X1 port map( A1 => A(29), A2 => n3, B1 => B(29), B2 => n2, ZN =>
                           n53);
   U68 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           Y(28));
   U69 : AOI22_X1 port map( A1 => G(28), A2 => n9, B1 => H(28), B2 => n10, ZN 
                           => n60);
   U70 : AOI22_X1 port map( A1 => E(28), A2 => n11, B1 => F(28), B2 => n12, ZN 
                           => n59);
   U71 : AOI22_X1 port map( A1 => C(28), A2 => n4, B1 => D(28), B2 => n1, ZN =>
                           n58);
   U72 : AOI22_X1 port map( A1 => A(28), A2 => n3, B1 => B(28), B2 => n2, ZN =>
                           n57);
   U73 : NAND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           Y(27));
   U74 : AOI22_X1 port map( A1 => G(27), A2 => n9, B1 => H(27), B2 => n10, ZN 
                           => n64);
   U75 : AOI22_X1 port map( A1 => E(27), A2 => n11, B1 => F(27), B2 => n12, ZN 
                           => n63);
   U76 : AOI22_X1 port map( A1 => C(27), A2 => n4, B1 => D(27), B2 => n1, ZN =>
                           n62);
   U77 : AOI22_X1 port map( A1 => A(27), A2 => n3, B1 => B(27), B2 => n2, ZN =>
                           n61);
   U78 : NAND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n68, ZN => 
                           Y(26));
   U79 : AOI22_X1 port map( A1 => G(26), A2 => n9, B1 => H(26), B2 => n10, ZN 
                           => n68);
   U80 : AOI22_X1 port map( A1 => E(26), A2 => n11, B1 => F(26), B2 => n12, ZN 
                           => n67);
   U81 : AOI22_X1 port map( A1 => C(26), A2 => n4, B1 => D(26), B2 => n1, ZN =>
                           n66);
   U82 : AOI22_X1 port map( A1 => A(26), A2 => n3, B1 => B(26), B2 => n2, ZN =>
                           n65);
   U83 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           Y(25));
   U84 : AOI22_X1 port map( A1 => G(25), A2 => n9, B1 => H(25), B2 => n10, ZN 
                           => n72);
   U85 : AOI22_X1 port map( A1 => E(25), A2 => n11, B1 => F(25), B2 => n12, ZN 
                           => n71);
   U86 : AOI22_X1 port map( A1 => C(25), A2 => n4, B1 => D(25), B2 => n1, ZN =>
                           n70);
   U87 : AOI22_X1 port map( A1 => A(25), A2 => n3, B1 => B(25), B2 => n2, ZN =>
                           n69);
   U88 : NAND4_X1 port map( A1 => n73, A2 => n74, A3 => n75, A4 => n76, ZN => 
                           Y(24));
   U89 : AOI22_X1 port map( A1 => G(24), A2 => n9, B1 => H(24), B2 => n10, ZN 
                           => n76);
   U90 : AOI22_X1 port map( A1 => E(24), A2 => n11, B1 => F(24), B2 => n12, ZN 
                           => n75);
   U91 : AOI22_X1 port map( A1 => C(24), A2 => n4, B1 => D(24), B2 => n1, ZN =>
                           n74);
   U92 : AOI22_X1 port map( A1 => A(24), A2 => n3, B1 => B(24), B2 => n2, ZN =>
                           n73);
   U93 : NAND4_X1 port map( A1 => n77, A2 => n78, A3 => n79, A4 => n80, ZN => 
                           Y(23));
   U94 : AOI22_X1 port map( A1 => G(23), A2 => n9, B1 => H(23), B2 => n10, ZN 
                           => n80);
   U95 : AOI22_X1 port map( A1 => E(23), A2 => n11, B1 => F(23), B2 => n12, ZN 
                           => n79);
   U96 : AOI22_X1 port map( A1 => C(23), A2 => n4, B1 => D(23), B2 => n1, ZN =>
                           n78);
   U97 : AOI22_X1 port map( A1 => A(23), A2 => n3, B1 => B(23), B2 => n2, ZN =>
                           n77);
   U98 : NAND4_X1 port map( A1 => n81, A2 => n82, A3 => n83, A4 => n84, ZN => 
                           Y(22));
   U99 : AOI22_X1 port map( A1 => G(22), A2 => n9, B1 => H(22), B2 => n10, ZN 
                           => n84);
   U100 : AOI22_X1 port map( A1 => E(22), A2 => n11, B1 => F(22), B2 => n12, ZN
                           => n83);
   U101 : AOI22_X1 port map( A1 => C(22), A2 => n4, B1 => D(22), B2 => n1, ZN 
                           => n82);
   U102 : AOI22_X1 port map( A1 => A(22), A2 => n3, B1 => B(22), B2 => n2, ZN 
                           => n81);
   U103 : NAND4_X1 port map( A1 => n85, A2 => n86, A3 => n87, A4 => n88, ZN => 
                           Y(21));
   U104 : AOI22_X1 port map( A1 => G(21), A2 => n9, B1 => H(21), B2 => n10, ZN 
                           => n88);
   U105 : AOI22_X1 port map( A1 => E(21), A2 => n11, B1 => F(21), B2 => n12, ZN
                           => n87);
   U106 : AOI22_X1 port map( A1 => C(21), A2 => n4, B1 => D(21), B2 => n1, ZN 
                           => n86);
   U107 : AOI22_X1 port map( A1 => A(21), A2 => n3, B1 => B(21), B2 => n2, ZN 
                           => n85);
   U108 : NAND4_X1 port map( A1 => n89, A2 => n90, A3 => n91, A4 => n92, ZN => 
                           Y(20));
   U109 : AOI22_X1 port map( A1 => G(20), A2 => n9, B1 => H(20), B2 => n10, ZN 
                           => n92);
   U110 : AOI22_X1 port map( A1 => E(20), A2 => n11, B1 => F(20), B2 => n12, ZN
                           => n91);
   U111 : AOI22_X1 port map( A1 => C(20), A2 => n4, B1 => D(20), B2 => n1, ZN 
                           => n90);
   U112 : AOI22_X1 port map( A1 => A(20), A2 => n3, B1 => B(20), B2 => n2, ZN 
                           => n89);
   U113 : NAND4_X1 port map( A1 => n93, A2 => n94, A3 => n95, A4 => n96, ZN => 
                           Y(1));
   U114 : AOI22_X1 port map( A1 => G(1), A2 => n9, B1 => H(1), B2 => n10, ZN =>
                           n96);
   U115 : AOI22_X1 port map( A1 => E(1), A2 => n11, B1 => F(1), B2 => n12, ZN 
                           => n95);
   U116 : AOI22_X1 port map( A1 => C(1), A2 => n4, B1 => D(1), B2 => n1, ZN => 
                           n94);
   U117 : AOI22_X1 port map( A1 => A(1), A2 => n3, B1 => B(1), B2 => n2, ZN => 
                           n93);
   U118 : NAND4_X1 port map( A1 => n97, A2 => n98, A3 => n99, A4 => n100, ZN =>
                           Y(19));
   U119 : AOI22_X1 port map( A1 => G(19), A2 => n9, B1 => H(19), B2 => n10, ZN 
                           => n100);
   U120 : AOI22_X1 port map( A1 => E(19), A2 => n11, B1 => F(19), B2 => n12, ZN
                           => n99);
   U121 : AOI22_X1 port map( A1 => C(19), A2 => n4, B1 => D(19), B2 => n1, ZN 
                           => n98);
   U122 : AOI22_X1 port map( A1 => A(19), A2 => n3, B1 => B(19), B2 => n2, ZN 
                           => n97);
   U123 : NAND4_X1 port map( A1 => n101, A2 => n102, A3 => n103, A4 => n104, ZN
                           => Y(18));
   U124 : AOI22_X1 port map( A1 => G(18), A2 => n9, B1 => H(18), B2 => n10, ZN 
                           => n104);
   U125 : AOI22_X1 port map( A1 => E(18), A2 => n11, B1 => F(18), B2 => n12, ZN
                           => n103);
   U126 : AOI22_X1 port map( A1 => C(18), A2 => n4, B1 => D(18), B2 => n1, ZN 
                           => n102);
   U127 : AOI22_X1 port map( A1 => A(18), A2 => n3, B1 => B(18), B2 => n2, ZN 
                           => n101);
   U128 : NAND4_X1 port map( A1 => n105, A2 => n106, A3 => n107, A4 => n108, ZN
                           => Y(17));
   U129 : AOI22_X1 port map( A1 => G(17), A2 => n9, B1 => H(17), B2 => n10, ZN 
                           => n108);
   U130 : AOI22_X1 port map( A1 => E(17), A2 => n11, B1 => F(17), B2 => n12, ZN
                           => n107);
   U131 : AOI22_X1 port map( A1 => C(17), A2 => n4, B1 => D(17), B2 => n1, ZN 
                           => n106);
   U132 : AOI22_X1 port map( A1 => A(17), A2 => n3, B1 => B(17), B2 => n2, ZN 
                           => n105);
   U133 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n111, A4 => n112, ZN
                           => Y(16));
   U134 : AOI22_X1 port map( A1 => G(16), A2 => n9, B1 => H(16), B2 => n10, ZN 
                           => n112);
   U135 : AOI22_X1 port map( A1 => E(16), A2 => n11, B1 => F(16), B2 => n12, ZN
                           => n111);
   U136 : AOI22_X1 port map( A1 => C(16), A2 => n4, B1 => D(16), B2 => n1, ZN 
                           => n110);
   U137 : AOI22_X1 port map( A1 => A(16), A2 => n3, B1 => B(16), B2 => n2, ZN 
                           => n109);
   U138 : NAND4_X1 port map( A1 => n113, A2 => n114, A3 => n115, A4 => n116, ZN
                           => Y(15));
   U139 : AOI22_X1 port map( A1 => G(15), A2 => n9, B1 => H(15), B2 => n10, ZN 
                           => n116);
   U140 : AOI22_X1 port map( A1 => E(15), A2 => n11, B1 => F(15), B2 => n12, ZN
                           => n115);
   U141 : AOI22_X1 port map( A1 => C(15), A2 => n4, B1 => D(15), B2 => n1, ZN 
                           => n114);
   U142 : AOI22_X1 port map( A1 => A(15), A2 => n3, B1 => B(15), B2 => n2, ZN 
                           => n113);
   U143 : NAND4_X1 port map( A1 => n117, A2 => n118, A3 => n119, A4 => n120, ZN
                           => Y(14));
   U144 : AOI22_X1 port map( A1 => G(14), A2 => n9, B1 => H(14), B2 => n10, ZN 
                           => n120);
   U145 : AOI22_X1 port map( A1 => E(14), A2 => n11, B1 => F(14), B2 => n12, ZN
                           => n119);
   U146 : AOI22_X1 port map( A1 => C(14), A2 => n4, B1 => D(14), B2 => n1, ZN 
                           => n118);
   U147 : AOI22_X1 port map( A1 => A(14), A2 => n3, B1 => B(14), B2 => n2, ZN 
                           => n117);
   U148 : NAND4_X1 port map( A1 => n121, A2 => n122, A3 => n123, A4 => n124, ZN
                           => Y(13));
   U149 : AOI22_X1 port map( A1 => G(13), A2 => n9, B1 => H(13), B2 => n10, ZN 
                           => n124);
   U150 : AOI22_X1 port map( A1 => E(13), A2 => n11, B1 => F(13), B2 => n12, ZN
                           => n123);
   U151 : AOI22_X1 port map( A1 => C(13), A2 => n4, B1 => D(13), B2 => n1, ZN 
                           => n122);
   U152 : AOI22_X1 port map( A1 => A(13), A2 => n3, B1 => B(13), B2 => n2, ZN 
                           => n121);
   U153 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => Y(12));
   U154 : AOI22_X1 port map( A1 => G(12), A2 => n9, B1 => H(12), B2 => n10, ZN 
                           => n128);
   U155 : AOI22_X1 port map( A1 => E(12), A2 => n11, B1 => F(12), B2 => n12, ZN
                           => n127);
   U156 : AOI22_X1 port map( A1 => C(12), A2 => n4, B1 => D(12), B2 => n1, ZN 
                           => n126);
   U157 : AOI22_X1 port map( A1 => A(12), A2 => n3, B1 => B(12), B2 => n2, ZN 
                           => n125);
   U158 : NAND4_X1 port map( A1 => n129, A2 => n130, A3 => n131, A4 => n132, ZN
                           => Y(11));
   U159 : AOI22_X1 port map( A1 => G(11), A2 => n9, B1 => H(11), B2 => n10, ZN 
                           => n132);
   U160 : AOI22_X1 port map( A1 => E(11), A2 => n11, B1 => F(11), B2 => n12, ZN
                           => n131);
   U161 : AOI22_X1 port map( A1 => C(11), A2 => n4, B1 => D(11), B2 => n1, ZN 
                           => n130);
   U162 : AOI22_X1 port map( A1 => A(11), A2 => n3, B1 => B(11), B2 => n2, ZN 
                           => n129);
   U163 : NAND4_X1 port map( A1 => n133, A2 => n134, A3 => n135, A4 => n136, ZN
                           => Y(10));
   U164 : AOI22_X1 port map( A1 => G(10), A2 => n9, B1 => H(10), B2 => n10, ZN 
                           => n136);
   U165 : AOI22_X1 port map( A1 => E(10), A2 => n11, B1 => F(10), B2 => n12, ZN
                           => n135);
   U166 : AOI22_X1 port map( A1 => C(10), A2 => n4, B1 => D(10), B2 => n1, ZN 
                           => n134);
   U167 : AOI22_X1 port map( A1 => A(10), A2 => n3, B1 => B(10), B2 => n2, ZN 
                           => n133);
   U168 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => Y(0));
   U169 : AOI22_X1 port map( A1 => G(0), A2 => n9, B1 => H(0), B2 => n10, ZN =>
                           n140);
   U170 : AOI22_X1 port map( A1 => E(0), A2 => n11, B1 => F(0), B2 => n12, ZN 
                           => n139);
   U171 : AOI22_X1 port map( A1 => C(0), A2 => n4, B1 => D(0), B2 => n1, ZN => 
                           n138);
   U172 : INV_X1 port map( A => S(1), ZN => n142);
   U173 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => n2, ZN => 
                           n137);
   U174 : INV_X1 port map( A => S(0), ZN => n141);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX81_N32_0 is

   port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX81_N32_0;

architecture SYN_BEHAVIORAL of MUX81_N32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142 : std_logic;

begin
   
   U1 : AND3_X2 port map( A1 => S(2), A2 => S(1), A3 => S(0), ZN => n10);
   U2 : AND3_X2 port map( A1 => S(2), A2 => n142, A3 => S(0), ZN => n12);
   U3 : AND3_X2 port map( A1 => S(1), A2 => n141, A3 => S(2), ZN => n9);
   U4 : AND3_X2 port map( A1 => n141, A2 => n142, A3 => S(2), ZN => n11);
   U5 : OR3_X1 port map( A1 => n142, A2 => S(2), A3 => n141, ZN => n14);
   U6 : INV_X2 port map( A => n14, ZN => n1);
   U7 : OR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n141, ZN => n16);
   U8 : INV_X2 port map( A => n16, ZN => n2);
   U9 : OR3_X1 port map( A1 => S(1), A2 => S(2), A3 => S(0), ZN => n15);
   U10 : INV_X2 port map( A => n15, ZN => n3);
   U11 : OR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n142, ZN => n13);
   U12 : INV_X2 port map( A => n13, ZN => n4);
   U13 : NAND4_X1 port map( A1 => n5, A2 => n6, A3 => n7, A4 => n8, ZN => Y(9))
                           ;
   U14 : AOI22_X1 port map( A1 => G(9), A2 => n9, B1 => H(9), B2 => n10, ZN => 
                           n8);
   U15 : AOI22_X1 port map( A1 => E(9), A2 => n11, B1 => F(9), B2 => n12, ZN =>
                           n7);
   U16 : AOI22_X1 port map( A1 => C(9), A2 => n4, B1 => D(9), B2 => n1, ZN => 
                           n6);
   U17 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => B(9), B2 => n2, ZN => 
                           n5);
   U18 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           Y(8));
   U19 : AOI22_X1 port map( A1 => G(8), A2 => n9, B1 => H(8), B2 => n10, ZN => 
                           n20);
   U20 : AOI22_X1 port map( A1 => E(8), A2 => n11, B1 => F(8), B2 => n12, ZN =>
                           n19);
   U21 : AOI22_X1 port map( A1 => C(8), A2 => n4, B1 => D(8), B2 => n1, ZN => 
                           n18);
   U22 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => n2, ZN => 
                           n17);
   U23 : NAND4_X1 port map( A1 => n21, A2 => n22, A3 => n23, A4 => n24, ZN => 
                           Y(7));
   U24 : AOI22_X1 port map( A1 => G(7), A2 => n9, B1 => H(7), B2 => n10, ZN => 
                           n24);
   U25 : AOI22_X1 port map( A1 => E(7), A2 => n11, B1 => F(7), B2 => n12, ZN =>
                           n23);
   U26 : AOI22_X1 port map( A1 => C(7), A2 => n4, B1 => D(7), B2 => n1, ZN => 
                           n22);
   U27 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => n2, ZN => 
                           n21);
   U28 : NAND4_X1 port map( A1 => n25, A2 => n26, A3 => n27, A4 => n28, ZN => 
                           Y(6));
   U29 : AOI22_X1 port map( A1 => G(6), A2 => n9, B1 => H(6), B2 => n10, ZN => 
                           n28);
   U30 : AOI22_X1 port map( A1 => E(6), A2 => n11, B1 => F(6), B2 => n12, ZN =>
                           n27);
   U31 : AOI22_X1 port map( A1 => C(6), A2 => n4, B1 => D(6), B2 => n1, ZN => 
                           n26);
   U32 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => n2, ZN => 
                           n25);
   U33 : NAND4_X1 port map( A1 => n29, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           Y(5));
   U34 : AOI22_X1 port map( A1 => G(5), A2 => n9, B1 => H(5), B2 => n10, ZN => 
                           n32);
   U35 : AOI22_X1 port map( A1 => E(5), A2 => n11, B1 => F(5), B2 => n12, ZN =>
                           n31);
   U36 : AOI22_X1 port map( A1 => C(5), A2 => n4, B1 => D(5), B2 => n1, ZN => 
                           n30);
   U37 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => n2, ZN => 
                           n29);
   U38 : NAND4_X1 port map( A1 => n33, A2 => n34, A3 => n35, A4 => n36, ZN => 
                           Y(4));
   U39 : AOI22_X1 port map( A1 => G(4), A2 => n9, B1 => H(4), B2 => n10, ZN => 
                           n36);
   U40 : AOI22_X1 port map( A1 => E(4), A2 => n11, B1 => F(4), B2 => n12, ZN =>
                           n35);
   U41 : AOI22_X1 port map( A1 => C(4), A2 => n4, B1 => D(4), B2 => n1, ZN => 
                           n34);
   U42 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => n2, ZN => 
                           n33);
   U43 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           Y(3));
   U44 : AOI22_X1 port map( A1 => G(3), A2 => n9, B1 => H(3), B2 => n10, ZN => 
                           n40);
   U45 : AOI22_X1 port map( A1 => E(3), A2 => n11, B1 => F(3), B2 => n12, ZN =>
                           n39);
   U46 : AOI22_X1 port map( A1 => C(3), A2 => n4, B1 => D(3), B2 => n1, ZN => 
                           n38);
   U47 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => n2, ZN => 
                           n37);
   U48 : NAND4_X1 port map( A1 => n41, A2 => n42, A3 => n43, A4 => n44, ZN => 
                           Y(31));
   U49 : AOI22_X1 port map( A1 => G(31), A2 => n9, B1 => H(31), B2 => n10, ZN 
                           => n44);
   U50 : AOI22_X1 port map( A1 => E(31), A2 => n11, B1 => F(31), B2 => n12, ZN 
                           => n43);
   U51 : AOI22_X1 port map( A1 => C(31), A2 => n4, B1 => D(31), B2 => n1, ZN =>
                           n42);
   U52 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => n2, ZN =>
                           n41);
   U53 : NAND4_X1 port map( A1 => n45, A2 => n46, A3 => n47, A4 => n48, ZN => 
                           Y(30));
   U54 : AOI22_X1 port map( A1 => G(30), A2 => n9, B1 => H(30), B2 => n10, ZN 
                           => n48);
   U55 : AOI22_X1 port map( A1 => E(30), A2 => n11, B1 => F(30), B2 => n12, ZN 
                           => n47);
   U56 : AOI22_X1 port map( A1 => C(30), A2 => n4, B1 => D(30), B2 => n1, ZN =>
                           n46);
   U57 : AOI22_X1 port map( A1 => A(30), A2 => n3, B1 => B(30), B2 => n2, ZN =>
                           n45);
   U58 : NAND4_X1 port map( A1 => n49, A2 => n50, A3 => n51, A4 => n52, ZN => 
                           Y(2));
   U59 : AOI22_X1 port map( A1 => G(2), A2 => n9, B1 => H(2), B2 => n10, ZN => 
                           n52);
   U60 : AOI22_X1 port map( A1 => E(2), A2 => n11, B1 => F(2), B2 => n12, ZN =>
                           n51);
   U61 : AOI22_X1 port map( A1 => C(2), A2 => n4, B1 => D(2), B2 => n1, ZN => 
                           n50);
   U62 : AOI22_X1 port map( A1 => A(2), A2 => n3, B1 => B(2), B2 => n2, ZN => 
                           n49);
   U63 : NAND4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           Y(29));
   U64 : AOI22_X1 port map( A1 => G(29), A2 => n9, B1 => H(29), B2 => n10, ZN 
                           => n56);
   U65 : AOI22_X1 port map( A1 => E(29), A2 => n11, B1 => F(29), B2 => n12, ZN 
                           => n55);
   U66 : AOI22_X1 port map( A1 => C(29), A2 => n4, B1 => D(29), B2 => n1, ZN =>
                           n54);
   U67 : AOI22_X1 port map( A1 => A(29), A2 => n3, B1 => B(29), B2 => n2, ZN =>
                           n53);
   U68 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           Y(28));
   U69 : AOI22_X1 port map( A1 => G(28), A2 => n9, B1 => H(28), B2 => n10, ZN 
                           => n60);
   U70 : AOI22_X1 port map( A1 => E(28), A2 => n11, B1 => F(28), B2 => n12, ZN 
                           => n59);
   U71 : AOI22_X1 port map( A1 => C(28), A2 => n4, B1 => D(28), B2 => n1, ZN =>
                           n58);
   U72 : AOI22_X1 port map( A1 => A(28), A2 => n3, B1 => B(28), B2 => n2, ZN =>
                           n57);
   U73 : NAND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           Y(27));
   U74 : AOI22_X1 port map( A1 => G(27), A2 => n9, B1 => H(27), B2 => n10, ZN 
                           => n64);
   U75 : AOI22_X1 port map( A1 => E(27), A2 => n11, B1 => F(27), B2 => n12, ZN 
                           => n63);
   U76 : AOI22_X1 port map( A1 => C(27), A2 => n4, B1 => D(27), B2 => n1, ZN =>
                           n62);
   U77 : AOI22_X1 port map( A1 => A(27), A2 => n3, B1 => B(27), B2 => n2, ZN =>
                           n61);
   U78 : NAND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n68, ZN => 
                           Y(26));
   U79 : AOI22_X1 port map( A1 => G(26), A2 => n9, B1 => H(26), B2 => n10, ZN 
                           => n68);
   U80 : AOI22_X1 port map( A1 => E(26), A2 => n11, B1 => F(26), B2 => n12, ZN 
                           => n67);
   U81 : AOI22_X1 port map( A1 => C(26), A2 => n4, B1 => D(26), B2 => n1, ZN =>
                           n66);
   U82 : AOI22_X1 port map( A1 => A(26), A2 => n3, B1 => B(26), B2 => n2, ZN =>
                           n65);
   U83 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           Y(25));
   U84 : AOI22_X1 port map( A1 => G(25), A2 => n9, B1 => H(25), B2 => n10, ZN 
                           => n72);
   U85 : AOI22_X1 port map( A1 => E(25), A2 => n11, B1 => F(25), B2 => n12, ZN 
                           => n71);
   U86 : AOI22_X1 port map( A1 => C(25), A2 => n4, B1 => D(25), B2 => n1, ZN =>
                           n70);
   U87 : AOI22_X1 port map( A1 => A(25), A2 => n3, B1 => B(25), B2 => n2, ZN =>
                           n69);
   U88 : NAND4_X1 port map( A1 => n73, A2 => n74, A3 => n75, A4 => n76, ZN => 
                           Y(24));
   U89 : AOI22_X1 port map( A1 => G(24), A2 => n9, B1 => H(24), B2 => n10, ZN 
                           => n76);
   U90 : AOI22_X1 port map( A1 => E(24), A2 => n11, B1 => F(24), B2 => n12, ZN 
                           => n75);
   U91 : AOI22_X1 port map( A1 => C(24), A2 => n4, B1 => D(24), B2 => n1, ZN =>
                           n74);
   U92 : AOI22_X1 port map( A1 => A(24), A2 => n3, B1 => B(24), B2 => n2, ZN =>
                           n73);
   U93 : NAND4_X1 port map( A1 => n77, A2 => n78, A3 => n79, A4 => n80, ZN => 
                           Y(23));
   U94 : AOI22_X1 port map( A1 => G(23), A2 => n9, B1 => H(23), B2 => n10, ZN 
                           => n80);
   U95 : AOI22_X1 port map( A1 => E(23), A2 => n11, B1 => F(23), B2 => n12, ZN 
                           => n79);
   U96 : AOI22_X1 port map( A1 => C(23), A2 => n4, B1 => D(23), B2 => n1, ZN =>
                           n78);
   U97 : AOI22_X1 port map( A1 => A(23), A2 => n3, B1 => B(23), B2 => n2, ZN =>
                           n77);
   U98 : NAND4_X1 port map( A1 => n81, A2 => n82, A3 => n83, A4 => n84, ZN => 
                           Y(22));
   U99 : AOI22_X1 port map( A1 => G(22), A2 => n9, B1 => H(22), B2 => n10, ZN 
                           => n84);
   U100 : AOI22_X1 port map( A1 => E(22), A2 => n11, B1 => F(22), B2 => n12, ZN
                           => n83);
   U101 : AOI22_X1 port map( A1 => C(22), A2 => n4, B1 => D(22), B2 => n1, ZN 
                           => n82);
   U102 : AOI22_X1 port map( A1 => A(22), A2 => n3, B1 => B(22), B2 => n2, ZN 
                           => n81);
   U103 : NAND4_X1 port map( A1 => n85, A2 => n86, A3 => n87, A4 => n88, ZN => 
                           Y(21));
   U104 : AOI22_X1 port map( A1 => G(21), A2 => n9, B1 => H(21), B2 => n10, ZN 
                           => n88);
   U105 : AOI22_X1 port map( A1 => E(21), A2 => n11, B1 => F(21), B2 => n12, ZN
                           => n87);
   U106 : AOI22_X1 port map( A1 => C(21), A2 => n4, B1 => D(21), B2 => n1, ZN 
                           => n86);
   U107 : AOI22_X1 port map( A1 => A(21), A2 => n3, B1 => B(21), B2 => n2, ZN 
                           => n85);
   U108 : NAND4_X1 port map( A1 => n89, A2 => n90, A3 => n91, A4 => n92, ZN => 
                           Y(20));
   U109 : AOI22_X1 port map( A1 => G(20), A2 => n9, B1 => H(20), B2 => n10, ZN 
                           => n92);
   U110 : AOI22_X1 port map( A1 => E(20), A2 => n11, B1 => F(20), B2 => n12, ZN
                           => n91);
   U111 : AOI22_X1 port map( A1 => C(20), A2 => n4, B1 => D(20), B2 => n1, ZN 
                           => n90);
   U112 : AOI22_X1 port map( A1 => A(20), A2 => n3, B1 => B(20), B2 => n2, ZN 
                           => n89);
   U113 : NAND4_X1 port map( A1 => n93, A2 => n94, A3 => n95, A4 => n96, ZN => 
                           Y(1));
   U114 : AOI22_X1 port map( A1 => G(1), A2 => n9, B1 => H(1), B2 => n10, ZN =>
                           n96);
   U115 : AOI22_X1 port map( A1 => E(1), A2 => n11, B1 => F(1), B2 => n12, ZN 
                           => n95);
   U116 : AOI22_X1 port map( A1 => C(1), A2 => n4, B1 => D(1), B2 => n1, ZN => 
                           n94);
   U117 : AOI22_X1 port map( A1 => A(1), A2 => n3, B1 => B(1), B2 => n2, ZN => 
                           n93);
   U118 : NAND4_X1 port map( A1 => n97, A2 => n98, A3 => n99, A4 => n100, ZN =>
                           Y(19));
   U119 : AOI22_X1 port map( A1 => G(19), A2 => n9, B1 => H(19), B2 => n10, ZN 
                           => n100);
   U120 : AOI22_X1 port map( A1 => E(19), A2 => n11, B1 => F(19), B2 => n12, ZN
                           => n99);
   U121 : AOI22_X1 port map( A1 => C(19), A2 => n4, B1 => D(19), B2 => n1, ZN 
                           => n98);
   U122 : AOI22_X1 port map( A1 => A(19), A2 => n3, B1 => B(19), B2 => n2, ZN 
                           => n97);
   U123 : NAND4_X1 port map( A1 => n101, A2 => n102, A3 => n103, A4 => n104, ZN
                           => Y(18));
   U124 : AOI22_X1 port map( A1 => G(18), A2 => n9, B1 => H(18), B2 => n10, ZN 
                           => n104);
   U125 : AOI22_X1 port map( A1 => E(18), A2 => n11, B1 => F(18), B2 => n12, ZN
                           => n103);
   U126 : AOI22_X1 port map( A1 => C(18), A2 => n4, B1 => D(18), B2 => n1, ZN 
                           => n102);
   U127 : AOI22_X1 port map( A1 => A(18), A2 => n3, B1 => B(18), B2 => n2, ZN 
                           => n101);
   U128 : NAND4_X1 port map( A1 => n105, A2 => n106, A3 => n107, A4 => n108, ZN
                           => Y(17));
   U129 : AOI22_X1 port map( A1 => G(17), A2 => n9, B1 => H(17), B2 => n10, ZN 
                           => n108);
   U130 : AOI22_X1 port map( A1 => E(17), A2 => n11, B1 => F(17), B2 => n12, ZN
                           => n107);
   U131 : AOI22_X1 port map( A1 => C(17), A2 => n4, B1 => D(17), B2 => n1, ZN 
                           => n106);
   U132 : AOI22_X1 port map( A1 => A(17), A2 => n3, B1 => B(17), B2 => n2, ZN 
                           => n105);
   U133 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n111, A4 => n112, ZN
                           => Y(16));
   U134 : AOI22_X1 port map( A1 => G(16), A2 => n9, B1 => H(16), B2 => n10, ZN 
                           => n112);
   U135 : AOI22_X1 port map( A1 => E(16), A2 => n11, B1 => F(16), B2 => n12, ZN
                           => n111);
   U136 : AOI22_X1 port map( A1 => C(16), A2 => n4, B1 => D(16), B2 => n1, ZN 
                           => n110);
   U137 : AOI22_X1 port map( A1 => A(16), A2 => n3, B1 => B(16), B2 => n2, ZN 
                           => n109);
   U138 : NAND4_X1 port map( A1 => n113, A2 => n114, A3 => n115, A4 => n116, ZN
                           => Y(15));
   U139 : AOI22_X1 port map( A1 => G(15), A2 => n9, B1 => H(15), B2 => n10, ZN 
                           => n116);
   U140 : AOI22_X1 port map( A1 => E(15), A2 => n11, B1 => F(15), B2 => n12, ZN
                           => n115);
   U141 : AOI22_X1 port map( A1 => C(15), A2 => n4, B1 => D(15), B2 => n1, ZN 
                           => n114);
   U142 : AOI22_X1 port map( A1 => A(15), A2 => n3, B1 => B(15), B2 => n2, ZN 
                           => n113);
   U143 : NAND4_X1 port map( A1 => n117, A2 => n118, A3 => n119, A4 => n120, ZN
                           => Y(14));
   U144 : AOI22_X1 port map( A1 => G(14), A2 => n9, B1 => H(14), B2 => n10, ZN 
                           => n120);
   U145 : AOI22_X1 port map( A1 => E(14), A2 => n11, B1 => F(14), B2 => n12, ZN
                           => n119);
   U146 : AOI22_X1 port map( A1 => C(14), A2 => n4, B1 => D(14), B2 => n1, ZN 
                           => n118);
   U147 : AOI22_X1 port map( A1 => A(14), A2 => n3, B1 => B(14), B2 => n2, ZN 
                           => n117);
   U148 : NAND4_X1 port map( A1 => n121, A2 => n122, A3 => n123, A4 => n124, ZN
                           => Y(13));
   U149 : AOI22_X1 port map( A1 => G(13), A2 => n9, B1 => H(13), B2 => n10, ZN 
                           => n124);
   U150 : AOI22_X1 port map( A1 => E(13), A2 => n11, B1 => F(13), B2 => n12, ZN
                           => n123);
   U151 : AOI22_X1 port map( A1 => C(13), A2 => n4, B1 => D(13), B2 => n1, ZN 
                           => n122);
   U152 : AOI22_X1 port map( A1 => A(13), A2 => n3, B1 => B(13), B2 => n2, ZN 
                           => n121);
   U153 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => Y(12));
   U154 : AOI22_X1 port map( A1 => G(12), A2 => n9, B1 => H(12), B2 => n10, ZN 
                           => n128);
   U155 : AOI22_X1 port map( A1 => E(12), A2 => n11, B1 => F(12), B2 => n12, ZN
                           => n127);
   U156 : AOI22_X1 port map( A1 => C(12), A2 => n4, B1 => D(12), B2 => n1, ZN 
                           => n126);
   U157 : AOI22_X1 port map( A1 => A(12), A2 => n3, B1 => B(12), B2 => n2, ZN 
                           => n125);
   U158 : NAND4_X1 port map( A1 => n129, A2 => n130, A3 => n131, A4 => n132, ZN
                           => Y(11));
   U159 : AOI22_X1 port map( A1 => G(11), A2 => n9, B1 => H(11), B2 => n10, ZN 
                           => n132);
   U160 : AOI22_X1 port map( A1 => E(11), A2 => n11, B1 => F(11), B2 => n12, ZN
                           => n131);
   U161 : AOI22_X1 port map( A1 => C(11), A2 => n4, B1 => D(11), B2 => n1, ZN 
                           => n130);
   U162 : AOI22_X1 port map( A1 => A(11), A2 => n3, B1 => B(11), B2 => n2, ZN 
                           => n129);
   U163 : NAND4_X1 port map( A1 => n133, A2 => n134, A3 => n135, A4 => n136, ZN
                           => Y(10));
   U164 : AOI22_X1 port map( A1 => G(10), A2 => n9, B1 => H(10), B2 => n10, ZN 
                           => n136);
   U165 : AOI22_X1 port map( A1 => E(10), A2 => n11, B1 => F(10), B2 => n12, ZN
                           => n135);
   U166 : AOI22_X1 port map( A1 => C(10), A2 => n4, B1 => D(10), B2 => n1, ZN 
                           => n134);
   U167 : AOI22_X1 port map( A1 => A(10), A2 => n3, B1 => B(10), B2 => n2, ZN 
                           => n133);
   U168 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => Y(0));
   U169 : AOI22_X1 port map( A1 => G(0), A2 => n9, B1 => H(0), B2 => n10, ZN =>
                           n140);
   U170 : AOI22_X1 port map( A1 => E(0), A2 => n11, B1 => F(0), B2 => n12, ZN 
                           => n139);
   U171 : AOI22_X1 port map( A1 => C(0), A2 => n4, B1 => D(0), B2 => n1, ZN => 
                           n138);
   U172 : INV_X1 port map( A => S(1), ZN => n142);
   U173 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => n2, ZN => 
                           n137);
   U174 : INV_X1 port map( A => S(0), ZN => n141);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_60;

architecture SYN_BEHAVIORAL of AND2_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_59;

architecture SYN_BEHAVIORAL of AND2_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_58;

architecture SYN_BEHAVIORAL of AND2_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_57;

architecture SYN_BEHAVIORAL of AND2_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_56;

architecture SYN_BEHAVIORAL of AND2_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_55;

architecture SYN_BEHAVIORAL of AND2_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_54;

architecture SYN_BEHAVIORAL of AND2_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_53;

architecture SYN_BEHAVIORAL of AND2_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_52;

architecture SYN_BEHAVIORAL of AND2_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_51;

architecture SYN_BEHAVIORAL of AND2_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_50;

architecture SYN_BEHAVIORAL of AND2_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_49;

architecture SYN_BEHAVIORAL of AND2_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_48;

architecture SYN_BEHAVIORAL of AND2_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_47;

architecture SYN_BEHAVIORAL of AND2_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_46;

architecture SYN_BEHAVIORAL of AND2_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_45;

architecture SYN_BEHAVIORAL of AND2_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_44;

architecture SYN_BEHAVIORAL of AND2_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_43;

architecture SYN_BEHAVIORAL of AND2_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_42;

architecture SYN_BEHAVIORAL of AND2_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_41;

architecture SYN_BEHAVIORAL of AND2_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_40;

architecture SYN_BEHAVIORAL of AND2_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_39;

architecture SYN_BEHAVIORAL of AND2_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_38;

architecture SYN_BEHAVIORAL of AND2_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_37;

architecture SYN_BEHAVIORAL of AND2_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_36;

architecture SYN_BEHAVIORAL of AND2_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_35;

architecture SYN_BEHAVIORAL of AND2_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_34;

architecture SYN_BEHAVIORAL of AND2_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_33;

architecture SYN_BEHAVIORAL of AND2_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_32;

architecture SYN_BEHAVIORAL of AND2_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_31;

architecture SYN_BEHAVIORAL of AND2_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_30;

architecture SYN_BEHAVIORAL of AND2_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_29;

architecture SYN_BEHAVIORAL of AND2_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_28;

architecture SYN_BEHAVIORAL of AND2_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_27;

architecture SYN_BEHAVIORAL of AND2_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_26;

architecture SYN_BEHAVIORAL of AND2_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_25;

architecture SYN_BEHAVIORAL of AND2_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_24;

architecture SYN_BEHAVIORAL of AND2_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_23;

architecture SYN_BEHAVIORAL of AND2_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_22;

architecture SYN_BEHAVIORAL of AND2_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_21;

architecture SYN_BEHAVIORAL of AND2_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_20;

architecture SYN_BEHAVIORAL of AND2_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_19;

architecture SYN_BEHAVIORAL of AND2_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_18;

architecture SYN_BEHAVIORAL of AND2_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_17;

architecture SYN_BEHAVIORAL of AND2_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_16;

architecture SYN_BEHAVIORAL of AND2_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_15;

architecture SYN_BEHAVIORAL of AND2_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_14;

architecture SYN_BEHAVIORAL of AND2_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_13;

architecture SYN_BEHAVIORAL of AND2_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_12;

architecture SYN_BEHAVIORAL of AND2_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_11;

architecture SYN_BEHAVIORAL of AND2_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_10;

architecture SYN_BEHAVIORAL of AND2_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_9;

architecture SYN_BEHAVIORAL of AND2_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_8;

architecture SYN_BEHAVIORAL of AND2_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_7;

architecture SYN_BEHAVIORAL of AND2_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_6;

architecture SYN_BEHAVIORAL of AND2_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_5;

architecture SYN_BEHAVIORAL of AND2_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_4;

architecture SYN_BEHAVIORAL of AND2_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_3;

architecture SYN_BEHAVIORAL of AND2_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_2;

architecture SYN_BEHAVIORAL of AND2_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_1;

architecture SYN_BEHAVIORAL of AND2_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_0;

architecture SYN_BEHAVIORAL of AND2_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_62;

architecture SYN_BEHAVIORAL of XNOR2_62 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_61;

architecture SYN_BEHAVIORAL of XNOR2_61 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_60;

architecture SYN_BEHAVIORAL of XNOR2_60 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_59;

architecture SYN_BEHAVIORAL of XNOR2_59 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_58;

architecture SYN_BEHAVIORAL of XNOR2_58 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_57;

architecture SYN_BEHAVIORAL of XNOR2_57 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_56;

architecture SYN_BEHAVIORAL of XNOR2_56 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_55;

architecture SYN_BEHAVIORAL of XNOR2_55 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_54;

architecture SYN_BEHAVIORAL of XNOR2_54 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_53;

architecture SYN_BEHAVIORAL of XNOR2_53 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_52;

architecture SYN_BEHAVIORAL of XNOR2_52 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_51;

architecture SYN_BEHAVIORAL of XNOR2_51 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_50;

architecture SYN_BEHAVIORAL of XNOR2_50 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_49;

architecture SYN_BEHAVIORAL of XNOR2_49 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_48;

architecture SYN_BEHAVIORAL of XNOR2_48 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_47;

architecture SYN_BEHAVIORAL of XNOR2_47 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_46;

architecture SYN_BEHAVIORAL of XNOR2_46 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_45;

architecture SYN_BEHAVIORAL of XNOR2_45 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_44;

architecture SYN_BEHAVIORAL of XNOR2_44 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_43;

architecture SYN_BEHAVIORAL of XNOR2_43 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_42;

architecture SYN_BEHAVIORAL of XNOR2_42 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_41;

architecture SYN_BEHAVIORAL of XNOR2_41 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_40;

architecture SYN_BEHAVIORAL of XNOR2_40 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_39;

architecture SYN_BEHAVIORAL of XNOR2_39 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_38;

architecture SYN_BEHAVIORAL of XNOR2_38 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_37;

architecture SYN_BEHAVIORAL of XNOR2_37 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_36;

architecture SYN_BEHAVIORAL of XNOR2_36 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_35;

architecture SYN_BEHAVIORAL of XNOR2_35 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_34;

architecture SYN_BEHAVIORAL of XNOR2_34 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_33;

architecture SYN_BEHAVIORAL of XNOR2_33 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_32;

architecture SYN_BEHAVIORAL of XNOR2_32 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_31;

architecture SYN_BEHAVIORAL of XNOR2_31 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_30;

architecture SYN_BEHAVIORAL of XNOR2_30 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_29;

architecture SYN_BEHAVIORAL of XNOR2_29 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_28;

architecture SYN_BEHAVIORAL of XNOR2_28 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_27;

architecture SYN_BEHAVIORAL of XNOR2_27 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_26;

architecture SYN_BEHAVIORAL of XNOR2_26 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_25;

architecture SYN_BEHAVIORAL of XNOR2_25 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_24;

architecture SYN_BEHAVIORAL of XNOR2_24 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_23;

architecture SYN_BEHAVIORAL of XNOR2_23 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_22;

architecture SYN_BEHAVIORAL of XNOR2_22 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_21;

architecture SYN_BEHAVIORAL of XNOR2_21 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_20;

architecture SYN_BEHAVIORAL of XNOR2_20 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_19;

architecture SYN_BEHAVIORAL of XNOR2_19 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_18;

architecture SYN_BEHAVIORAL of XNOR2_18 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_17;

architecture SYN_BEHAVIORAL of XNOR2_17 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_16;

architecture SYN_BEHAVIORAL of XNOR2_16 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_15;

architecture SYN_BEHAVIORAL of XNOR2_15 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_14;

architecture SYN_BEHAVIORAL of XNOR2_14 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_13;

architecture SYN_BEHAVIORAL of XNOR2_13 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_12;

architecture SYN_BEHAVIORAL of XNOR2_12 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_11;

architecture SYN_BEHAVIORAL of XNOR2_11 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_10;

architecture SYN_BEHAVIORAL of XNOR2_10 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_9;

architecture SYN_BEHAVIORAL of XNOR2_9 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_8;

architecture SYN_BEHAVIORAL of XNOR2_8 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_7;

architecture SYN_BEHAVIORAL of XNOR2_7 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_6;

architecture SYN_BEHAVIORAL of XNOR2_6 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_5;

architecture SYN_BEHAVIORAL of XNOR2_5 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_4;

architecture SYN_BEHAVIORAL of XNOR2_4 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_3;

architecture SYN_BEHAVIORAL of XNOR2_3 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_2;

architecture SYN_BEHAVIORAL of XNOR2_2 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_1;

architecture SYN_BEHAVIORAL of XNOR2_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_0;

architecture SYN_BEHAVIORAL of XNOR2_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_30 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_30;

architecture SYN_BEHAVIORAL of FFD_30 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1220 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1220);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_29 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_29;

architecture SYN_BEHAVIORAL of FFD_29 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1221 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1221);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_28 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_28;

architecture SYN_BEHAVIORAL of FFD_28 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1222 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1222);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_27 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_27;

architecture SYN_BEHAVIORAL of FFD_27 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1223 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1223);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_26 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_26;

architecture SYN_BEHAVIORAL of FFD_26 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1224 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1224);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_25 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_25;

architecture SYN_BEHAVIORAL of FFD_25 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1225 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1225);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_24 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_24;

architecture SYN_BEHAVIORAL of FFD_24 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1226 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1226);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_23 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_23;

architecture SYN_BEHAVIORAL of FFD_23 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1227 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1227);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_22 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_22;

architecture SYN_BEHAVIORAL of FFD_22 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1228 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1228);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_21 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_21;

architecture SYN_BEHAVIORAL of FFD_21 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1229 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1229);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_20 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_20;

architecture SYN_BEHAVIORAL of FFD_20 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1230 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1230);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_19 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_19;

architecture SYN_BEHAVIORAL of FFD_19 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1231 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1231);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_18 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_18;

architecture SYN_BEHAVIORAL of FFD_18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1232 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1232);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_17 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_17;

architecture SYN_BEHAVIORAL of FFD_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1233 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1233);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_16 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_16;

architecture SYN_BEHAVIORAL of FFD_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1234 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1234);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_15 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_15;

architecture SYN_BEHAVIORAL of FFD_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1235 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1235);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_14 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_14;

architecture SYN_BEHAVIORAL of FFD_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1236 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1236);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_13 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_13;

architecture SYN_BEHAVIORAL of FFD_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1237 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1237);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_12 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_12;

architecture SYN_BEHAVIORAL of FFD_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1238 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1238);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_11 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_11;

architecture SYN_BEHAVIORAL of FFD_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1239 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1239);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_10 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_10;

architecture SYN_BEHAVIORAL of FFD_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1240 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1240);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_9 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_9;

architecture SYN_BEHAVIORAL of FFD_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1241 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1241);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_8 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_8;

architecture SYN_BEHAVIORAL of FFD_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1242 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1242);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_7 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_7;

architecture SYN_BEHAVIORAL of FFD_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1243 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1243);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_6 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_6;

architecture SYN_BEHAVIORAL of FFD_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1244 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1244);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_5 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_5;

architecture SYN_BEHAVIORAL of FFD_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1245 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1245);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_4 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_4;

architecture SYN_BEHAVIORAL of FFD_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1246 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1246);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_3 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_3;

architecture SYN_BEHAVIORAL of FFD_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1247 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1247);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_2 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_2;

architecture SYN_BEHAVIORAL of FFD_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1248 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1248);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_1 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_1;

architecture SYN_BEHAVIORAL of FFD_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1249 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1249);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_0 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_0;

architecture SYN_BEHAVIORAL of FFD_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1250 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1250);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n2);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_223 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_223;

architecture SYN_BEHAVIORAL of LD_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_222 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_222;

architecture SYN_BEHAVIORAL of LD_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_221 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_221;

architecture SYN_BEHAVIORAL of LD_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_220 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_220;

architecture SYN_BEHAVIORAL of LD_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_219 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_219;

architecture SYN_BEHAVIORAL of LD_219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_218 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_218;

architecture SYN_BEHAVIORAL of LD_218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_217 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_217;

architecture SYN_BEHAVIORAL of LD_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_216 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_216;

architecture SYN_BEHAVIORAL of LD_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_215 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_215;

architecture SYN_BEHAVIORAL of LD_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_214 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_214;

architecture SYN_BEHAVIORAL of LD_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_213 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_213;

architecture SYN_BEHAVIORAL of LD_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_212 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_212;

architecture SYN_BEHAVIORAL of LD_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_211 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_211;

architecture SYN_BEHAVIORAL of LD_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_210 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_210;

architecture SYN_BEHAVIORAL of LD_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_209 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_209;

architecture SYN_BEHAVIORAL of LD_209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_208 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_208;

architecture SYN_BEHAVIORAL of LD_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_207 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_207;

architecture SYN_BEHAVIORAL of LD_207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_206 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_206;

architecture SYN_BEHAVIORAL of LD_206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_205 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_205;

architecture SYN_BEHAVIORAL of LD_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_204 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_204;

architecture SYN_BEHAVIORAL of LD_204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_203 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_203;

architecture SYN_BEHAVIORAL of LD_203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_202 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_202;

architecture SYN_BEHAVIORAL of LD_202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_201 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_201;

architecture SYN_BEHAVIORAL of LD_201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_200 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_200;

architecture SYN_BEHAVIORAL of LD_200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_199 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_199;

architecture SYN_BEHAVIORAL of LD_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_198 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_198;

architecture SYN_BEHAVIORAL of LD_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_197 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_197;

architecture SYN_BEHAVIORAL of LD_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_196 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_196;

architecture SYN_BEHAVIORAL of LD_196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_195 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_195;

architecture SYN_BEHAVIORAL of LD_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_194 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_194;

architecture SYN_BEHAVIORAL of LD_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_193 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_193;

architecture SYN_BEHAVIORAL of LD_193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_192 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_192;

architecture SYN_BEHAVIORAL of LD_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_191 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_191;

architecture SYN_BEHAVIORAL of LD_191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_190 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_190;

architecture SYN_BEHAVIORAL of LD_190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_189 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_189;

architecture SYN_BEHAVIORAL of LD_189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_188 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_188;

architecture SYN_BEHAVIORAL of LD_188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_187 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_187;

architecture SYN_BEHAVIORAL of LD_187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_186 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_186;

architecture SYN_BEHAVIORAL of LD_186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_185 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_185;

architecture SYN_BEHAVIORAL of LD_185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_184 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_184;

architecture SYN_BEHAVIORAL of LD_184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_183 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_183;

architecture SYN_BEHAVIORAL of LD_183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_182 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_182;

architecture SYN_BEHAVIORAL of LD_182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_181 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_181;

architecture SYN_BEHAVIORAL of LD_181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_180 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_180;

architecture SYN_BEHAVIORAL of LD_180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_179 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_179;

architecture SYN_BEHAVIORAL of LD_179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_178 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_178;

architecture SYN_BEHAVIORAL of LD_178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_177 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_177;

architecture SYN_BEHAVIORAL of LD_177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_176 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_176;

architecture SYN_BEHAVIORAL of LD_176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_175 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_175;

architecture SYN_BEHAVIORAL of LD_175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_174 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_174;

architecture SYN_BEHAVIORAL of LD_174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_173 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_173;

architecture SYN_BEHAVIORAL of LD_173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_172 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_172;

architecture SYN_BEHAVIORAL of LD_172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_171 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_171;

architecture SYN_BEHAVIORAL of LD_171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_170 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_170;

architecture SYN_BEHAVIORAL of LD_170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_169 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_169;

architecture SYN_BEHAVIORAL of LD_169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_168 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_168;

architecture SYN_BEHAVIORAL of LD_168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_167 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_167;

architecture SYN_BEHAVIORAL of LD_167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_166 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_166;

architecture SYN_BEHAVIORAL of LD_166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_165 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_165;

architecture SYN_BEHAVIORAL of LD_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_164 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_164;

architecture SYN_BEHAVIORAL of LD_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_163 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_163;

architecture SYN_BEHAVIORAL of LD_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_162 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_162;

architecture SYN_BEHAVIORAL of LD_162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_161 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_161;

architecture SYN_BEHAVIORAL of LD_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_160 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_160;

architecture SYN_BEHAVIORAL of LD_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_159 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_159;

architecture SYN_BEHAVIORAL of LD_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_158 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_158;

architecture SYN_BEHAVIORAL of LD_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_157 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_157;

architecture SYN_BEHAVIORAL of LD_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_156 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_156;

architecture SYN_BEHAVIORAL of LD_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_155 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_155;

architecture SYN_BEHAVIORAL of LD_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_154 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_154;

architecture SYN_BEHAVIORAL of LD_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_153 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_153;

architecture SYN_BEHAVIORAL of LD_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_152 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_152;

architecture SYN_BEHAVIORAL of LD_152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_151 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_151;

architecture SYN_BEHAVIORAL of LD_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_150 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_150;

architecture SYN_BEHAVIORAL of LD_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_149 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_149;

architecture SYN_BEHAVIORAL of LD_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_148 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_148;

architecture SYN_BEHAVIORAL of LD_148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_147 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_147;

architecture SYN_BEHAVIORAL of LD_147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_146 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_146;

architecture SYN_BEHAVIORAL of LD_146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_145 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_145;

architecture SYN_BEHAVIORAL of LD_145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_144 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_144;

architecture SYN_BEHAVIORAL of LD_144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_143 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_143;

architecture SYN_BEHAVIORAL of LD_143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_142 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_142;

architecture SYN_BEHAVIORAL of LD_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_141 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_141;

architecture SYN_BEHAVIORAL of LD_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_140 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_140;

architecture SYN_BEHAVIORAL of LD_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_139 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_139;

architecture SYN_BEHAVIORAL of LD_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_138 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_138;

architecture SYN_BEHAVIORAL of LD_138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_137 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_137;

architecture SYN_BEHAVIORAL of LD_137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_136 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_136;

architecture SYN_BEHAVIORAL of LD_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_135 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_135;

architecture SYN_BEHAVIORAL of LD_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_134 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_134;

architecture SYN_BEHAVIORAL of LD_134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_133 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_133;

architecture SYN_BEHAVIORAL of LD_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_132 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_132;

architecture SYN_BEHAVIORAL of LD_132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_131 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_131;

architecture SYN_BEHAVIORAL of LD_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_130 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_130;

architecture SYN_BEHAVIORAL of LD_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_129 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_129;

architecture SYN_BEHAVIORAL of LD_129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_128 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_128;

architecture SYN_BEHAVIORAL of LD_128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_127 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_127;

architecture SYN_BEHAVIORAL of LD_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_126 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_126;

architecture SYN_BEHAVIORAL of LD_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_125 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_125;

architecture SYN_BEHAVIORAL of LD_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_124 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_124;

architecture SYN_BEHAVIORAL of LD_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_123 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_123;

architecture SYN_BEHAVIORAL of LD_123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_122 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_122;

architecture SYN_BEHAVIORAL of LD_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_121 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_121;

architecture SYN_BEHAVIORAL of LD_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_120 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_120;

architecture SYN_BEHAVIORAL of LD_120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_119 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_119;

architecture SYN_BEHAVIORAL of LD_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_118 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_118;

architecture SYN_BEHAVIORAL of LD_118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_117 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_117;

architecture SYN_BEHAVIORAL of LD_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_116 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_116;

architecture SYN_BEHAVIORAL of LD_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_115 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_115;

architecture SYN_BEHAVIORAL of LD_115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_114 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_114;

architecture SYN_BEHAVIORAL of LD_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_113 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_113;

architecture SYN_BEHAVIORAL of LD_113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_112 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_112;

architecture SYN_BEHAVIORAL of LD_112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_111 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_111;

architecture SYN_BEHAVIORAL of LD_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_110 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_110;

architecture SYN_BEHAVIORAL of LD_110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_109 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_109;

architecture SYN_BEHAVIORAL of LD_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_108 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_108;

architecture SYN_BEHAVIORAL of LD_108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_107 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_107;

architecture SYN_BEHAVIORAL of LD_107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_106 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_106;

architecture SYN_BEHAVIORAL of LD_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_105 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_105;

architecture SYN_BEHAVIORAL of LD_105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_104 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_104;

architecture SYN_BEHAVIORAL of LD_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_103 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_103;

architecture SYN_BEHAVIORAL of LD_103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_102 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_102;

architecture SYN_BEHAVIORAL of LD_102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_101 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_101;

architecture SYN_BEHAVIORAL of LD_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_100 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_100;

architecture SYN_BEHAVIORAL of LD_100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_99 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_99;

architecture SYN_BEHAVIORAL of LD_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_98 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_98;

architecture SYN_BEHAVIORAL of LD_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_97 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_97;

architecture SYN_BEHAVIORAL of LD_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_96 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_96;

architecture SYN_BEHAVIORAL of LD_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_95 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_95;

architecture SYN_BEHAVIORAL of LD_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_94 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_94;

architecture SYN_BEHAVIORAL of LD_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_93 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_93;

architecture SYN_BEHAVIORAL of LD_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_92 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_92;

architecture SYN_BEHAVIORAL of LD_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_91 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_91;

architecture SYN_BEHAVIORAL of LD_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_90 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_90;

architecture SYN_BEHAVIORAL of LD_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_89 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_89;

architecture SYN_BEHAVIORAL of LD_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_88 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_88;

architecture SYN_BEHAVIORAL of LD_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_87 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_87;

architecture SYN_BEHAVIORAL of LD_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_86 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_86;

architecture SYN_BEHAVIORAL of LD_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_85 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_85;

architecture SYN_BEHAVIORAL of LD_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_84 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_84;

architecture SYN_BEHAVIORAL of LD_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_83 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_83;

architecture SYN_BEHAVIORAL of LD_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_82 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_82;

architecture SYN_BEHAVIORAL of LD_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_81 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_81;

architecture SYN_BEHAVIORAL of LD_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_80 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_80;

architecture SYN_BEHAVIORAL of LD_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_79 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_79;

architecture SYN_BEHAVIORAL of LD_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_78 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_78;

architecture SYN_BEHAVIORAL of LD_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_77 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_77;

architecture SYN_BEHAVIORAL of LD_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_76 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_76;

architecture SYN_BEHAVIORAL of LD_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_75 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_75;

architecture SYN_BEHAVIORAL of LD_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_74 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_74;

architecture SYN_BEHAVIORAL of LD_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_73 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_73;

architecture SYN_BEHAVIORAL of LD_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_72 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_72;

architecture SYN_BEHAVIORAL of LD_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_71 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_71;

architecture SYN_BEHAVIORAL of LD_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_70 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_70;

architecture SYN_BEHAVIORAL of LD_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_69 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_69;

architecture SYN_BEHAVIORAL of LD_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_68 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_68;

architecture SYN_BEHAVIORAL of LD_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_67 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_67;

architecture SYN_BEHAVIORAL of LD_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_66 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_66;

architecture SYN_BEHAVIORAL of LD_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_65 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_65;

architecture SYN_BEHAVIORAL of LD_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_64 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_64;

architecture SYN_BEHAVIORAL of LD_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_63 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_63;

architecture SYN_BEHAVIORAL of LD_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_62 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_62;

architecture SYN_BEHAVIORAL of LD_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_61 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_61;

architecture SYN_BEHAVIORAL of LD_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_60 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_60;

architecture SYN_BEHAVIORAL of LD_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_59 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_59;

architecture SYN_BEHAVIORAL of LD_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_58 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_58;

architecture SYN_BEHAVIORAL of LD_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_57 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_57;

architecture SYN_BEHAVIORAL of LD_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_56 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_56;

architecture SYN_BEHAVIORAL of LD_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_55 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_55;

architecture SYN_BEHAVIORAL of LD_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_54 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_54;

architecture SYN_BEHAVIORAL of LD_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_53 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_53;

architecture SYN_BEHAVIORAL of LD_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_52 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_52;

architecture SYN_BEHAVIORAL of LD_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_51 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_51;

architecture SYN_BEHAVIORAL of LD_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_50 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_50;

architecture SYN_BEHAVIORAL of LD_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_49 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_49;

architecture SYN_BEHAVIORAL of LD_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_48 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_48;

architecture SYN_BEHAVIORAL of LD_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_47 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_47;

architecture SYN_BEHAVIORAL of LD_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_46 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_46;

architecture SYN_BEHAVIORAL of LD_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_45 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_45;

architecture SYN_BEHAVIORAL of LD_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_44 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_44;

architecture SYN_BEHAVIORAL of LD_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_43 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_43;

architecture SYN_BEHAVIORAL of LD_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_42 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_42;

architecture SYN_BEHAVIORAL of LD_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_41 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_41;

architecture SYN_BEHAVIORAL of LD_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_40 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_40;

architecture SYN_BEHAVIORAL of LD_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_39 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_39;

architecture SYN_BEHAVIORAL of LD_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_38 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_38;

architecture SYN_BEHAVIORAL of LD_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_37 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_37;

architecture SYN_BEHAVIORAL of LD_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_36 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_36;

architecture SYN_BEHAVIORAL of LD_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_35 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_35;

architecture SYN_BEHAVIORAL of LD_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_34 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_34;

architecture SYN_BEHAVIORAL of LD_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_33 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_33;

architecture SYN_BEHAVIORAL of LD_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_32 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_32;

architecture SYN_BEHAVIORAL of LD_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_31 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_31;

architecture SYN_BEHAVIORAL of LD_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_30 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_30;

architecture SYN_BEHAVIORAL of LD_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_29 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_29;

architecture SYN_BEHAVIORAL of LD_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_28 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_28;

architecture SYN_BEHAVIORAL of LD_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_27 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_27;

architecture SYN_BEHAVIORAL of LD_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_26 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_26;

architecture SYN_BEHAVIORAL of LD_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_25 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_25;

architecture SYN_BEHAVIORAL of LD_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_24 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_24;

architecture SYN_BEHAVIORAL of LD_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_23 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_23;

architecture SYN_BEHAVIORAL of LD_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_22 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_22;

architecture SYN_BEHAVIORAL of LD_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_21 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_21;

architecture SYN_BEHAVIORAL of LD_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_20 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_20;

architecture SYN_BEHAVIORAL of LD_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_19 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_19;

architecture SYN_BEHAVIORAL of LD_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_18 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_18;

architecture SYN_BEHAVIORAL of LD_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_17 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_17;

architecture SYN_BEHAVIORAL of LD_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_16 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_16;

architecture SYN_BEHAVIORAL of LD_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_15 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_15;

architecture SYN_BEHAVIORAL of LD_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_14 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_14;

architecture SYN_BEHAVIORAL of LD_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_13 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_13;

architecture SYN_BEHAVIORAL of LD_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_12 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_12;

architecture SYN_BEHAVIORAL of LD_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_11 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_11;

architecture SYN_BEHAVIORAL of LD_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_10 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_10;

architecture SYN_BEHAVIORAL of LD_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_9 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_9;

architecture SYN_BEHAVIORAL of LD_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_8 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_8;

architecture SYN_BEHAVIORAL of LD_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_7 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_7;

architecture SYN_BEHAVIORAL of LD_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_6 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_6;

architecture SYN_BEHAVIORAL of LD_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_5 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_5;

architecture SYN_BEHAVIORAL of LD_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_4 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_4;

architecture SYN_BEHAVIORAL of LD_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_3 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_3;

architecture SYN_BEHAVIORAL of LD_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_2 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_2;

architecture SYN_BEHAVIORAL of LD_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_1 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_1;

architecture SYN_BEHAVIORAL of LD_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_0 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_0;

architecture SYN_BEHAVIORAL of LD_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX41_N32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX41_N32_0;

architecture SYN_BEHAVIORAL of MUX41_N32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n1);
   U2 : OR2_X1 port map( A1 => n71, A2 => S(1), ZN => n2);
   U3 : INV_X2 port map( A => n2, ZN => n3);
   U4 : INV_X2 port map( A => n1, ZN => n4);
   U5 : AND2_X2 port map( A1 => S(0), A2 => S(1), ZN => n8);
   U6 : AND2_X2 port map( A1 => S(1), A2 => n71, ZN => n7);
   U7 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Y(9));
   U8 : AOI22_X1 port map( A1 => C(9), A2 => n7, B1 => D(9), B2 => n8, ZN => n6
                           );
   U9 : AOI22_X1 port map( A1 => A(9), A2 => n4, B1 => B(9), B2 => n3, ZN => n5
                           );
   U10 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => Y(8));
   U11 : AOI22_X1 port map( A1 => C(8), A2 => n7, B1 => D(8), B2 => n8, ZN => 
                           n10);
   U12 : AOI22_X1 port map( A1 => A(8), A2 => n4, B1 => B(8), B2 => n3, ZN => 
                           n9);
   U13 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => Y(7));
   U14 : AOI22_X1 port map( A1 => C(7), A2 => n7, B1 => D(7), B2 => n8, ZN => 
                           n12);
   U15 : AOI22_X1 port map( A1 => A(7), A2 => n4, B1 => B(7), B2 => n3, ZN => 
                           n11);
   U16 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => Y(6));
   U17 : AOI22_X1 port map( A1 => C(6), A2 => n7, B1 => D(6), B2 => n8, ZN => 
                           n14);
   U18 : AOI22_X1 port map( A1 => A(6), A2 => n4, B1 => B(6), B2 => n3, ZN => 
                           n13);
   U19 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => Y(5));
   U20 : AOI22_X1 port map( A1 => C(5), A2 => n7, B1 => D(5), B2 => n8, ZN => 
                           n16);
   U21 : AOI22_X1 port map( A1 => A(5), A2 => n4, B1 => B(5), B2 => n3, ZN => 
                           n15);
   U22 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => Y(4));
   U23 : AOI22_X1 port map( A1 => C(4), A2 => n7, B1 => D(4), B2 => n8, ZN => 
                           n18);
   U24 : AOI22_X1 port map( A1 => A(4), A2 => n4, B1 => B(4), B2 => n3, ZN => 
                           n17);
   U25 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => Y(3));
   U26 : AOI22_X1 port map( A1 => C(3), A2 => n7, B1 => D(3), B2 => n8, ZN => 
                           n20);
   U27 : AOI22_X1 port map( A1 => A(3), A2 => n4, B1 => B(3), B2 => n3, ZN => 
                           n19);
   U28 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => Y(31));
   U29 : AOI22_X1 port map( A1 => C(31), A2 => n7, B1 => D(31), B2 => n8, ZN =>
                           n22);
   U30 : AOI22_X1 port map( A1 => A(31), A2 => n4, B1 => B(31), B2 => n3, ZN =>
                           n21);
   U31 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => Y(30));
   U32 : AOI22_X1 port map( A1 => C(30), A2 => n7, B1 => D(30), B2 => n8, ZN =>
                           n24);
   U33 : AOI22_X1 port map( A1 => A(30), A2 => n4, B1 => B(30), B2 => n3, ZN =>
                           n23);
   U34 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => Y(2));
   U35 : AOI22_X1 port map( A1 => C(2), A2 => n7, B1 => D(2), B2 => n8, ZN => 
                           n26);
   U36 : AOI22_X1 port map( A1 => A(2), A2 => n4, B1 => B(2), B2 => n3, ZN => 
                           n25);
   U37 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => Y(29));
   U38 : AOI22_X1 port map( A1 => C(29), A2 => n7, B1 => D(29), B2 => n8, ZN =>
                           n28);
   U39 : AOI22_X1 port map( A1 => A(29), A2 => n4, B1 => B(29), B2 => n3, ZN =>
                           n27);
   U40 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => Y(28));
   U41 : AOI22_X1 port map( A1 => C(28), A2 => n7, B1 => D(28), B2 => n8, ZN =>
                           n30);
   U42 : AOI22_X1 port map( A1 => A(28), A2 => n4, B1 => B(28), B2 => n3, ZN =>
                           n29);
   U43 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => Y(27));
   U44 : AOI22_X1 port map( A1 => C(27), A2 => n7, B1 => D(27), B2 => n8, ZN =>
                           n32);
   U45 : AOI22_X1 port map( A1 => A(27), A2 => n4, B1 => B(27), B2 => n3, ZN =>
                           n31);
   U46 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => Y(26));
   U47 : AOI22_X1 port map( A1 => C(26), A2 => n7, B1 => D(26), B2 => n8, ZN =>
                           n34);
   U48 : AOI22_X1 port map( A1 => A(26), A2 => n4, B1 => B(26), B2 => n3, ZN =>
                           n33);
   U49 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => Y(25));
   U50 : AOI22_X1 port map( A1 => C(25), A2 => n7, B1 => D(25), B2 => n8, ZN =>
                           n36);
   U51 : AOI22_X1 port map( A1 => A(25), A2 => n4, B1 => B(25), B2 => n3, ZN =>
                           n35);
   U52 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => Y(24));
   U53 : AOI22_X1 port map( A1 => C(24), A2 => n7, B1 => D(24), B2 => n8, ZN =>
                           n38);
   U54 : AOI22_X1 port map( A1 => A(24), A2 => n4, B1 => B(24), B2 => n3, ZN =>
                           n37);
   U55 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => Y(23));
   U56 : AOI22_X1 port map( A1 => C(23), A2 => n7, B1 => D(23), B2 => n8, ZN =>
                           n40);
   U57 : AOI22_X1 port map( A1 => A(23), A2 => n4, B1 => B(23), B2 => n3, ZN =>
                           n39);
   U58 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => Y(22));
   U59 : AOI22_X1 port map( A1 => C(22), A2 => n7, B1 => D(22), B2 => n8, ZN =>
                           n42);
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n4, B1 => B(22), B2 => n3, ZN =>
                           n41);
   U61 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => Y(21));
   U62 : AOI22_X1 port map( A1 => C(21), A2 => n7, B1 => D(21), B2 => n8, ZN =>
                           n44);
   U63 : AOI22_X1 port map( A1 => A(21), A2 => n4, B1 => B(21), B2 => n3, ZN =>
                           n43);
   U64 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => Y(20));
   U65 : AOI22_X1 port map( A1 => C(20), A2 => n7, B1 => D(20), B2 => n8, ZN =>
                           n46);
   U66 : AOI22_X1 port map( A1 => A(20), A2 => n4, B1 => B(20), B2 => n3, ZN =>
                           n45);
   U67 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => Y(1));
   U68 : AOI22_X1 port map( A1 => C(1), A2 => n7, B1 => D(1), B2 => n8, ZN => 
                           n48);
   U69 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n3, ZN => 
                           n47);
   U70 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => Y(19));
   U71 : AOI22_X1 port map( A1 => C(19), A2 => n7, B1 => D(19), B2 => n8, ZN =>
                           n50);
   U72 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n3, ZN =>
                           n49);
   U73 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => Y(18));
   U74 : AOI22_X1 port map( A1 => C(18), A2 => n7, B1 => D(18), B2 => n8, ZN =>
                           n52);
   U75 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n3, ZN =>
                           n51);
   U76 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => Y(17));
   U77 : AOI22_X1 port map( A1 => C(17), A2 => n7, B1 => D(17), B2 => n8, ZN =>
                           n54);
   U78 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n3, ZN =>
                           n53);
   U79 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => Y(16));
   U80 : AOI22_X1 port map( A1 => C(16), A2 => n7, B1 => D(16), B2 => n8, ZN =>
                           n56);
   U81 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n3, ZN =>
                           n55);
   U82 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => Y(15));
   U83 : AOI22_X1 port map( A1 => C(15), A2 => n7, B1 => D(15), B2 => n8, ZN =>
                           n58);
   U84 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n3, ZN =>
                           n57);
   U85 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => Y(14));
   U86 : AOI22_X1 port map( A1 => C(14), A2 => n7, B1 => D(14), B2 => n8, ZN =>
                           n60);
   U87 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n3, ZN =>
                           n59);
   U88 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => Y(13));
   U89 : AOI22_X1 port map( A1 => C(13), A2 => n7, B1 => D(13), B2 => n8, ZN =>
                           n62);
   U90 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n3, ZN =>
                           n61);
   U91 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => Y(12));
   U92 : AOI22_X1 port map( A1 => C(12), A2 => n7, B1 => D(12), B2 => n8, ZN =>
                           n64);
   U93 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n3, ZN =>
                           n63);
   U94 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => Y(11));
   U95 : AOI22_X1 port map( A1 => C(11), A2 => n7, B1 => D(11), B2 => n8, ZN =>
                           n66);
   U96 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n3, ZN =>
                           n65);
   U97 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => Y(10));
   U98 : AOI22_X1 port map( A1 => C(10), A2 => n7, B1 => D(10), B2 => n8, ZN =>
                           n68);
   U99 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n3, ZN =>
                           n67);
   U100 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => Y(0));
   U101 : AOI22_X1 port map( A1 => C(0), A2 => n7, B1 => D(0), B2 => n8, ZN => 
                           n70);
   U102 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n3, ZN => 
                           n69);
   U103 : INV_X1 port map( A => S(0), ZN => n71);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_5 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_5;

architecture SYN_STRUCTURAL of LDR_N32_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_160
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_161
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_162
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_163
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_164
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_165
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_166
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_167
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_168
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_169
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_170
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_171
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_172
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_173
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_174
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_175
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_176
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_177
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_178
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_179
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_180
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_181
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_182
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_183
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_184
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_185
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_186
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_187
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_188
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_189
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_190
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_191
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_191 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_190 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_189 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_188 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_187 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_186 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_185 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_184 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_183 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_182 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_181 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_180 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_179 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_178 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_177 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_176 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_175 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_174 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_173 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_172 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_171 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_170 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_169 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9))
                           ;
   LDI_8 : LD_168 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8))
                           ;
   LDI_7 : LD_167 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7))
                           ;
   LDI_6 : LD_166 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6))
                           ;
   LDI_5 : LD_165 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5))
                           ;
   LDI_4 : LD_164 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4))
                           ;
   LDI_3 : LD_163 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3))
                           ;
   LDI_2 : LD_162 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2))
                           ;
   LDI_1 : LD_161 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1))
                           ;
   LDI_0 : LD_160 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0))
                           ;
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_4 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_4;

architecture SYN_STRUCTURAL of LDR_N32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_128
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_129
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_130
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_131
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_132
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_133
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_134
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_135
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_136
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_137
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_138
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_139
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_140
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_141
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_142
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_143
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_144
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_145
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_146
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_147
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_148
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_149
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_150
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_151
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_152
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_153
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_154
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_155
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_156
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_157
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_158
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_159
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_159 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_158 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_157 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_156 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_155 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_154 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_153 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_152 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_151 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_150 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_149 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_148 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_147 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_146 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_145 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_144 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_143 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_142 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_141 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_140 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_139 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_138 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_137 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9))
                           ;
   LDI_8 : LD_136 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8))
                           ;
   LDI_7 : LD_135 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7))
                           ;
   LDI_6 : LD_134 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6))
                           ;
   LDI_5 : LD_133 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5))
                           ;
   LDI_4 : LD_132 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4))
                           ;
   LDI_3 : LD_131 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3))
                           ;
   LDI_2 : LD_130 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2))
                           ;
   LDI_1 : LD_129 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1))
                           ;
   LDI_0 : LD_128 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0))
                           ;
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_3 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_3;

architecture SYN_STRUCTURAL of LDR_N32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_96
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_97
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_98
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_99
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_100
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_101
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_102
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_103
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_104
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_105
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_106
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_107
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_108
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_109
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_110
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_111
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_112
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_113
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_114
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_115
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_116
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_117
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_118
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_119
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_120
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_121
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_122
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_123
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_124
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_125
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_126
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_127
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_127 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_126 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_125 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_124 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_123 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_122 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_121 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_120 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_119 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_118 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_117 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_116 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_115 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_114 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_113 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_112 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_111 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_110 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_109 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_108 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_107 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_106 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_105 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9))
                           ;
   LDI_8 : LD_104 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8))
                           ;
   LDI_7 : LD_103 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7))
                           ;
   LDI_6 : LD_102 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6))
                           ;
   LDI_5 : LD_101 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5))
                           ;
   LDI_4 : LD_100 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4))
                           ;
   LDI_3 : LD_99 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3));
   LDI_2 : LD_98 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2));
   LDI_1 : LD_97 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1));
   LDI_0 : LD_96 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_2 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_2;

architecture SYN_STRUCTURAL of LDR_N32_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_64
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_65
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_66
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_67
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_68
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_69
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_70
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_71
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_72
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_73
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_74
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_75
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_76
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_77
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_78
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_79
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_80
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_81
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_82
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_83
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_84
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_85
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_86
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_87
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_88
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_89
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_90
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_91
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_92
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_93
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_94
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_95
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_95 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_94 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_93 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_92 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_91 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_90 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_89 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_88 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_87 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_86 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_85 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_84 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_83 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_82 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_81 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_80 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_79 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_78 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_77 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_76 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_75 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_74 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_73 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9));
   LDI_8 : LD_72 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8));
   LDI_7 : LD_71 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7));
   LDI_6 : LD_70 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6));
   LDI_5 : LD_69 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5));
   LDI_4 : LD_68 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4));
   LDI_3 : LD_67 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3));
   LDI_2 : LD_66 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2));
   LDI_1 : LD_65 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1));
   LDI_0 : LD_64 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_1 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_1;

architecture SYN_STRUCTURAL of LDR_N32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_32
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_33
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_34
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_35
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_36
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_37
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_38
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_39
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_40
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_41
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_42
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_43
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_44
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_45
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_46
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_47
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_48
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_49
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_50
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_51
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_52
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_53
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_54
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_55
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_56
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_57
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_58
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_59
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_60
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_61
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_62
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_63
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_63 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_62 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_61 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_60 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_59 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_58 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_57 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_56 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_55 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_54 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_53 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_52 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_51 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_50 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_49 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_48 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_47 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_46 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_45 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_44 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_43 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_42 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_41 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9));
   LDI_8 : LD_40 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8));
   LDI_7 : LD_39 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7));
   LDI_6 : LD_38 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6));
   LDI_5 : LD_37 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5));
   LDI_4 : LD_36 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4));
   LDI_3 : LD_35 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3));
   LDI_2 : LD_34 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2));
   LDI_1 : LD_33 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1));
   LDI_0 : LD_32 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_0 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_0;

architecture SYN_STRUCTURAL of LDR_N32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_0
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_1
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_2
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_3
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_4
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_5
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_6
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_7
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_8
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_9
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_10
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_11
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_12
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_13
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_14
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_15
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_16
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_17
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_18
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_19
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_20
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_21
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_22
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_23
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_24
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_25
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_26
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_27
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_28
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_29
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_30
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_31
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_31 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_30 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_29 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_28 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_27 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_26 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_25 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_24 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_23 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_22 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_21 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_20 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_19 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_18 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_17 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_16 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_15 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_14 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_13 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_12 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_11 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_10 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_9 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9));
   LDI_8 : LD_8 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8));
   LDI_7 : LD_7 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7));
   LDI_6 : LD_6 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6));
   LDI_5 : LD_5 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5));
   LDI_4 : LD_4 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4));
   LDI_3 : LD_3 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3));
   LDI_2 : LD_2 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2));
   LDI_1 : LD_1 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1));
   LDI_0 : LD_0 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_3;

architecture SYN_BEHAVIORAL of MUX21_N32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => S, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => S, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => S, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => S, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => S, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => S, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => S, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => S, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => S, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => S, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => S, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => S, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => S, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => S, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => S, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => S, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => S, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => S, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => S, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => S, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => S, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => S, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => S, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => S, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => S, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => S, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => S, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => S, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_2;

architecture SYN_BEHAVIORAL of MUX21_N32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => S, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => S, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => S, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => S, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => S, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => S, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => S, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => S, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => S, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => S, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => S, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => S, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => S, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => S, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => S, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => S, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => S, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => S, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => S, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => S, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => S, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => S, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => S, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => S, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => S, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => S, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => S, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => S, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_1;

architecture SYN_BEHAVIORAL of MUX21_N32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => S, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => S, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => S, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => S, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => S, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => S, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => S, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => S, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => S, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => S, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => S, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => S, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => S, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => S, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => S, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => S, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => S, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => S, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => S, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => S, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => S, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => S, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => S, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => S, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => S, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => S, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => S, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => S, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_0;

architecture SYN_BEHAVIORAL of MUX21_N32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => S, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => S, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => S, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => S, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => S, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => S, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => S, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => S, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => S, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => S, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => S, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => S, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => S, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => S, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => S, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => S, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => S, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => S, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => S, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => S, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => S, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => S, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => S, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => S, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => S, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => S, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => S, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => S, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_319 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_319;

architecture SYN_BEHAVIORAL of MUX21_L_319 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_318 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_318;

architecture SYN_BEHAVIORAL of MUX21_L_318 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_317 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_317;

architecture SYN_BEHAVIORAL of MUX21_L_317 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_316 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_316;

architecture SYN_BEHAVIORAL of MUX21_L_316 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_315 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_315;

architecture SYN_BEHAVIORAL of MUX21_L_315 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_314 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_314;

architecture SYN_BEHAVIORAL of MUX21_L_314 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_313 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_313;

architecture SYN_BEHAVIORAL of MUX21_L_313 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_312 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_312;

architecture SYN_BEHAVIORAL of MUX21_L_312 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_311 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_311;

architecture SYN_BEHAVIORAL of MUX21_L_311 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_310 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_310;

architecture SYN_BEHAVIORAL of MUX21_L_310 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_309 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_309;

architecture SYN_BEHAVIORAL of MUX21_L_309 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_308 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_308;

architecture SYN_BEHAVIORAL of MUX21_L_308 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_307 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_307;

architecture SYN_BEHAVIORAL of MUX21_L_307 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_306 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_306;

architecture SYN_BEHAVIORAL of MUX21_L_306 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_305 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_305;

architecture SYN_BEHAVIORAL of MUX21_L_305 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_304 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_304;

architecture SYN_BEHAVIORAL of MUX21_L_304 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_303 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_303;

architecture SYN_BEHAVIORAL of MUX21_L_303 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_302 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_302;

architecture SYN_BEHAVIORAL of MUX21_L_302 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_301 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_301;

architecture SYN_BEHAVIORAL of MUX21_L_301 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_300 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_300;

architecture SYN_BEHAVIORAL of MUX21_L_300 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_299 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_299;

architecture SYN_BEHAVIORAL of MUX21_L_299 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_298 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_298;

architecture SYN_BEHAVIORAL of MUX21_L_298 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_297 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_297;

architecture SYN_BEHAVIORAL of MUX21_L_297 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_296 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_296;

architecture SYN_BEHAVIORAL of MUX21_L_296 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_295 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_295;

architecture SYN_BEHAVIORAL of MUX21_L_295 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_294 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_294;

architecture SYN_BEHAVIORAL of MUX21_L_294 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_293 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_293;

architecture SYN_BEHAVIORAL of MUX21_L_293 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_292 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_292;

architecture SYN_BEHAVIORAL of MUX21_L_292 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_291 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_291;

architecture SYN_BEHAVIORAL of MUX21_L_291 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_290 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_290;

architecture SYN_BEHAVIORAL of MUX21_L_290 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_289 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_289;

architecture SYN_BEHAVIORAL of MUX21_L_289 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_288 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_288;

architecture SYN_BEHAVIORAL of MUX21_L_288 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_287 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_287;

architecture SYN_BEHAVIORAL of MUX21_L_287 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_286 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_286;

architecture SYN_BEHAVIORAL of MUX21_L_286 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_285 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_285;

architecture SYN_BEHAVIORAL of MUX21_L_285 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_284 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_284;

architecture SYN_BEHAVIORAL of MUX21_L_284 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_283 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_283;

architecture SYN_BEHAVIORAL of MUX21_L_283 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_282 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_282;

architecture SYN_BEHAVIORAL of MUX21_L_282 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_281 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_281;

architecture SYN_BEHAVIORAL of MUX21_L_281 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_280 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_280;

architecture SYN_BEHAVIORAL of MUX21_L_280 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_279 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_279;

architecture SYN_BEHAVIORAL of MUX21_L_279 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_278 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_278;

architecture SYN_BEHAVIORAL of MUX21_L_278 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_277 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_277;

architecture SYN_BEHAVIORAL of MUX21_L_277 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_276 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_276;

architecture SYN_BEHAVIORAL of MUX21_L_276 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_275 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_275;

architecture SYN_BEHAVIORAL of MUX21_L_275 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_274 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_274;

architecture SYN_BEHAVIORAL of MUX21_L_274 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_273 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_273;

architecture SYN_BEHAVIORAL of MUX21_L_273 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_272 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_272;

architecture SYN_BEHAVIORAL of MUX21_L_272 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_271 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_271;

architecture SYN_BEHAVIORAL of MUX21_L_271 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_270 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_270;

architecture SYN_BEHAVIORAL of MUX21_L_270 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_269 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_269;

architecture SYN_BEHAVIORAL of MUX21_L_269 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_268 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_268;

architecture SYN_BEHAVIORAL of MUX21_L_268 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_267 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_267;

architecture SYN_BEHAVIORAL of MUX21_L_267 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_266 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_266;

architecture SYN_BEHAVIORAL of MUX21_L_266 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_265 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_265;

architecture SYN_BEHAVIORAL of MUX21_L_265 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_264 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_264;

architecture SYN_BEHAVIORAL of MUX21_L_264 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_263 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_263;

architecture SYN_BEHAVIORAL of MUX21_L_263 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_262 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_262;

architecture SYN_BEHAVIORAL of MUX21_L_262 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_261 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_261;

architecture SYN_BEHAVIORAL of MUX21_L_261 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_260 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_260;

architecture SYN_BEHAVIORAL of MUX21_L_260 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_259 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_259;

architecture SYN_BEHAVIORAL of MUX21_L_259 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_258 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_258;

architecture SYN_BEHAVIORAL of MUX21_L_258 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_257 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_257;

architecture SYN_BEHAVIORAL of MUX21_L_257 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_256 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_256;

architecture SYN_BEHAVIORAL of MUX21_L_256 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_255 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_255;

architecture SYN_BEHAVIORAL of MUX21_L_255 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_254 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_254;

architecture SYN_BEHAVIORAL of MUX21_L_254 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_253 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_253;

architecture SYN_BEHAVIORAL of MUX21_L_253 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_252 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_252;

architecture SYN_BEHAVIORAL of MUX21_L_252 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_251 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_251;

architecture SYN_BEHAVIORAL of MUX21_L_251 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_250 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_250;

architecture SYN_BEHAVIORAL of MUX21_L_250 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_249 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_249;

architecture SYN_BEHAVIORAL of MUX21_L_249 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_248 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_248;

architecture SYN_BEHAVIORAL of MUX21_L_248 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_247 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_247;

architecture SYN_BEHAVIORAL of MUX21_L_247 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_246 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_246;

architecture SYN_BEHAVIORAL of MUX21_L_246 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_245 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_245;

architecture SYN_BEHAVIORAL of MUX21_L_245 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_244 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_244;

architecture SYN_BEHAVIORAL of MUX21_L_244 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_243 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_243;

architecture SYN_BEHAVIORAL of MUX21_L_243 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_242 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_242;

architecture SYN_BEHAVIORAL of MUX21_L_242 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_241 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_241;

architecture SYN_BEHAVIORAL of MUX21_L_241 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_240 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_240;

architecture SYN_BEHAVIORAL of MUX21_L_240 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_239 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_239;

architecture SYN_BEHAVIORAL of MUX21_L_239 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_238 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_238;

architecture SYN_BEHAVIORAL of MUX21_L_238 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_237 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_237;

architecture SYN_BEHAVIORAL of MUX21_L_237 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_236 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_236;

architecture SYN_BEHAVIORAL of MUX21_L_236 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_235 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_235;

architecture SYN_BEHAVIORAL of MUX21_L_235 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_234 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_234;

architecture SYN_BEHAVIORAL of MUX21_L_234 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_233 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_233;

architecture SYN_BEHAVIORAL of MUX21_L_233 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_232 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_232;

architecture SYN_BEHAVIORAL of MUX21_L_232 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_231 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_231;

architecture SYN_BEHAVIORAL of MUX21_L_231 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_230 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_230;

architecture SYN_BEHAVIORAL of MUX21_L_230 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_229 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_229;

architecture SYN_BEHAVIORAL of MUX21_L_229 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_228 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_228;

architecture SYN_BEHAVIORAL of MUX21_L_228 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_227 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_227;

architecture SYN_BEHAVIORAL of MUX21_L_227 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_226 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_226;

architecture SYN_BEHAVIORAL of MUX21_L_226 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_225 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_225;

architecture SYN_BEHAVIORAL of MUX21_L_225 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_224 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_224;

architecture SYN_BEHAVIORAL of MUX21_L_224 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_223 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_223;

architecture SYN_BEHAVIORAL of MUX21_L_223 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_222 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_222;

architecture SYN_BEHAVIORAL of MUX21_L_222 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_221 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_221;

architecture SYN_BEHAVIORAL of MUX21_L_221 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_220 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_220;

architecture SYN_BEHAVIORAL of MUX21_L_220 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_219 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_219;

architecture SYN_BEHAVIORAL of MUX21_L_219 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_218 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_218;

architecture SYN_BEHAVIORAL of MUX21_L_218 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_217 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_217;

architecture SYN_BEHAVIORAL of MUX21_L_217 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_216 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_216;

architecture SYN_BEHAVIORAL of MUX21_L_216 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_215 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_215;

architecture SYN_BEHAVIORAL of MUX21_L_215 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_214 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_214;

architecture SYN_BEHAVIORAL of MUX21_L_214 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_213 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_213;

architecture SYN_BEHAVIORAL of MUX21_L_213 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_212 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_212;

architecture SYN_BEHAVIORAL of MUX21_L_212 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_211 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_211;

architecture SYN_BEHAVIORAL of MUX21_L_211 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_210 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_210;

architecture SYN_BEHAVIORAL of MUX21_L_210 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_209 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_209;

architecture SYN_BEHAVIORAL of MUX21_L_209 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_208 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_208;

architecture SYN_BEHAVIORAL of MUX21_L_208 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_207 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_207;

architecture SYN_BEHAVIORAL of MUX21_L_207 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_206 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_206;

architecture SYN_BEHAVIORAL of MUX21_L_206 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_205 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_205;

architecture SYN_BEHAVIORAL of MUX21_L_205 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_204 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_204;

architecture SYN_BEHAVIORAL of MUX21_L_204 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_203 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_203;

architecture SYN_BEHAVIORAL of MUX21_L_203 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_202 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_202;

architecture SYN_BEHAVIORAL of MUX21_L_202 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_201 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_201;

architecture SYN_BEHAVIORAL of MUX21_L_201 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_200 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_200;

architecture SYN_BEHAVIORAL of MUX21_L_200 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_199 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_199;

architecture SYN_BEHAVIORAL of MUX21_L_199 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_198 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_198;

architecture SYN_BEHAVIORAL of MUX21_L_198 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_197 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_197;

architecture SYN_BEHAVIORAL of MUX21_L_197 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_196 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_196;

architecture SYN_BEHAVIORAL of MUX21_L_196 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_195 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_195;

architecture SYN_BEHAVIORAL of MUX21_L_195 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_194 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_194;

architecture SYN_BEHAVIORAL of MUX21_L_194 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_193 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_193;

architecture SYN_BEHAVIORAL of MUX21_L_193 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_192 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_192;

architecture SYN_BEHAVIORAL of MUX21_L_192 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_191 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_191;

architecture SYN_BEHAVIORAL of MUX21_L_191 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_190 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_190;

architecture SYN_BEHAVIORAL of MUX21_L_190 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_189 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_189;

architecture SYN_BEHAVIORAL of MUX21_L_189 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_188 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_188;

architecture SYN_BEHAVIORAL of MUX21_L_188 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_187 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_187;

architecture SYN_BEHAVIORAL of MUX21_L_187 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_186 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_186;

architecture SYN_BEHAVIORAL of MUX21_L_186 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_185 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_185;

architecture SYN_BEHAVIORAL of MUX21_L_185 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_184 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_184;

architecture SYN_BEHAVIORAL of MUX21_L_184 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_183 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_183;

architecture SYN_BEHAVIORAL of MUX21_L_183 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_182 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_182;

architecture SYN_BEHAVIORAL of MUX21_L_182 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_181 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_181;

architecture SYN_BEHAVIORAL of MUX21_L_181 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_180 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_180;

architecture SYN_BEHAVIORAL of MUX21_L_180 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_179 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_179;

architecture SYN_BEHAVIORAL of MUX21_L_179 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_178 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_178;

architecture SYN_BEHAVIORAL of MUX21_L_178 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_177 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_177;

architecture SYN_BEHAVIORAL of MUX21_L_177 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_176 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_176;

architecture SYN_BEHAVIORAL of MUX21_L_176 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_175 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_175;

architecture SYN_BEHAVIORAL of MUX21_L_175 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_174 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_174;

architecture SYN_BEHAVIORAL of MUX21_L_174 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_173 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_173;

architecture SYN_BEHAVIORAL of MUX21_L_173 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_172 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_172;

architecture SYN_BEHAVIORAL of MUX21_L_172 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_171 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_171;

architecture SYN_BEHAVIORAL of MUX21_L_171 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_170 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_170;

architecture SYN_BEHAVIORAL of MUX21_L_170 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_169 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_169;

architecture SYN_BEHAVIORAL of MUX21_L_169 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_168 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_168;

architecture SYN_BEHAVIORAL of MUX21_L_168 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_167 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_167;

architecture SYN_BEHAVIORAL of MUX21_L_167 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_166 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_166;

architecture SYN_BEHAVIORAL of MUX21_L_166 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_165 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_165;

architecture SYN_BEHAVIORAL of MUX21_L_165 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_164 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_164;

architecture SYN_BEHAVIORAL of MUX21_L_164 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_163 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_163;

architecture SYN_BEHAVIORAL of MUX21_L_163 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_162 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_162;

architecture SYN_BEHAVIORAL of MUX21_L_162 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_161 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_161;

architecture SYN_BEHAVIORAL of MUX21_L_161 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_160 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_160;

architecture SYN_BEHAVIORAL of MUX21_L_160 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_159 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_159;

architecture SYN_BEHAVIORAL of MUX21_L_159 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_158 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_158;

architecture SYN_BEHAVIORAL of MUX21_L_158 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_157 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_157;

architecture SYN_BEHAVIORAL of MUX21_L_157 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_156 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_156;

architecture SYN_BEHAVIORAL of MUX21_L_156 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_155 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_155;

architecture SYN_BEHAVIORAL of MUX21_L_155 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_154 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_154;

architecture SYN_BEHAVIORAL of MUX21_L_154 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_153 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_153;

architecture SYN_BEHAVIORAL of MUX21_L_153 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_152 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_152;

architecture SYN_BEHAVIORAL of MUX21_L_152 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_151 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_151;

architecture SYN_BEHAVIORAL of MUX21_L_151 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_150 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_150;

architecture SYN_BEHAVIORAL of MUX21_L_150 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_149 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_149;

architecture SYN_BEHAVIORAL of MUX21_L_149 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_148 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_148;

architecture SYN_BEHAVIORAL of MUX21_L_148 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_147 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_147;

architecture SYN_BEHAVIORAL of MUX21_L_147 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_146 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_146;

architecture SYN_BEHAVIORAL of MUX21_L_146 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_145 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_145;

architecture SYN_BEHAVIORAL of MUX21_L_145 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_144 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_144;

architecture SYN_BEHAVIORAL of MUX21_L_144 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_143 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_143;

architecture SYN_BEHAVIORAL of MUX21_L_143 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_142 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_142;

architecture SYN_BEHAVIORAL of MUX21_L_142 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_141 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_141;

architecture SYN_BEHAVIORAL of MUX21_L_141 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_140 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_140;

architecture SYN_BEHAVIORAL of MUX21_L_140 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_139 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_139;

architecture SYN_BEHAVIORAL of MUX21_L_139 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_138 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_138;

architecture SYN_BEHAVIORAL of MUX21_L_138 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_137 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_137;

architecture SYN_BEHAVIORAL of MUX21_L_137 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_136 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_136;

architecture SYN_BEHAVIORAL of MUX21_L_136 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_135 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_135;

architecture SYN_BEHAVIORAL of MUX21_L_135 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_134 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_134;

architecture SYN_BEHAVIORAL of MUX21_L_134 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_133 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_133;

architecture SYN_BEHAVIORAL of MUX21_L_133 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_132 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_132;

architecture SYN_BEHAVIORAL of MUX21_L_132 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_131 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_131;

architecture SYN_BEHAVIORAL of MUX21_L_131 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_130 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_130;

architecture SYN_BEHAVIORAL of MUX21_L_130 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_129 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_129;

architecture SYN_BEHAVIORAL of MUX21_L_129 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_128 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_128;

architecture SYN_BEHAVIORAL of MUX21_L_128 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_127 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_127;

architecture SYN_BEHAVIORAL of MUX21_L_127 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_126 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_126;

architecture SYN_BEHAVIORAL of MUX21_L_126 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_125 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_125;

architecture SYN_BEHAVIORAL of MUX21_L_125 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_124 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_124;

architecture SYN_BEHAVIORAL of MUX21_L_124 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_123 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_123;

architecture SYN_BEHAVIORAL of MUX21_L_123 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_122 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_122;

architecture SYN_BEHAVIORAL of MUX21_L_122 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_121 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_121;

architecture SYN_BEHAVIORAL of MUX21_L_121 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_120 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_120;

architecture SYN_BEHAVIORAL of MUX21_L_120 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_119 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_119;

architecture SYN_BEHAVIORAL of MUX21_L_119 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_118 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_118;

architecture SYN_BEHAVIORAL of MUX21_L_118 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_117 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_117;

architecture SYN_BEHAVIORAL of MUX21_L_117 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_116 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_116;

architecture SYN_BEHAVIORAL of MUX21_L_116 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_115 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_115;

architecture SYN_BEHAVIORAL of MUX21_L_115 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_114 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_114;

architecture SYN_BEHAVIORAL of MUX21_L_114 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_113 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_113;

architecture SYN_BEHAVIORAL of MUX21_L_113 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_112 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_112;

architecture SYN_BEHAVIORAL of MUX21_L_112 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_111 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_111;

architecture SYN_BEHAVIORAL of MUX21_L_111 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_110 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_110;

architecture SYN_BEHAVIORAL of MUX21_L_110 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_109 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_109;

architecture SYN_BEHAVIORAL of MUX21_L_109 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_108 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_108;

architecture SYN_BEHAVIORAL of MUX21_L_108 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_107 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_107;

architecture SYN_BEHAVIORAL of MUX21_L_107 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_106 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_106;

architecture SYN_BEHAVIORAL of MUX21_L_106 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_105 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_105;

architecture SYN_BEHAVIORAL of MUX21_L_105 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_104 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_104;

architecture SYN_BEHAVIORAL of MUX21_L_104 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_103 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_103;

architecture SYN_BEHAVIORAL of MUX21_L_103 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_102 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_102;

architecture SYN_BEHAVIORAL of MUX21_L_102 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_101 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_101;

architecture SYN_BEHAVIORAL of MUX21_L_101 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_100 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_100;

architecture SYN_BEHAVIORAL of MUX21_L_100 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_99 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_99;

architecture SYN_BEHAVIORAL of MUX21_L_99 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_98 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_98;

architecture SYN_BEHAVIORAL of MUX21_L_98 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_97 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_97;

architecture SYN_BEHAVIORAL of MUX21_L_97 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_96 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_96;

architecture SYN_BEHAVIORAL of MUX21_L_96 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_95 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_95;

architecture SYN_BEHAVIORAL of MUX21_L_95 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_94 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_94;

architecture SYN_BEHAVIORAL of MUX21_L_94 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_93 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_93;

architecture SYN_BEHAVIORAL of MUX21_L_93 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_92 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_92;

architecture SYN_BEHAVIORAL of MUX21_L_92 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_91 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_91;

architecture SYN_BEHAVIORAL of MUX21_L_91 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_90 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_90;

architecture SYN_BEHAVIORAL of MUX21_L_90 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_89 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_89;

architecture SYN_BEHAVIORAL of MUX21_L_89 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_88 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_88;

architecture SYN_BEHAVIORAL of MUX21_L_88 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_87 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_87;

architecture SYN_BEHAVIORAL of MUX21_L_87 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_86 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_86;

architecture SYN_BEHAVIORAL of MUX21_L_86 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_85 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_85;

architecture SYN_BEHAVIORAL of MUX21_L_85 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_84 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_84;

architecture SYN_BEHAVIORAL of MUX21_L_84 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_83 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_83;

architecture SYN_BEHAVIORAL of MUX21_L_83 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_82 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_82;

architecture SYN_BEHAVIORAL of MUX21_L_82 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_81 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_81;

architecture SYN_BEHAVIORAL of MUX21_L_81 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_80 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_80;

architecture SYN_BEHAVIORAL of MUX21_L_80 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_79 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_79;

architecture SYN_BEHAVIORAL of MUX21_L_79 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_78 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_78;

architecture SYN_BEHAVIORAL of MUX21_L_78 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_77 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_77;

architecture SYN_BEHAVIORAL of MUX21_L_77 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_76 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_76;

architecture SYN_BEHAVIORAL of MUX21_L_76 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_75 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_75;

architecture SYN_BEHAVIORAL of MUX21_L_75 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_74 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_74;

architecture SYN_BEHAVIORAL of MUX21_L_74 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_73 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_73;

architecture SYN_BEHAVIORAL of MUX21_L_73 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_72 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_72;

architecture SYN_BEHAVIORAL of MUX21_L_72 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_71 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_71;

architecture SYN_BEHAVIORAL of MUX21_L_71 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_70 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_70;

architecture SYN_BEHAVIORAL of MUX21_L_70 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_69 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_69;

architecture SYN_BEHAVIORAL of MUX21_L_69 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_68 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_68;

architecture SYN_BEHAVIORAL of MUX21_L_68 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_67 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_67;

architecture SYN_BEHAVIORAL of MUX21_L_67 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_66 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_66;

architecture SYN_BEHAVIORAL of MUX21_L_66 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_65 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_65;

architecture SYN_BEHAVIORAL of MUX21_L_65 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_64 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_64;

architecture SYN_BEHAVIORAL of MUX21_L_64 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_63 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_63;

architecture SYN_BEHAVIORAL of MUX21_L_63 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_62 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_62;

architecture SYN_BEHAVIORAL of MUX21_L_62 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_61 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_61;

architecture SYN_BEHAVIORAL of MUX21_L_61 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_60 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_60;

architecture SYN_BEHAVIORAL of MUX21_L_60 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_59 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_59;

architecture SYN_BEHAVIORAL of MUX21_L_59 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_58 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_58;

architecture SYN_BEHAVIORAL of MUX21_L_58 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_57 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_57;

architecture SYN_BEHAVIORAL of MUX21_L_57 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_56 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_56;

architecture SYN_BEHAVIORAL of MUX21_L_56 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_55 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_55;

architecture SYN_BEHAVIORAL of MUX21_L_55 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_54 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_54;

architecture SYN_BEHAVIORAL of MUX21_L_54 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_53 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_53;

architecture SYN_BEHAVIORAL of MUX21_L_53 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_52 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_52;

architecture SYN_BEHAVIORAL of MUX21_L_52 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_51 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_51;

architecture SYN_BEHAVIORAL of MUX21_L_51 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_50 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_50;

architecture SYN_BEHAVIORAL of MUX21_L_50 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_49 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_49;

architecture SYN_BEHAVIORAL of MUX21_L_49 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_48 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_48;

architecture SYN_BEHAVIORAL of MUX21_L_48 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_47 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_47;

architecture SYN_BEHAVIORAL of MUX21_L_47 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_46 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_46;

architecture SYN_BEHAVIORAL of MUX21_L_46 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_45 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_45;

architecture SYN_BEHAVIORAL of MUX21_L_45 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_44 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_44;

architecture SYN_BEHAVIORAL of MUX21_L_44 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_43 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_43;

architecture SYN_BEHAVIORAL of MUX21_L_43 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_42 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_42;

architecture SYN_BEHAVIORAL of MUX21_L_42 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_41 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_41;

architecture SYN_BEHAVIORAL of MUX21_L_41 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_40 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_40;

architecture SYN_BEHAVIORAL of MUX21_L_40 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_39 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_39;

architecture SYN_BEHAVIORAL of MUX21_L_39 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_38 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_38;

architecture SYN_BEHAVIORAL of MUX21_L_38 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_37 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_37;

architecture SYN_BEHAVIORAL of MUX21_L_37 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_36 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_36;

architecture SYN_BEHAVIORAL of MUX21_L_36 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_35 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_35;

architecture SYN_BEHAVIORAL of MUX21_L_35 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_34 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_34;

architecture SYN_BEHAVIORAL of MUX21_L_34 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_33 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_33;

architecture SYN_BEHAVIORAL of MUX21_L_33 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_32 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_32;

architecture SYN_BEHAVIORAL of MUX21_L_32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_31;

architecture SYN_BEHAVIORAL of MUX21_L_31 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_30;

architecture SYN_BEHAVIORAL of MUX21_L_30 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_29;

architecture SYN_BEHAVIORAL of MUX21_L_29 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_28;

architecture SYN_BEHAVIORAL of MUX21_L_28 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_27;

architecture SYN_BEHAVIORAL of MUX21_L_27 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_26;

architecture SYN_BEHAVIORAL of MUX21_L_26 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_25;

architecture SYN_BEHAVIORAL of MUX21_L_25 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_24;

architecture SYN_BEHAVIORAL of MUX21_L_24 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_23;

architecture SYN_BEHAVIORAL of MUX21_L_23 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_22;

architecture SYN_BEHAVIORAL of MUX21_L_22 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_21;

architecture SYN_BEHAVIORAL of MUX21_L_21 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_20;

architecture SYN_BEHAVIORAL of MUX21_L_20 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_19;

architecture SYN_BEHAVIORAL of MUX21_L_19 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_18;

architecture SYN_BEHAVIORAL of MUX21_L_18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_17;

architecture SYN_BEHAVIORAL of MUX21_L_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_16;

architecture SYN_BEHAVIORAL of MUX21_L_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_15;

architecture SYN_BEHAVIORAL of MUX21_L_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_14;

architecture SYN_BEHAVIORAL of MUX21_L_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_13;

architecture SYN_BEHAVIORAL of MUX21_L_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_12;

architecture SYN_BEHAVIORAL of MUX21_L_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_11;

architecture SYN_BEHAVIORAL of MUX21_L_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_10;

architecture SYN_BEHAVIORAL of MUX21_L_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_9;

architecture SYN_BEHAVIORAL of MUX21_L_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_8;

architecture SYN_BEHAVIORAL of MUX21_L_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_7;

architecture SYN_BEHAVIORAL of MUX21_L_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_6;

architecture SYN_BEHAVIORAL of MUX21_L_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_5;

architecture SYN_BEHAVIORAL of MUX21_L_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_4;

architecture SYN_BEHAVIORAL of MUX21_L_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_3;

architecture SYN_BEHAVIORAL of MUX21_L_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_2;

architecture SYN_BEHAVIORAL of MUX21_L_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_1;

architecture SYN_BEHAVIORAL of MUX21_L_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_0;

architecture SYN_BEHAVIORAL of MUX21_L_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end MUX21_N4_7;

architecture SYN_BEHAVIORAL of MUX21_N4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_BEHAVIORAL of RCA_N4_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(3));
   U2 : XNOR2_X1 port map( A => A(3), B => B(3), ZN => n2);
   U3 : XOR2_X1 port map( A => n3, B => n4, Z => S(2));
   U4 : XOR2_X1 port map( A => B(2), B => A(2), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => n6, ZN => S(1));
   U6 : XNOR2_X1 port map( A => B(1), B => n7, ZN => n6);
   U7 : XOR2_X1 port map( A => A(0), B => n8, Z => S(0));
   U8 : XOR2_X1 port map( A => Ci, B => B(0), Z => n8);
   U9 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11, ZN => Co);
   U10 : OAI21_X1 port map( B1 => n1, B2 => A(3), A => B(3), ZN => n11);
   U11 : INV_X1 port map( A => n10, ZN => n1);
   U12 : OAI21_X1 port map( B1 => A(2), B2 => n3, A => n12, ZN => n10);
   U13 : INV_X1 port map( A => n13, ZN => n12);
   U14 : AOI21_X1 port map( B1 => n3, B2 => A(2), A => B(2), ZN => n13);
   U15 : AOI21_X1 port map( B1 => n7, B2 => n5, A => n14, ZN => n3);
   U16 : AOI21_X1 port map( B1 => n15, B2 => A(1), A => B(1), ZN => n14);
   U17 : INV_X1 port map( A => n5, ZN => n15);
   U18 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => n16, ZN => n5);
   U19 : INV_X1 port map( A => n17, ZN => n16);
   U20 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n17);
   U21 : INV_X1 port map( A => A(1), ZN => n7);
   U22 : INV_X1 port map( A => A(3), ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ENCODER_7 is

   port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end ENCODER_7;

architecture SYN_BEHAVIORAL of ENCODER_7 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : AND3_X1 port map( A1 => B(2), A2 => n1, A3 => n2, ZN => Y(2));
   U4 : INV_X1 port map( A => n3, ZN => Y(1));
   U5 : MUX2_X1 port map( A => n1, B => n2, S => B(2), Z => n3);
   U6 : AOI21_X1 port map( B1 => n2, B2 => n1, A => B(2), ZN => Y(0));
   U7 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n1);
   U8 : XNOR2_X1 port map( A => B(0), B => B(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_6;

architecture SYN_STRUCTURAL of CSB_N4_6 is

   component MUX21_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1251, 
      n_1252 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1251);
   RCA1 : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1252);
   MUX : MUX21_N4_6 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CSB_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_N4_7;

architecture SYN_STRUCTURAL of CSB_N4_7 is

   component MUX21_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, SUM0_3_port, SUM0_2_port, SUM0_1_port, 
      SUM0_0_port, SUM1_3_port, SUM1_2_port, SUM1_1_port, SUM1_0_port, n_1253, 
      n_1254 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => SUM0_3_port, 
                           S(2) => SUM0_2_port, S(1) => SUM0_1_port, S(0) => 
                           SUM0_0_port, Co => n_1253);
   RCA1 : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => SUM1_3_port, 
                           S(2) => SUM1_2_port, S(1) => SUM1_1_port, S(0) => 
                           SUM1_0_port, Co => n_1254);
   MUX : MUX21_N4_7 port map( A(3) => SUM0_3_port, A(2) => SUM0_2_port, A(1) =>
                           SUM0_1_port, A(0) => SUM0_0_port, B(3) => 
                           SUM1_3_port, B(2) => SUM1_2_port, B(1) => 
                           SUM1_1_port, B(0) => SUM1_0_port, S => Ci, Y(3) => 
                           S(3), Y(2) => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_BLOCK_33 is

   port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);

end PG_BLOCK_33;

architecture SYN_BEHAVIORAL of PG_BLOCK_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pkj, A2 => Pik, ZN => Pij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity GENERATE_BLOCK_8 is

   port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);

end GENERATE_BLOCK_8;

architecture SYN_BEHAVIORAL of GENERATE_BLOCK_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gkj, A => Gik, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_ROW_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  P, G : 
         out std_logic_vector (31 downto 0));

end PG_ROW_N32;

architecture SYN_BEHAVIORAL of PG_ROW_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B(9), B => A(9), Z => P(9));
   U2 : XOR2_X1 port map( A => B(8), B => A(8), Z => P(8));
   U3 : XOR2_X1 port map( A => B(7), B => A(7), Z => P(7));
   U4 : XOR2_X1 port map( A => B(6), B => A(6), Z => P(6));
   U5 : XOR2_X1 port map( A => B(5), B => A(5), Z => P(5));
   U6 : XOR2_X1 port map( A => B(4), B => A(4), Z => P(4));
   U7 : XOR2_X1 port map( A => B(3), B => A(3), Z => P(3));
   U8 : XOR2_X1 port map( A => B(31), B => A(31), Z => P(31));
   U9 : XOR2_X1 port map( A => B(30), B => A(30), Z => P(30));
   U10 : XOR2_X1 port map( A => B(2), B => A(2), Z => P(2));
   U11 : XOR2_X1 port map( A => B(29), B => A(29), Z => P(29));
   U12 : XOR2_X1 port map( A => B(28), B => A(28), Z => P(28));
   U13 : XOR2_X1 port map( A => B(27), B => A(27), Z => P(27));
   U14 : XOR2_X1 port map( A => B(26), B => A(26), Z => P(26));
   U15 : XOR2_X1 port map( A => B(25), B => A(25), Z => P(25));
   U16 : XOR2_X1 port map( A => B(24), B => A(24), Z => P(24));
   U17 : XOR2_X1 port map( A => B(23), B => A(23), Z => P(23));
   U18 : XOR2_X1 port map( A => B(22), B => A(22), Z => P(22));
   U19 : XOR2_X1 port map( A => B(21), B => A(21), Z => P(21));
   U20 : XOR2_X1 port map( A => B(20), B => A(20), Z => P(20));
   U21 : XOR2_X1 port map( A => B(1), B => A(1), Z => P(1));
   U22 : XOR2_X1 port map( A => B(19), B => A(19), Z => P(19));
   U23 : XOR2_X1 port map( A => B(18), B => A(18), Z => P(18));
   U24 : XOR2_X1 port map( A => B(17), B => A(17), Z => P(17));
   U25 : XOR2_X1 port map( A => B(16), B => A(16), Z => P(16));
   U26 : XOR2_X1 port map( A => B(15), B => A(15), Z => P(15));
   U27 : XOR2_X1 port map( A => B(14), B => A(14), Z => P(14));
   U28 : XOR2_X1 port map( A => B(13), B => A(13), Z => P(13));
   U29 : XOR2_X1 port map( A => B(12), B => A(12), Z => P(12));
   U30 : XOR2_X1 port map( A => B(11), B => A(11), Z => P(11));
   U31 : XOR2_X1 port map( A => B(10), B => A(10), Z => P(10));
   U32 : XNOR2_X1 port map( A => n1, B => A(0), ZN => P(0));
   U33 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => G(9));
   U34 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => G(8));
   U35 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => G(7));
   U36 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => G(6));
   U37 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => G(5));
   U38 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => G(4));
   U39 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => G(3));
   U40 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => G(31));
   U41 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => G(30));
   U42 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => G(2));
   U43 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => G(29));
   U44 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => G(28));
   U45 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => G(27));
   U46 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => G(26));
   U47 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => G(25));
   U48 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => G(24));
   U49 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => G(23));
   U50 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => G(22));
   U51 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => G(21));
   U52 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => G(20));
   U53 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => G(1));
   U54 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => G(19));
   U55 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => G(18));
   U56 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => G(17));
   U57 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => G(16));
   U58 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => G(15));
   U59 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => G(14));
   U60 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => G(13));
   U61 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => G(12));
   U62 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => G(11));
   U63 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => G(10));
   U64 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => G(0));
   U65 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n3);
   U66 : INV_X1 port map( A => A(0), ZN => n2);
   U67 : INV_X1 port map( A => B(0), ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_N32_2;

architecture SYN_BEHAVIORAL of RCA_N32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n2, ZN => S(9));
   U2 : XOR2_X1 port map( A => B(9), B => A(9), Z => n2);
   U3 : XNOR2_X1 port map( A => n3, B => n4, ZN => S(8));
   U4 : XNOR2_X1 port map( A => A(8), B => B(8), ZN => n4);
   U5 : XOR2_X1 port map( A => n5, B => n6, Z => S(7));
   U6 : XNOR2_X1 port map( A => B(7), B => n7, ZN => n6);
   U7 : XNOR2_X1 port map( A => n8, B => n9, ZN => S(6));
   U8 : XNOR2_X1 port map( A => A(6), B => B(6), ZN => n9);
   U9 : XOR2_X1 port map( A => n10, B => n11, Z => S(5));
   U10 : XOR2_X1 port map( A => B(5), B => A(5), Z => n11);
   U11 : XNOR2_X1 port map( A => n12, B => n13, ZN => S(4));
   U12 : XNOR2_X1 port map( A => A(4), B => B(4), ZN => n13);
   U13 : XNOR2_X1 port map( A => n14, B => n15, ZN => S(3));
   U14 : XNOR2_X1 port map( A => B(3), B => n16, ZN => n15);
   U15 : XOR2_X1 port map( A => n17, B => n18, Z => S(31));
   U16 : XOR2_X1 port map( A => B(31), B => A(31), Z => n18);
   U17 : XNOR2_X1 port map( A => n19, B => n20, ZN => S(30));
   U18 : XNOR2_X1 port map( A => B(30), B => n21, ZN => n20);
   U19 : XNOR2_X1 port map( A => n22, B => n23, ZN => S(2));
   U20 : XOR2_X1 port map( A => B(2), B => A(2), Z => n23);
   U21 : XOR2_X1 port map( A => n24, B => n25, Z => S(29));
   U22 : XOR2_X1 port map( A => B(29), B => A(29), Z => n25);
   U23 : XNOR2_X1 port map( A => n26, B => n27, ZN => S(28));
   U24 : XNOR2_X1 port map( A => B(28), B => n28, ZN => n27);
   U25 : XNOR2_X1 port map( A => n29, B => n30, ZN => S(27));
   U26 : XOR2_X1 port map( A => B(27), B => A(27), Z => n30);
   U27 : XOR2_X1 port map( A => n31, B => n32, Z => S(26));
   U28 : XOR2_X1 port map( A => B(26), B => A(26), Z => n32);
   U29 : XNOR2_X1 port map( A => n33, B => n34, ZN => S(25));
   U30 : XNOR2_X1 port map( A => B(25), B => n35, ZN => n34);
   U31 : XOR2_X1 port map( A => n36, B => n37, Z => S(24));
   U32 : XOR2_X1 port map( A => B(24), B => A(24), Z => n37);
   U33 : XNOR2_X1 port map( A => n38, B => n39, ZN => S(23));
   U34 : XNOR2_X1 port map( A => B(23), B => n40, ZN => n39);
   U35 : XOR2_X1 port map( A => n41, B => n42, Z => S(22));
   U36 : XOR2_X1 port map( A => B(22), B => A(22), Z => n42);
   U37 : XNOR2_X1 port map( A => n43, B => n44, ZN => S(21));
   U38 : XNOR2_X1 port map( A => B(21), B => n45, ZN => n44);
   U39 : XOR2_X1 port map( A => n46, B => n47, Z => S(20));
   U40 : XOR2_X1 port map( A => B(20), B => A(20), Z => n47);
   U41 : XNOR2_X1 port map( A => n48, B => n49, ZN => S(1));
   U42 : XOR2_X1 port map( A => B(1), B => A(1), Z => n49);
   U43 : XNOR2_X1 port map( A => n50, B => n51, ZN => S(19));
   U44 : XNOR2_X1 port map( A => B(19), B => n52, ZN => n51);
   U45 : XNOR2_X1 port map( A => n53, B => n54, ZN => S(18));
   U46 : XNOR2_X1 port map( A => B(18), B => n55, ZN => n54);
   U47 : XOR2_X1 port map( A => n56, B => n57, Z => S(17));
   U48 : XOR2_X1 port map( A => B(17), B => A(17), Z => n57);
   U49 : XNOR2_X1 port map( A => n58, B => n59, ZN => S(16));
   U50 : XNOR2_X1 port map( A => B(16), B => n60, ZN => n59);
   U51 : XOR2_X1 port map( A => n61, B => n62, Z => S(15));
   U52 : XOR2_X1 port map( A => B(15), B => A(15), Z => n62);
   U53 : XNOR2_X1 port map( A => n63, B => n64, ZN => S(14));
   U54 : XOR2_X1 port map( A => B(14), B => A(14), Z => n64);
   U55 : XOR2_X1 port map( A => n65, B => n66, Z => S(13));
   U56 : XOR2_X1 port map( A => B(13), B => A(13), Z => n66);
   U57 : XNOR2_X1 port map( A => n67, B => n68, ZN => S(12));
   U58 : XNOR2_X1 port map( A => A(12), B => B(12), ZN => n68);
   U59 : XOR2_X1 port map( A => n69, B => n70, Z => S(11));
   U60 : XOR2_X1 port map( A => B(11), B => A(11), Z => n70);
   U61 : XNOR2_X1 port map( A => n71, B => n72, ZN => S(10));
   U62 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => n72);
   U63 : XOR2_X1 port map( A => A(0), B => n73, Z => S(0));
   U64 : XOR2_X1 port map( A => Ci, B => B(0), Z => n73);
   U65 : INV_X1 port map( A => n74, ZN => Co);
   U66 : AOI22_X1 port map( A1 => A(31), A2 => n17, B1 => n75, B2 => B(31), ZN 
                           => n74);
   U67 : OR2_X1 port map( A1 => n17, A2 => A(31), ZN => n75);
   U68 : AOI21_X1 port map( B1 => n21, B2 => n19, A => n76, ZN => n17);
   U69 : AOI21_X1 port map( B1 => n77, B2 => A(30), A => B(30), ZN => n76);
   U70 : INV_X1 port map( A => n19, ZN => n77);
   U71 : AOI22_X1 port map( A1 => n24, A2 => A(29), B1 => n78, B2 => B(29), ZN 
                           => n19);
   U72 : OR2_X1 port map( A1 => A(29), A2 => n24, ZN => n78);
   U73 : OAI21_X1 port map( B1 => n26, B2 => n28, A => n79, ZN => n24);
   U74 : OAI21_X1 port map( B1 => n80, B2 => A(28), A => B(28), ZN => n79);
   U75 : INV_X1 port map( A => n26, ZN => n80);
   U76 : INV_X1 port map( A => A(28), ZN => n28);
   U77 : OAI21_X1 port map( B1 => A(27), B2 => n81, A => n82, ZN => n26);
   U78 : INV_X1 port map( A => n83, ZN => n82);
   U79 : AOI21_X1 port map( B1 => n81, B2 => A(27), A => B(27), ZN => n83);
   U80 : INV_X1 port map( A => n29, ZN => n81);
   U81 : AOI22_X1 port map( A1 => n31, A2 => A(26), B1 => n84, B2 => B(26), ZN 
                           => n29);
   U82 : OR2_X1 port map( A1 => n31, A2 => A(26), ZN => n84);
   U83 : AOI21_X1 port map( B1 => n35, B2 => n33, A => n85, ZN => n31);
   U84 : AOI21_X1 port map( B1 => n86, B2 => A(25), A => B(25), ZN => n85);
   U85 : INV_X1 port map( A => n33, ZN => n86);
   U86 : AOI21_X1 port map( B1 => n36, B2 => A(24), A => n87, ZN => n33);
   U87 : INV_X1 port map( A => n88, ZN => n87);
   U88 : OAI21_X1 port map( B1 => n36, B2 => A(24), A => B(24), ZN => n88);
   U89 : AOI21_X1 port map( B1 => n40, B2 => n38, A => n89, ZN => n36);
   U90 : AOI21_X1 port map( B1 => n90, B2 => A(23), A => B(23), ZN => n89);
   U91 : INV_X1 port map( A => n38, ZN => n90);
   U92 : AOI21_X1 port map( B1 => n41, B2 => A(22), A => n91, ZN => n38);
   U93 : INV_X1 port map( A => n92, ZN => n91);
   U94 : OAI21_X1 port map( B1 => n41, B2 => A(22), A => B(22), ZN => n92);
   U95 : AOI21_X1 port map( B1 => n45, B2 => n43, A => n93, ZN => n41);
   U96 : AOI21_X1 port map( B1 => n94, B2 => A(21), A => B(21), ZN => n93);
   U97 : INV_X1 port map( A => n43, ZN => n94);
   U98 : AOI22_X1 port map( A1 => n46, A2 => A(20), B1 => n95, B2 => B(20), ZN 
                           => n43);
   U99 : OR2_X1 port map( A1 => n46, A2 => A(20), ZN => n95);
   U100 : AOI21_X1 port map( B1 => n52, B2 => n50, A => n96, ZN => n46);
   U101 : AOI21_X1 port map( B1 => n97, B2 => A(19), A => B(19), ZN => n96);
   U102 : INV_X1 port map( A => n97, ZN => n50);
   U103 : OAI21_X1 port map( B1 => n53, B2 => n55, A => n98, ZN => n97);
   U104 : OAI21_X1 port map( B1 => n99, B2 => A(18), A => B(18), ZN => n98);
   U105 : INV_X1 port map( A => n53, ZN => n99);
   U106 : INV_X1 port map( A => A(18), ZN => n55);
   U107 : OAI21_X1 port map( B1 => A(17), B2 => n56, A => n100, ZN => n53);
   U108 : INV_X1 port map( A => n101, ZN => n100);
   U109 : AOI21_X1 port map( B1 => n56, B2 => A(17), A => B(17), ZN => n101);
   U110 : OAI21_X1 port map( B1 => n58, B2 => n60, A => n102, ZN => n56);
   U111 : OAI21_X1 port map( B1 => n103, B2 => A(16), A => B(16), ZN => n102);
   U112 : INV_X1 port map( A => n58, ZN => n103);
   U113 : INV_X1 port map( A => A(16), ZN => n60);
   U114 : OAI21_X1 port map( B1 => A(15), B2 => n61, A => n104, ZN => n58);
   U115 : INV_X1 port map( A => n105, ZN => n104);
   U116 : AOI21_X1 port map( B1 => n61, B2 => A(15), A => B(15), ZN => n105);
   U117 : OAI21_X1 port map( B1 => n63, B2 => n106, A => n107, ZN => n61);
   U118 : OAI21_X1 port map( B1 => n108, B2 => A(14), A => B(14), ZN => n107);
   U119 : INV_X1 port map( A => n63, ZN => n108);
   U120 : INV_X1 port map( A => A(14), ZN => n106);
   U121 : OAI21_X1 port map( B1 => A(13), B2 => n65, A => n109, ZN => n63);
   U122 : INV_X1 port map( A => n110, ZN => n109);
   U123 : AOI21_X1 port map( B1 => n65, B2 => A(13), A => B(13), ZN => n110);
   U124 : OAI21_X1 port map( B1 => n111, B2 => n112, A => n113, ZN => n65);
   U125 : OAI21_X1 port map( B1 => n67, B2 => A(12), A => B(12), ZN => n113);
   U126 : INV_X1 port map( A => n111, ZN => n67);
   U127 : INV_X1 port map( A => A(12), ZN => n112);
   U128 : OAI21_X1 port map( B1 => A(11), B2 => n69, A => n114, ZN => n111);
   U129 : INV_X1 port map( A => n115, ZN => n114);
   U130 : AOI21_X1 port map( B1 => n69, B2 => A(11), A => B(11), ZN => n115);
   U131 : OAI21_X1 port map( B1 => n116, B2 => n117, A => n118, ZN => n69);
   U132 : OAI21_X1 port map( B1 => n71, B2 => A(10), A => B(10), ZN => n118);
   U133 : INV_X1 port map( A => A(10), ZN => n117);
   U134 : INV_X1 port map( A => n71, ZN => n116);
   U135 : AOI21_X1 port map( B1 => n119, B2 => n1, A => n120, ZN => n71);
   U136 : AOI21_X1 port map( B1 => n121, B2 => A(9), A => B(9), ZN => n120);
   U137 : INV_X1 port map( A => n1, ZN => n121);
   U138 : AOI21_X1 port map( B1 => n3, B2 => A(8), A => n122, ZN => n1);
   U139 : INV_X1 port map( A => n123, ZN => n122);
   U140 : OAI21_X1 port map( B1 => n3, B2 => A(8), A => B(8), ZN => n123);
   U141 : AOI21_X1 port map( B1 => n7, B2 => n124, A => n125, ZN => n3);
   U142 : AOI21_X1 port map( B1 => n5, B2 => A(7), A => B(7), ZN => n125);
   U143 : INV_X1 port map( A => n124, ZN => n5);
   U144 : AOI21_X1 port map( B1 => n8, B2 => A(6), A => n126, ZN => n124);
   U145 : INV_X1 port map( A => n127, ZN => n126);
   U146 : OAI21_X1 port map( B1 => n8, B2 => A(6), A => B(6), ZN => n127);
   U147 : AOI21_X1 port map( B1 => n128, B2 => n129, A => n130, ZN => n8);
   U148 : AOI21_X1 port map( B1 => n10, B2 => A(5), A => B(5), ZN => n130);
   U149 : INV_X1 port map( A => n129, ZN => n10);
   U150 : AOI21_X1 port map( B1 => n12, B2 => A(4), A => n131, ZN => n129);
   U151 : INV_X1 port map( A => n132, ZN => n131);
   U152 : OAI21_X1 port map( B1 => n12, B2 => A(4), A => B(4), ZN => n132);
   U153 : AOI21_X1 port map( B1 => n16, B2 => n14, A => n133, ZN => n12);
   U154 : AOI21_X1 port map( B1 => n134, B2 => A(3), A => B(3), ZN => n133);
   U155 : INV_X1 port map( A => n14, ZN => n134);
   U156 : OAI22_X1 port map( A1 => A(2), A2 => n135, B1 => B(2), B2 => n136, ZN
                           => n14);
   U157 : AND2_X1 port map( A1 => n135, A2 => A(2), ZN => n136);
   U158 : INV_X1 port map( A => n22, ZN => n135);
   U159 : OAI22_X1 port map( A1 => A(1), A2 => n137, B1 => B(1), B2 => n138, ZN
                           => n22);
   U160 : AND2_X1 port map( A1 => n137, A2 => A(1), ZN => n138);
   U161 : INV_X1 port map( A => n48, ZN => n137);
   U162 : OAI21_X1 port map( B1 => B(0), B2 => A(0), A => n139, ZN => n48);
   U163 : INV_X1 port map( A => n140, ZN => n139);
   U164 : AOI21_X1 port map( B1 => A(0), B2 => B(0), A => Ci, ZN => n140);
   U165 : INV_X1 port map( A => A(3), ZN => n16);
   U166 : INV_X1 port map( A => A(5), ZN => n128);
   U167 : INV_X1 port map( A => A(7), ZN => n7);
   U168 : INV_X1 port map( A => A(9), ZN => n119);
   U169 : INV_X1 port map( A => A(19), ZN => n52);
   U170 : INV_X1 port map( A => A(21), ZN => n45);
   U171 : INV_X1 port map( A => A(23), ZN => n40);
   U172 : INV_X1 port map( A => A(25), ZN => n35);
   U173 : INV_X1 port map( A => A(30), ZN => n21);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX81_N32_3 is

   port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX81_N32_3;

architecture SYN_BEHAVIORAL of MUX81_N32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142 : std_logic;

begin
   
   U1 : OR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n142, ZN => n1);
   U2 : OR3_X1 port map( A1 => S(1), A2 => S(2), A3 => S(0), ZN => n2);
   U3 : OR3_X1 port map( A1 => n142, A2 => S(2), A3 => n141, ZN => n3);
   U4 : OR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n141, ZN => n4);
   U5 : AND3_X2 port map( A1 => S(2), A2 => S(1), A3 => S(0), ZN => n14);
   U6 : AND3_X2 port map( A1 => S(2), A2 => n142, A3 => S(0), ZN => n16);
   U7 : AND3_X2 port map( A1 => S(1), A2 => n141, A3 => S(2), ZN => n13);
   U8 : AND3_X2 port map( A1 => n141, A2 => n142, A3 => S(2), ZN => n15);
   U9 : INV_X2 port map( A => n3, ZN => n5);
   U10 : INV_X2 port map( A => n4, ZN => n6);
   U11 : INV_X2 port map( A => n1, ZN => n7);
   U12 : INV_X2 port map( A => n2, ZN => n8);
   U13 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => 
                           Y(9));
   U14 : AOI22_X1 port map( A1 => G(9), A2 => n13, B1 => H(9), B2 => n14, ZN =>
                           n12);
   U15 : AOI22_X1 port map( A1 => E(9), A2 => n15, B1 => F(9), B2 => n16, ZN =>
                           n11);
   U16 : AOI22_X1 port map( A1 => C(9), A2 => n7, B1 => D(9), B2 => n5, ZN => 
                           n10);
   U17 : AOI22_X1 port map( A1 => A(9), A2 => n8, B1 => B(9), B2 => n6, ZN => 
                           n9);
   U18 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           Y(8));
   U19 : AOI22_X1 port map( A1 => G(8), A2 => n13, B1 => H(8), B2 => n14, ZN =>
                           n20);
   U20 : AOI22_X1 port map( A1 => E(8), A2 => n15, B1 => F(8), B2 => n16, ZN =>
                           n19);
   U21 : AOI22_X1 port map( A1 => C(8), A2 => n7, B1 => D(8), B2 => n5, ZN => 
                           n18);
   U22 : AOI22_X1 port map( A1 => A(8), A2 => n8, B1 => B(8), B2 => n6, ZN => 
                           n17);
   U23 : NAND4_X1 port map( A1 => n21, A2 => n22, A3 => n23, A4 => n24, ZN => 
                           Y(7));
   U24 : AOI22_X1 port map( A1 => G(7), A2 => n13, B1 => H(7), B2 => n14, ZN =>
                           n24);
   U25 : AOI22_X1 port map( A1 => E(7), A2 => n15, B1 => F(7), B2 => n16, ZN =>
                           n23);
   U26 : AOI22_X1 port map( A1 => C(7), A2 => n7, B1 => D(7), B2 => n5, ZN => 
                           n22);
   U27 : AOI22_X1 port map( A1 => A(7), A2 => n8, B1 => B(7), B2 => n6, ZN => 
                           n21);
   U28 : NAND4_X1 port map( A1 => n25, A2 => n26, A3 => n27, A4 => n28, ZN => 
                           Y(6));
   U29 : AOI22_X1 port map( A1 => G(6), A2 => n13, B1 => H(6), B2 => n14, ZN =>
                           n28);
   U30 : AOI22_X1 port map( A1 => E(6), A2 => n15, B1 => F(6), B2 => n16, ZN =>
                           n27);
   U31 : AOI22_X1 port map( A1 => C(6), A2 => n7, B1 => D(6), B2 => n5, ZN => 
                           n26);
   U32 : AOI22_X1 port map( A1 => A(6), A2 => n8, B1 => B(6), B2 => n6, ZN => 
                           n25);
   U33 : NAND4_X1 port map( A1 => n29, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           Y(5));
   U34 : AOI22_X1 port map( A1 => G(5), A2 => n13, B1 => H(5), B2 => n14, ZN =>
                           n32);
   U35 : AOI22_X1 port map( A1 => E(5), A2 => n15, B1 => F(5), B2 => n16, ZN =>
                           n31);
   U36 : AOI22_X1 port map( A1 => C(5), A2 => n7, B1 => D(5), B2 => n5, ZN => 
                           n30);
   U37 : AOI22_X1 port map( A1 => A(5), A2 => n8, B1 => B(5), B2 => n6, ZN => 
                           n29);
   U38 : NAND4_X1 port map( A1 => n33, A2 => n34, A3 => n35, A4 => n36, ZN => 
                           Y(4));
   U39 : AOI22_X1 port map( A1 => G(4), A2 => n13, B1 => H(4), B2 => n14, ZN =>
                           n36);
   U40 : AOI22_X1 port map( A1 => E(4), A2 => n15, B1 => F(4), B2 => n16, ZN =>
                           n35);
   U41 : AOI22_X1 port map( A1 => C(4), A2 => n7, B1 => D(4), B2 => n5, ZN => 
                           n34);
   U42 : AOI22_X1 port map( A1 => A(4), A2 => n8, B1 => B(4), B2 => n6, ZN => 
                           n33);
   U43 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           Y(3));
   U44 : AOI22_X1 port map( A1 => G(3), A2 => n13, B1 => H(3), B2 => n14, ZN =>
                           n40);
   U45 : AOI22_X1 port map( A1 => E(3), A2 => n15, B1 => F(3), B2 => n16, ZN =>
                           n39);
   U46 : AOI22_X1 port map( A1 => C(3), A2 => n7, B1 => D(3), B2 => n5, ZN => 
                           n38);
   U47 : AOI22_X1 port map( A1 => A(3), A2 => n8, B1 => B(3), B2 => n6, ZN => 
                           n37);
   U48 : NAND4_X1 port map( A1 => n41, A2 => n42, A3 => n43, A4 => n44, ZN => 
                           Y(31));
   U49 : AOI22_X1 port map( A1 => G(31), A2 => n13, B1 => H(31), B2 => n14, ZN 
                           => n44);
   U50 : AOI22_X1 port map( A1 => E(31), A2 => n15, B1 => F(31), B2 => n16, ZN 
                           => n43);
   U51 : AOI22_X1 port map( A1 => C(31), A2 => n7, B1 => D(31), B2 => n5, ZN =>
                           n42);
   U52 : AOI22_X1 port map( A1 => A(31), A2 => n8, B1 => B(31), B2 => n6, ZN =>
                           n41);
   U53 : NAND4_X1 port map( A1 => n45, A2 => n46, A3 => n47, A4 => n48, ZN => 
                           Y(30));
   U54 : AOI22_X1 port map( A1 => G(30), A2 => n13, B1 => H(30), B2 => n14, ZN 
                           => n48);
   U55 : AOI22_X1 port map( A1 => E(30), A2 => n15, B1 => F(30), B2 => n16, ZN 
                           => n47);
   U56 : AOI22_X1 port map( A1 => C(30), A2 => n7, B1 => D(30), B2 => n5, ZN =>
                           n46);
   U57 : AOI22_X1 port map( A1 => A(30), A2 => n8, B1 => B(30), B2 => n6, ZN =>
                           n45);
   U58 : NAND4_X1 port map( A1 => n49, A2 => n50, A3 => n51, A4 => n52, ZN => 
                           Y(2));
   U59 : AOI22_X1 port map( A1 => G(2), A2 => n13, B1 => H(2), B2 => n14, ZN =>
                           n52);
   U60 : AOI22_X1 port map( A1 => E(2), A2 => n15, B1 => F(2), B2 => n16, ZN =>
                           n51);
   U61 : AOI22_X1 port map( A1 => C(2), A2 => n7, B1 => D(2), B2 => n5, ZN => 
                           n50);
   U62 : AOI22_X1 port map( A1 => A(2), A2 => n8, B1 => B(2), B2 => n6, ZN => 
                           n49);
   U63 : NAND4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           Y(29));
   U64 : AOI22_X1 port map( A1 => G(29), A2 => n13, B1 => H(29), B2 => n14, ZN 
                           => n56);
   U65 : AOI22_X1 port map( A1 => E(29), A2 => n15, B1 => F(29), B2 => n16, ZN 
                           => n55);
   U66 : AOI22_X1 port map( A1 => C(29), A2 => n7, B1 => D(29), B2 => n5, ZN =>
                           n54);
   U67 : AOI22_X1 port map( A1 => A(29), A2 => n8, B1 => B(29), B2 => n6, ZN =>
                           n53);
   U68 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           Y(28));
   U69 : AOI22_X1 port map( A1 => G(28), A2 => n13, B1 => H(28), B2 => n14, ZN 
                           => n60);
   U70 : AOI22_X1 port map( A1 => E(28), A2 => n15, B1 => F(28), B2 => n16, ZN 
                           => n59);
   U71 : AOI22_X1 port map( A1 => C(28), A2 => n7, B1 => D(28), B2 => n5, ZN =>
                           n58);
   U72 : AOI22_X1 port map( A1 => A(28), A2 => n8, B1 => B(28), B2 => n6, ZN =>
                           n57);
   U73 : NAND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           Y(27));
   U74 : AOI22_X1 port map( A1 => G(27), A2 => n13, B1 => H(27), B2 => n14, ZN 
                           => n64);
   U75 : AOI22_X1 port map( A1 => E(27), A2 => n15, B1 => F(27), B2 => n16, ZN 
                           => n63);
   U76 : AOI22_X1 port map( A1 => C(27), A2 => n7, B1 => D(27), B2 => n5, ZN =>
                           n62);
   U77 : AOI22_X1 port map( A1 => A(27), A2 => n8, B1 => B(27), B2 => n6, ZN =>
                           n61);
   U78 : NAND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n68, ZN => 
                           Y(26));
   U79 : AOI22_X1 port map( A1 => G(26), A2 => n13, B1 => H(26), B2 => n14, ZN 
                           => n68);
   U80 : AOI22_X1 port map( A1 => E(26), A2 => n15, B1 => F(26), B2 => n16, ZN 
                           => n67);
   U81 : AOI22_X1 port map( A1 => C(26), A2 => n7, B1 => D(26), B2 => n5, ZN =>
                           n66);
   U82 : AOI22_X1 port map( A1 => A(26), A2 => n8, B1 => B(26), B2 => n6, ZN =>
                           n65);
   U83 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           Y(25));
   U84 : AOI22_X1 port map( A1 => G(25), A2 => n13, B1 => H(25), B2 => n14, ZN 
                           => n72);
   U85 : AOI22_X1 port map( A1 => E(25), A2 => n15, B1 => F(25), B2 => n16, ZN 
                           => n71);
   U86 : AOI22_X1 port map( A1 => C(25), A2 => n7, B1 => D(25), B2 => n5, ZN =>
                           n70);
   U87 : AOI22_X1 port map( A1 => A(25), A2 => n8, B1 => B(25), B2 => n6, ZN =>
                           n69);
   U88 : NAND4_X1 port map( A1 => n73, A2 => n74, A3 => n75, A4 => n76, ZN => 
                           Y(24));
   U89 : AOI22_X1 port map( A1 => G(24), A2 => n13, B1 => H(24), B2 => n14, ZN 
                           => n76);
   U90 : AOI22_X1 port map( A1 => E(24), A2 => n15, B1 => F(24), B2 => n16, ZN 
                           => n75);
   U91 : AOI22_X1 port map( A1 => C(24), A2 => n7, B1 => D(24), B2 => n5, ZN =>
                           n74);
   U92 : AOI22_X1 port map( A1 => A(24), A2 => n8, B1 => B(24), B2 => n6, ZN =>
                           n73);
   U93 : NAND4_X1 port map( A1 => n77, A2 => n78, A3 => n79, A4 => n80, ZN => 
                           Y(23));
   U94 : AOI22_X1 port map( A1 => G(23), A2 => n13, B1 => H(23), B2 => n14, ZN 
                           => n80);
   U95 : AOI22_X1 port map( A1 => E(23), A2 => n15, B1 => F(23), B2 => n16, ZN 
                           => n79);
   U96 : AOI22_X1 port map( A1 => C(23), A2 => n7, B1 => D(23), B2 => n5, ZN =>
                           n78);
   U97 : AOI22_X1 port map( A1 => A(23), A2 => n8, B1 => B(23), B2 => n6, ZN =>
                           n77);
   U98 : NAND4_X1 port map( A1 => n81, A2 => n82, A3 => n83, A4 => n84, ZN => 
                           Y(22));
   U99 : AOI22_X1 port map( A1 => G(22), A2 => n13, B1 => H(22), B2 => n14, ZN 
                           => n84);
   U100 : AOI22_X1 port map( A1 => E(22), A2 => n15, B1 => F(22), B2 => n16, ZN
                           => n83);
   U101 : AOI22_X1 port map( A1 => C(22), A2 => n7, B1 => D(22), B2 => n5, ZN 
                           => n82);
   U102 : AOI22_X1 port map( A1 => A(22), A2 => n8, B1 => B(22), B2 => n6, ZN 
                           => n81);
   U103 : NAND4_X1 port map( A1 => n85, A2 => n86, A3 => n87, A4 => n88, ZN => 
                           Y(21));
   U104 : AOI22_X1 port map( A1 => G(21), A2 => n13, B1 => H(21), B2 => n14, ZN
                           => n88);
   U105 : AOI22_X1 port map( A1 => E(21), A2 => n15, B1 => F(21), B2 => n16, ZN
                           => n87);
   U106 : AOI22_X1 port map( A1 => C(21), A2 => n7, B1 => D(21), B2 => n5, ZN 
                           => n86);
   U107 : AOI22_X1 port map( A1 => A(21), A2 => n8, B1 => B(21), B2 => n6, ZN 
                           => n85);
   U108 : NAND4_X1 port map( A1 => n89, A2 => n90, A3 => n91, A4 => n92, ZN => 
                           Y(20));
   U109 : AOI22_X1 port map( A1 => G(20), A2 => n13, B1 => H(20), B2 => n14, ZN
                           => n92);
   U110 : AOI22_X1 port map( A1 => E(20), A2 => n15, B1 => F(20), B2 => n16, ZN
                           => n91);
   U111 : AOI22_X1 port map( A1 => C(20), A2 => n7, B1 => D(20), B2 => n5, ZN 
                           => n90);
   U112 : AOI22_X1 port map( A1 => A(20), A2 => n8, B1 => B(20), B2 => n6, ZN 
                           => n89);
   U113 : NAND4_X1 port map( A1 => n93, A2 => n94, A3 => n95, A4 => n96, ZN => 
                           Y(1));
   U114 : AOI22_X1 port map( A1 => G(1), A2 => n13, B1 => H(1), B2 => n14, ZN 
                           => n96);
   U115 : AOI22_X1 port map( A1 => E(1), A2 => n15, B1 => F(1), B2 => n16, ZN 
                           => n95);
   U116 : AOI22_X1 port map( A1 => C(1), A2 => n7, B1 => D(1), B2 => n5, ZN => 
                           n94);
   U117 : AOI22_X1 port map( A1 => A(1), A2 => n8, B1 => B(1), B2 => n6, ZN => 
                           n93);
   U118 : NAND4_X1 port map( A1 => n97, A2 => n98, A3 => n99, A4 => n100, ZN =>
                           Y(19));
   U119 : AOI22_X1 port map( A1 => G(19), A2 => n13, B1 => H(19), B2 => n14, ZN
                           => n100);
   U120 : AOI22_X1 port map( A1 => E(19), A2 => n15, B1 => F(19), B2 => n16, ZN
                           => n99);
   U121 : AOI22_X1 port map( A1 => C(19), A2 => n7, B1 => D(19), B2 => n5, ZN 
                           => n98);
   U122 : AOI22_X1 port map( A1 => A(19), A2 => n8, B1 => B(19), B2 => n6, ZN 
                           => n97);
   U123 : NAND4_X1 port map( A1 => n101, A2 => n102, A3 => n103, A4 => n104, ZN
                           => Y(18));
   U124 : AOI22_X1 port map( A1 => G(18), A2 => n13, B1 => H(18), B2 => n14, ZN
                           => n104);
   U125 : AOI22_X1 port map( A1 => E(18), A2 => n15, B1 => F(18), B2 => n16, ZN
                           => n103);
   U126 : AOI22_X1 port map( A1 => C(18), A2 => n7, B1 => D(18), B2 => n5, ZN 
                           => n102);
   U127 : AOI22_X1 port map( A1 => A(18), A2 => n8, B1 => B(18), B2 => n6, ZN 
                           => n101);
   U128 : NAND4_X1 port map( A1 => n105, A2 => n106, A3 => n107, A4 => n108, ZN
                           => Y(17));
   U129 : AOI22_X1 port map( A1 => G(17), A2 => n13, B1 => H(17), B2 => n14, ZN
                           => n108);
   U130 : AOI22_X1 port map( A1 => E(17), A2 => n15, B1 => F(17), B2 => n16, ZN
                           => n107);
   U131 : AOI22_X1 port map( A1 => C(17), A2 => n7, B1 => D(17), B2 => n5, ZN 
                           => n106);
   U132 : AOI22_X1 port map( A1 => A(17), A2 => n8, B1 => B(17), B2 => n6, ZN 
                           => n105);
   U133 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n111, A4 => n112, ZN
                           => Y(16));
   U134 : AOI22_X1 port map( A1 => G(16), A2 => n13, B1 => H(16), B2 => n14, ZN
                           => n112);
   U135 : AOI22_X1 port map( A1 => E(16), A2 => n15, B1 => F(16), B2 => n16, ZN
                           => n111);
   U136 : AOI22_X1 port map( A1 => C(16), A2 => n7, B1 => D(16), B2 => n5, ZN 
                           => n110);
   U137 : AOI22_X1 port map( A1 => A(16), A2 => n8, B1 => B(16), B2 => n6, ZN 
                           => n109);
   U138 : NAND4_X1 port map( A1 => n113, A2 => n114, A3 => n115, A4 => n116, ZN
                           => Y(15));
   U139 : AOI22_X1 port map( A1 => G(15), A2 => n13, B1 => H(15), B2 => n14, ZN
                           => n116);
   U140 : AOI22_X1 port map( A1 => E(15), A2 => n15, B1 => F(15), B2 => n16, ZN
                           => n115);
   U141 : AOI22_X1 port map( A1 => C(15), A2 => n7, B1 => D(15), B2 => n5, ZN 
                           => n114);
   U142 : AOI22_X1 port map( A1 => A(15), A2 => n8, B1 => B(15), B2 => n6, ZN 
                           => n113);
   U143 : NAND4_X1 port map( A1 => n117, A2 => n118, A3 => n119, A4 => n120, ZN
                           => Y(14));
   U144 : AOI22_X1 port map( A1 => G(14), A2 => n13, B1 => H(14), B2 => n14, ZN
                           => n120);
   U145 : AOI22_X1 port map( A1 => E(14), A2 => n15, B1 => F(14), B2 => n16, ZN
                           => n119);
   U146 : AOI22_X1 port map( A1 => C(14), A2 => n7, B1 => D(14), B2 => n5, ZN 
                           => n118);
   U147 : AOI22_X1 port map( A1 => A(14), A2 => n8, B1 => B(14), B2 => n6, ZN 
                           => n117);
   U148 : NAND4_X1 port map( A1 => n121, A2 => n122, A3 => n123, A4 => n124, ZN
                           => Y(13));
   U149 : AOI22_X1 port map( A1 => G(13), A2 => n13, B1 => H(13), B2 => n14, ZN
                           => n124);
   U150 : AOI22_X1 port map( A1 => E(13), A2 => n15, B1 => F(13), B2 => n16, ZN
                           => n123);
   U151 : AOI22_X1 port map( A1 => C(13), A2 => n7, B1 => D(13), B2 => n5, ZN 
                           => n122);
   U152 : AOI22_X1 port map( A1 => A(13), A2 => n8, B1 => B(13), B2 => n6, ZN 
                           => n121);
   U153 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => Y(12));
   U154 : AOI22_X1 port map( A1 => G(12), A2 => n13, B1 => H(12), B2 => n14, ZN
                           => n128);
   U155 : AOI22_X1 port map( A1 => E(12), A2 => n15, B1 => F(12), B2 => n16, ZN
                           => n127);
   U156 : AOI22_X1 port map( A1 => C(12), A2 => n7, B1 => D(12), B2 => n5, ZN 
                           => n126);
   U157 : AOI22_X1 port map( A1 => A(12), A2 => n8, B1 => B(12), B2 => n6, ZN 
                           => n125);
   U158 : NAND4_X1 port map( A1 => n129, A2 => n130, A3 => n131, A4 => n132, ZN
                           => Y(11));
   U159 : AOI22_X1 port map( A1 => G(11), A2 => n13, B1 => H(11), B2 => n14, ZN
                           => n132);
   U160 : AOI22_X1 port map( A1 => E(11), A2 => n15, B1 => F(11), B2 => n16, ZN
                           => n131);
   U161 : AOI22_X1 port map( A1 => C(11), A2 => n7, B1 => D(11), B2 => n5, ZN 
                           => n130);
   U162 : AOI22_X1 port map( A1 => A(11), A2 => n8, B1 => B(11), B2 => n6, ZN 
                           => n129);
   U163 : NAND4_X1 port map( A1 => n133, A2 => n134, A3 => n135, A4 => n136, ZN
                           => Y(10));
   U164 : AOI22_X1 port map( A1 => G(10), A2 => n13, B1 => H(10), B2 => n14, ZN
                           => n136);
   U165 : AOI22_X1 port map( A1 => E(10), A2 => n15, B1 => F(10), B2 => n16, ZN
                           => n135);
   U166 : AOI22_X1 port map( A1 => C(10), A2 => n7, B1 => D(10), B2 => n5, ZN 
                           => n134);
   U167 : AOI22_X1 port map( A1 => A(10), A2 => n8, B1 => B(10), B2 => n6, ZN 
                           => n133);
   U168 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => Y(0));
   U169 : AOI22_X1 port map( A1 => G(0), A2 => n13, B1 => H(0), B2 => n14, ZN 
                           => n140);
   U170 : AOI22_X1 port map( A1 => E(0), A2 => n15, B1 => F(0), B2 => n16, ZN 
                           => n139);
   U171 : AOI22_X1 port map( A1 => C(0), A2 => n7, B1 => D(0), B2 => n5, ZN => 
                           n138);
   U172 : INV_X1 port map( A => S(1), ZN => n142);
   U173 : AOI22_X1 port map( A1 => A(0), A2 => n8, B1 => B(0), B2 => n6, ZN => 
                           n137);
   U174 : INV_X1 port map( A => S(0), ZN => n141);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BOOTH_ENCODER_N16 is

   port( B : in std_logic_vector (15 downto 0);  Bo : out std_logic_vector (23 
         downto 0));

end BOOTH_ENCODER_N16;

architecture SYN_STRUCTURAL of BOOTH_ENCODER_N16 is

   component ENCODER_0
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_1
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_2
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_3
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_4
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_5
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_6
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component ENCODER_7
      port( B : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   ENC_0 : ENCODER_7 port map( B(2) => B(1), B(1) => B(0), B(0) => 
                           X_Logic0_port, Y(2) => Bo(2), Y(1) => Bo(1), Y(0) =>
                           Bo(0));
   ENC_1 : ENCODER_6 port map( B(2) => B(3), B(1) => B(2), B(0) => B(1), Y(2) 
                           => Bo(5), Y(1) => Bo(4), Y(0) => Bo(3));
   ENC_2 : ENCODER_5 port map( B(2) => B(5), B(1) => B(4), B(0) => B(3), Y(2) 
                           => Bo(8), Y(1) => Bo(7), Y(0) => Bo(6));
   ENC_3 : ENCODER_4 port map( B(2) => B(7), B(1) => B(6), B(0) => B(5), Y(2) 
                           => Bo(11), Y(1) => Bo(10), Y(0) => Bo(9));
   ENC_4 : ENCODER_3 port map( B(2) => B(9), B(1) => B(8), B(0) => B(7), Y(2) 
                           => Bo(14), Y(1) => Bo(13), Y(0) => Bo(12));
   ENC_5 : ENCODER_2 port map( B(2) => B(11), B(1) => B(10), B(0) => B(9), Y(2)
                           => Bo(17), Y(1) => Bo(16), Y(0) => Bo(15));
   ENC_6 : ENCODER_1 port map( B(2) => B(13), B(1) => B(12), B(0) => B(11), 
                           Y(2) => Bo(20), Y(1) => Bo(19), Y(0) => Bo(18));
   ENC_7 : ENCODER_0 port map( B(2) => B(15), B(1) => B(14), B(0) => B(13), 
                           Y(2) => Bo(23), Y(1) => Bo(22), Y(0) => Bo(21));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GENERATOR_N32_NB8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_N32_NB8;

architecture SYN_STRUCTURAL of SUM_GENERATOR_N32_NB8 is

   component CSB_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_1 : CSB_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => Ci(0), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   CSBI_2 : CSB_N4_6 port map( A(3) => A(7), A(2) => A(6), A(1) => A(5), A(0) 
                           => A(4), B(3) => B(7), B(2) => B(6), B(1) => B(5), 
                           B(0) => B(4), Ci => Ci(1), S(3) => S(7), S(2) => 
                           S(6), S(1) => S(5), S(0) => S(4));
   CSBI_3 : CSB_N4_5 port map( A(3) => A(11), A(2) => A(10), A(1) => A(9), A(0)
                           => A(8), B(3) => B(11), B(2) => B(10), B(1) => B(9),
                           B(0) => B(8), Ci => Ci(2), S(3) => S(11), S(2) => 
                           S(10), S(1) => S(9), S(0) => S(8));
   CSBI_4 : CSB_N4_4 port map( A(3) => A(15), A(2) => A(14), A(1) => A(13), 
                           A(0) => A(12), B(3) => B(15), B(2) => B(14), B(1) =>
                           B(13), B(0) => B(12), Ci => Ci(3), S(3) => S(15), 
                           S(2) => S(14), S(1) => S(13), S(0) => S(12));
   CSBI_5 : CSB_N4_3 port map( A(3) => A(19), A(2) => A(18), A(1) => A(17), 
                           A(0) => A(16), B(3) => B(19), B(2) => B(18), B(1) =>
                           B(17), B(0) => B(16), Ci => Ci(4), S(3) => S(19), 
                           S(2) => S(18), S(1) => S(17), S(0) => S(16));
   CSBI_6 : CSB_N4_2 port map( A(3) => A(23), A(2) => A(22), A(1) => A(21), 
                           A(0) => A(20), B(3) => B(23), B(2) => B(22), B(1) =>
                           B(21), B(0) => B(20), Ci => Ci(5), S(3) => S(23), 
                           S(2) => S(22), S(1) => S(21), S(0) => S(20));
   CSBI_7 : CSB_N4_1 port map( A(3) => A(27), A(2) => A(26), A(1) => A(25), 
                           A(0) => A(24), B(3) => B(27), B(2) => B(26), B(1) =>
                           B(25), B(0) => B(24), Ci => Ci(6), S(3) => S(27), 
                           S(2) => S(26), S(1) => S(25), S(0) => S(24));
   CSBI_8 : CSB_N4_0 port map( A(3) => A(31), A(2) => A(30), A(1) => A(29), 
                           A(0) => A(28), B(3) => B(31), B(2) => B(30), B(1) =>
                           B(29), B(0) => B(28), Ci => Ci(7), S(3) => S(31), 
                           S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CARRY_GENERATOR_N32_NB8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_N32_NB8;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_N32_NB8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component PG_BLOCK_0
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_0
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_1
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_1
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_2
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_2
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_3
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_3
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_4
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_5
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_6
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_4
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_7
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_5
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_8
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_9
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_10
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_11
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_6
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_12
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_13
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_14
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_15
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_16
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_17
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_18
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_7
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_BLOCK_19
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_20
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_21
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_22
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_23
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_24
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_25
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_26
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_27
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_28
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_29
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_30
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_31
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_32
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component PG_BLOCK_33
      port( Gik, Gkj, Pik, Pkj : in std_logic;  Gij, Pij : out std_logic);
   end component;
   
   component GENERATE_BLOCK_8
      port( Gik, Gkj, Pik : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_ROW_N32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  P, G
            : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port,
      Co_2_port, Co_1_port, Co_0_port, G_4_31_port, G_4_27_port, G_4_23_port, 
      G_3_31_port, G_3_27_port, G_3_19_port, G_3_15_port, G_3_11_port, 
      G_2_31_port, G_2_23_port, G_2_15_port, G_2_7_port, G_1_31_port, 
      G_1_29_port, G_1_27_port, G_1_25_port, G_1_23_port, G_1_21_port, 
      G_1_19_port, G_1_17_port, G_1_15_port, G_1_13_port, G_1_11_port, 
      G_1_9_port, G_1_7_port, G_1_5_port, G_1_3_port, G_1_1_port, G_0_31_port, 
      G_0_30_port, G_0_29_port, G_0_28_port, G_0_27_port, G_0_26_port, 
      G_0_25_port, G_0_24_port, G_0_23_port, G_0_22_port, G_0_21_port, 
      G_0_20_port, G_0_19_port, G_0_18_port, G_0_17_port, G_0_16_port, 
      G_0_15_port, G_0_14_port, G_0_13_port, G_0_12_port, G_0_11_port, 
      G_0_10_port, G_0_9_port, G_0_8_port, G_0_7_port, G_0_6_port, G_0_5_port, 
      G_0_4_port, G_0_3_port, G_0_2_port, G_0_1_port, G_0_0_port, P_5_15_port, 
      P_4_31_port, P_4_27_port, P_4_23_port, P_4_7_port, P_3_31_port, 
      P_3_27_port, P_3_19_port, P_3_15_port, P_3_11_port, P_2_31_port, 
      P_2_23_port, P_2_15_port, P_2_7_port, P_1_31_port, P_1_29_port, 
      P_1_27_port, P_1_25_port, P_1_23_port, P_1_21_port, P_1_19_port, 
      P_1_17_port, P_1_15_port, P_1_13_port, P_1_11_port, P_1_9_port, 
      P_1_7_port, P_1_5_port, P_1_3_port, P_0_31_port, P_0_30_port, P_0_29_port
      , P_0_28_port, P_0_27_port, P_0_26_port, P_0_25_port, P_0_24_port, 
      P_0_23_port, P_0_22_port, P_0_21_port, P_0_20_port, P_0_19_port, 
      P_0_18_port, P_0_17_port, P_0_16_port, P_0_15_port, P_0_14_port, 
      P_0_13_port, P_0_12_port, P_0_11_port, P_0_10_port, P_0_9_port, 
      P_0_8_port, P_0_7_port, P_0_6_port, P_0_5_port, P_0_4_port, P_0_3_port, 
      P_0_2_port, P_0_1_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12
      , n13, n14, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   X_Logic0_port <= '0';
   PG_ROW_INSTANCE : PG_ROW_N32 port map( A(31) => A(31), A(30) => A(30), A(29)
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => Ci, P(31) => P_0_31_port, P(30) => 
                           P_0_30_port, P(29) => P_0_29_port, P(28) => 
                           P_0_28_port, P(27) => P_0_27_port, P(26) => 
                           P_0_26_port, P(25) => P_0_25_port, P(24) => 
                           P_0_24_port, P(23) => P_0_23_port, P(22) => 
                           P_0_22_port, P(21) => P_0_21_port, P(20) => 
                           P_0_20_port, P(19) => P_0_19_port, P(18) => 
                           P_0_18_port, P(17) => P_0_17_port, P(16) => 
                           P_0_16_port, P(15) => P_0_15_port, P(14) => 
                           P_0_14_port, P(13) => P_0_13_port, P(12) => 
                           P_0_12_port, P(11) => P_0_11_port, P(10) => 
                           P_0_10_port, P(9) => P_0_9_port, P(8) => P_0_8_port,
                           P(7) => P_0_7_port, P(6) => P_0_6_port, P(5) => 
                           P_0_5_port, P(4) => P_0_4_port, P(3) => P_0_3_port, 
                           P(2) => P_0_2_port, P(1) => P_0_1_port, P(0) => 
                           n_1255, G(31) => G_0_31_port, G(30) => G_0_30_port, 
                           G(29) => G_0_29_port, G(28) => G_0_28_port, G(27) =>
                           G_0_27_port, G(26) => G_0_26_port, G(25) => 
                           G_0_25_port, G(24) => G_0_24_port, G(23) => 
                           G_0_23_port, G(22) => G_0_22_port, G(21) => 
                           G_0_21_port, G(20) => G_0_20_port, G(19) => 
                           G_0_19_port, G(18) => G_0_18_port, G(17) => 
                           G_0_17_port, G(16) => G_0_16_port, G(15) => 
                           G_0_15_port, G(14) => G_0_14_port, G(13) => 
                           G_0_13_port, G(12) => G_0_12_port, G(11) => 
                           G_0_11_port, G(10) => G_0_10_port, G(9) => 
                           G_0_9_port, G(8) => G_0_8_port, G(7) => G_0_7_port, 
                           G(6) => G_0_6_port, G(5) => G_0_5_port, G(4) => 
                           G_0_4_port, G(3) => G_0_3_port, G(2) => G_0_2_port, 
                           G(1) => G_0_1_port, G(0) => G_0_0_port);
   G_BLOCK_INSTANCE_1_1 : GENERATE_BLOCK_8 port map( Gik => G_0_1_port, Gkj => 
                           G_0_0_port, Pik => P_0_1_port, Gij => G_1_1_port);
   PG_BLOCK_REG_INSTANCE_1_3 : PG_BLOCK_33 port map( Gik => G_0_3_port, Gkj => 
                           G_0_2_port, Pik => P_0_3_port, Pkj => P_0_2_port, 
                           Gij => G_1_3_port, Pij => P_1_3_port);
   PG_BLOCK_REG_INSTANCE_1_5 : PG_BLOCK_32 port map( Gik => G_0_5_port, Gkj => 
                           G_0_4_port, Pik => P_0_5_port, Pkj => P_0_4_port, 
                           Gij => G_1_5_port, Pij => P_1_5_port);
   PG_BLOCK_REG_INSTANCE_1_7 : PG_BLOCK_31 port map( Gik => G_0_7_port, Gkj => 
                           G_0_6_port, Pik => P_0_7_port, Pkj => P_0_6_port, 
                           Gij => G_1_7_port, Pij => P_1_7_port);
   PG_BLOCK_REG_INSTANCE_1_9 : PG_BLOCK_30 port map( Gik => G_0_9_port, Gkj => 
                           G_0_8_port, Pik => P_0_9_port, Pkj => P_0_8_port, 
                           Gij => G_1_9_port, Pij => P_1_9_port);
   PG_BLOCK_REG_INSTANCE_1_11 : PG_BLOCK_29 port map( Gik => G_0_11_port, Gkj 
                           => G_0_10_port, Pik => P_0_11_port, Pkj => 
                           P_0_10_port, Gij => G_1_11_port, Pij => P_1_11_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_13 : PG_BLOCK_28 port map( Gik => G_0_13_port, Gkj 
                           => G_0_12_port, Pik => P_0_13_port, Pkj => 
                           P_0_12_port, Gij => G_1_13_port, Pij => P_1_13_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_15 : PG_BLOCK_27 port map( Gik => G_0_15_port, Gkj 
                           => G_0_14_port, Pik => P_0_15_port, Pkj => 
                           P_0_14_port, Gij => G_1_15_port, Pij => P_1_15_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_17 : PG_BLOCK_26 port map( Gik => G_0_17_port, Gkj 
                           => G_0_16_port, Pik => P_0_17_port, Pkj => 
                           P_0_16_port, Gij => G_1_17_port, Pij => P_1_17_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_19 : PG_BLOCK_25 port map( Gik => G_0_19_port, Gkj 
                           => G_0_18_port, Pik => P_0_19_port, Pkj => 
                           P_0_18_port, Gij => G_1_19_port, Pij => P_1_19_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_21 : PG_BLOCK_24 port map( Gik => G_0_21_port, Gkj 
                           => G_0_20_port, Pik => P_0_21_port, Pkj => 
                           P_0_20_port, Gij => G_1_21_port, Pij => P_1_21_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_23 : PG_BLOCK_23 port map( Gik => G_0_23_port, Gkj 
                           => G_0_22_port, Pik => P_0_23_port, Pkj => 
                           P_0_22_port, Gij => G_1_23_port, Pij => P_1_23_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_25 : PG_BLOCK_22 port map( Gik => G_0_25_port, Gkj 
                           => G_0_24_port, Pik => P_0_25_port, Pkj => 
                           P_0_24_port, Gij => G_1_25_port, Pij => P_1_25_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_27 : PG_BLOCK_21 port map( Gik => G_0_27_port, Gkj 
                           => G_0_26_port, Pik => P_0_27_port, Pkj => 
                           P_0_26_port, Gij => G_1_27_port, Pij => P_1_27_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_29 : PG_BLOCK_20 port map( Gik => G_0_29_port, Gkj 
                           => G_0_28_port, Pik => P_0_29_port, Pkj => 
                           P_0_28_port, Gij => G_1_29_port, Pij => P_1_29_port)
                           ;
   PG_BLOCK_REG_INSTANCE_1_31 : PG_BLOCK_19 port map( Gik => G_0_31_port, Gkj 
                           => G_0_30_port, Pik => P_0_31_port, Pkj => 
                           P_0_30_port, Gij => G_1_31_port, Pij => P_1_31_port)
                           ;
   G_BLOCK_INSTANCE_2_3 : GENERATE_BLOCK_7 port map( Gik => G_1_3_port, Gkj => 
                           G_1_1_port, Pik => P_1_3_port, Gij => Co_0_port);
   PG_BLOCK_REG_INSTANCE_2_7 : PG_BLOCK_18 port map( Gik => G_1_7_port, Gkj => 
                           G_1_5_port, Pik => P_1_7_port, Pkj => P_1_5_port, 
                           Gij => G_2_7_port, Pij => P_2_7_port);
   PG_BLOCK_REG_INSTANCE_2_11 : PG_BLOCK_17 port map( Gik => G_1_11_port, Gkj 
                           => G_1_9_port, Pik => P_1_11_port, Pkj => P_1_9_port
                           , Gij => G_3_11_port, Pij => P_3_11_port);
   PG_BLOCK_REG_INSTANCE_2_15 : PG_BLOCK_16 port map( Gik => G_1_15_port, Gkj 
                           => G_1_13_port, Pik => P_1_15_port, Pkj => 
                           P_1_13_port, Gij => G_2_15_port, Pij => P_2_15_port)
                           ;
   PG_BLOCK_REG_INSTANCE_2_19 : PG_BLOCK_15 port map( Gik => G_1_19_port, Gkj 
                           => G_1_17_port, Pik => P_1_19_port, Pkj => 
                           P_1_17_port, Gij => G_3_19_port, Pij => P_3_19_port)
                           ;
   PG_BLOCK_REG_INSTANCE_2_23 : PG_BLOCK_14 port map( Gik => G_1_23_port, Gkj 
                           => G_1_21_port, Pik => P_1_23_port, Pkj => 
                           P_1_21_port, Gij => G_2_23_port, Pij => P_2_23_port)
                           ;
   PG_BLOCK_REG_INSTANCE_2_27 : PG_BLOCK_13 port map( Gik => G_1_27_port, Gkj 
                           => G_1_25_port, Pik => P_1_27_port, Pkj => 
                           P_1_25_port, Gij => G_3_27_port, Pij => P_3_27_port)
                           ;
   PG_BLOCK_REG_INSTANCE_2_31 : PG_BLOCK_12 port map( Gik => G_1_31_port, Gkj 
                           => G_1_29_port, Pik => P_1_31_port, Pkj => 
                           P_1_29_port, Gij => G_2_31_port, Pij => P_2_31_port)
                           ;
   G_BLOCK_INSTANCE_3_7 : GENERATE_BLOCK_6 port map( Gik => G_2_7_port, Gkj => 
                           Co_0_port, Pik => P_2_7_port, Gij => n1);
   PG_BLOCK_REG_INSTANCE_3_7 : PG_BLOCK_11 port map( Gik => G_2_7_port, Gkj => 
                           Co_0_port, Pik => P_2_7_port, Pkj => X_Logic0_port, 
                           Gij => n2, Pij => P_4_7_port);
   PG_BLOCK_REG_INSTANCE_3_15 : PG_BLOCK_10 port map( Gik => G_2_15_port, Gkj 
                           => G_3_11_port, Pik => P_2_15_port, Pkj => 
                           P_3_11_port, Gij => G_3_15_port, Pij => P_3_15_port)
                           ;
   PG_BLOCK_REG_INSTANCE_3_23 : PG_BLOCK_9 port map( Gik => G_2_23_port, Gkj =>
                           G_3_19_port, Pik => P_2_23_port, Pkj => P_3_19_port,
                           Gij => G_4_23_port, Pij => P_4_23_port);
   PG_BLOCK_REG_INSTANCE_3_31 : PG_BLOCK_8 port map( Gik => G_2_31_port, Gkj =>
                           G_3_27_port, Pik => P_2_31_port, Pkj => P_3_27_port,
                           Gij => G_3_31_port, Pij => P_3_31_port);
   G_BLOCK_INSTANCE_4_11 : GENERATE_BLOCK_5 port map( Gik => G_3_11_port, Gkj 
                           => Co_1_port, Pik => P_3_11_port, Gij => n3);
   PG_BLOCK_REG_INSTANCE_4_11 : PG_BLOCK_7 port map( Gik => G_3_11_port, Gkj =>
                           Co_1_port, Pik => P_3_11_port, Pkj => P_4_7_port, 
                           Gij => n4, Pij => n_1256);
   G_BLOCK_INSTANCE_4_15 : GENERATE_BLOCK_4 port map( Gik => G_3_15_port, Gkj 
                           => Co_1_port, Pik => P_3_15_port, Gij => n5);
   PG_BLOCK_REG_INSTANCE_4_15 : PG_BLOCK_6 port map( Gik => G_3_15_port, Gkj =>
                           Co_1_port, Pik => P_3_15_port, Pkj => P_4_7_port, 
                           Gij => n6, Pij => P_5_15_port);
   PG_BLOCK_REG_INSTANCE_4_27 : PG_BLOCK_5 port map( Gik => G_3_27_port, Gkj =>
                           G_4_23_port, Pik => P_3_27_port, Pkj => P_4_23_port,
                           Gij => G_4_27_port, Pij => P_4_27_port);
   PG_BLOCK_REG_INSTANCE_4_31 : PG_BLOCK_4 port map( Gik => G_3_31_port, Gkj =>
                           G_4_23_port, Pik => P_3_31_port, Pkj => P_4_23_port,
                           Gij => G_4_31_port, Pij => P_4_31_port);
   G_BLOCK_INSTANCE_5_19 : GENERATE_BLOCK_3 port map( Gik => G_3_19_port, Gkj 
                           => Co_3_port, Pik => P_3_19_port, Gij => n7);
   PG_BLOCK_REG_INSTANCE_5_19 : PG_BLOCK_3 port map( Gik => G_3_19_port, Gkj =>
                           Co_3_port, Pik => P_3_19_port, Pkj => P_5_15_port, 
                           Gij => n8, Pij => n_1257);
   G_BLOCK_INSTANCE_5_23 : GENERATE_BLOCK_2 port map( Gik => G_4_23_port, Gkj 
                           => Co_3_port, Pik => P_4_23_port, Gij => n9);
   PG_BLOCK_REG_INSTANCE_5_23 : PG_BLOCK_2 port map( Gik => G_4_23_port, Gkj =>
                           Co_3_port, Pik => P_4_23_port, Pkj => P_5_15_port, 
                           Gij => n10, Pij => n_1258);
   G_BLOCK_INSTANCE_5_27 : GENERATE_BLOCK_1 port map( Gik => G_4_27_port, Gkj 
                           => Co_3_port, Pik => P_4_27_port, Gij => n11);
   PG_BLOCK_REG_INSTANCE_5_27 : PG_BLOCK_1 port map( Gik => G_4_27_port, Gkj =>
                           Co_3_port, Pik => P_4_27_port, Pkj => P_5_15_port, 
                           Gij => n12, Pij => n_1259);
   G_BLOCK_INSTANCE_5_31 : GENERATE_BLOCK_0 port map( Gik => G_4_31_port, Gkj 
                           => Co_3_port, Pik => P_4_31_port, Gij => n13);
   PG_BLOCK_REG_INSTANCE_5_31 : PG_BLOCK_0 port map( Gik => G_4_31_port, Gkj =>
                           Co_3_port, Pik => P_4_31_port, Pkj => P_5_15_port, 
                           Gij => n14, Pij => n_1260);
   U2 : AND2_X1 port map( A1 => n14, A2 => n13, ZN => Co_7_port);
   U3 : AND2_X1 port map( A1 => n12, A2 => n11, ZN => Co_6_port);
   U4 : AND2_X1 port map( A1 => n10, A2 => n9, ZN => Co_5_port);
   U5 : AND2_X1 port map( A1 => n8, A2 => n7, ZN => Co_4_port);
   U6 : AND2_X1 port map( A1 => n6, A2 => n5, ZN => Co_3_port);
   U7 : AND2_X1 port map( A1 => n4, A2 => n3, ZN => Co_2_port);
   U8 : AND2_X1 port map( A1 => n2, A2 => n1, ZN => Co_1_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end AND2_61;

architecture SYN_BEHAVIORAL of AND2_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity XNOR2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end XNOR2_63;

architecture SYN_BEHAVIORAL of XNOR2_63 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ZERO_DETECTOR_N32_0 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic);

end ZERO_DETECTOR_N32_0;

architecture SYN_STRUCTURAL of ZERO_DETECTOR_N32_0 is

   component AND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, M_4_1_port, M_4_0_port, M_3_3_port, M_3_2_port, 
      M_3_1_port, M_3_0_port, M_2_7_port, M_2_6_port, M_2_5_port, M_2_4_port, 
      M_2_3_port, M_2_2_port, M_2_1_port, M_2_0_port, M_1_15_port, M_1_14_port,
      M_1_13_port, M_1_12_port, M_1_11_port, M_1_10_port, M_1_9_port, 
      M_1_8_port, M_1_7_port, M_1_6_port, M_1_5_port, M_1_4_port, M_1_3_port, 
      M_1_2_port, M_1_1_port, M_1_0_port, M_0_31_port, M_0_30_port, M_0_29_port
      , M_0_28_port, M_0_27_port, M_0_26_port, M_0_25_port, M_0_24_port, 
      M_0_23_port, M_0_22_port, M_0_21_port, M_0_20_port, M_0_19_port, 
      M_0_18_port, M_0_17_port, M_0_16_port, M_0_15_port, M_0_14_port, 
      M_0_13_port, M_0_12_port, M_0_11_port, M_0_10_port, M_0_9_port, 
      M_0_8_port, M_0_7_port, M_0_6_port, M_0_5_port, M_0_4_port, M_0_3_port, 
      M_0_2_port, M_0_1_port, M_0_0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   XOR0_i_0_0 : XNOR2_31 port map( A => A(0), B => X_Logic0_port, Y => 
                           M_0_0_port);
   XOR0_i_0_1 : XNOR2_30 port map( A => A(1), B => X_Logic0_port, Y => 
                           M_0_1_port);
   XOR0_i_0_2 : XNOR2_29 port map( A => A(2), B => X_Logic0_port, Y => 
                           M_0_2_port);
   XOR0_i_0_3 : XNOR2_28 port map( A => A(3), B => X_Logic0_port, Y => 
                           M_0_3_port);
   XOR0_i_0_4 : XNOR2_27 port map( A => A(4), B => X_Logic0_port, Y => 
                           M_0_4_port);
   XOR0_i_0_5 : XNOR2_26 port map( A => A(5), B => X_Logic0_port, Y => 
                           M_0_5_port);
   XOR0_i_0_6 : XNOR2_25 port map( A => A(6), B => X_Logic0_port, Y => 
                           M_0_6_port);
   XOR0_i_0_7 : XNOR2_24 port map( A => A(7), B => X_Logic0_port, Y => 
                           M_0_7_port);
   XOR0_i_0_8 : XNOR2_23 port map( A => A(8), B => X_Logic0_port, Y => 
                           M_0_8_port);
   XOR0_i_0_9 : XNOR2_22 port map( A => A(9), B => X_Logic0_port, Y => 
                           M_0_9_port);
   XOR0_i_0_10 : XNOR2_21 port map( A => A(10), B => X_Logic0_port, Y => 
                           M_0_10_port);
   XOR0_i_0_11 : XNOR2_20 port map( A => A(11), B => X_Logic0_port, Y => 
                           M_0_11_port);
   XOR0_i_0_12 : XNOR2_19 port map( A => A(12), B => X_Logic0_port, Y => 
                           M_0_12_port);
   XOR0_i_0_13 : XNOR2_18 port map( A => A(13), B => X_Logic0_port, Y => 
                           M_0_13_port);
   XOR0_i_0_14 : XNOR2_17 port map( A => A(14), B => X_Logic0_port, Y => 
                           M_0_14_port);
   XOR0_i_0_15 : XNOR2_16 port map( A => A(15), B => X_Logic0_port, Y => 
                           M_0_15_port);
   XOR0_i_0_16 : XNOR2_15 port map( A => A(16), B => X_Logic0_port, Y => 
                           M_0_16_port);
   XOR0_i_0_17 : XNOR2_14 port map( A => A(17), B => X_Logic0_port, Y => 
                           M_0_17_port);
   XOR0_i_0_18 : XNOR2_13 port map( A => A(18), B => X_Logic0_port, Y => 
                           M_0_18_port);
   XOR0_i_0_19 : XNOR2_12 port map( A => A(19), B => X_Logic0_port, Y => 
                           M_0_19_port);
   XOR0_i_0_20 : XNOR2_11 port map( A => A(20), B => X_Logic0_port, Y => 
                           M_0_20_port);
   XOR0_i_0_21 : XNOR2_10 port map( A => A(21), B => X_Logic0_port, Y => 
                           M_0_21_port);
   XOR0_i_0_22 : XNOR2_9 port map( A => A(22), B => X_Logic0_port, Y => 
                           M_0_22_port);
   XOR0_i_0_23 : XNOR2_8 port map( A => A(23), B => X_Logic0_port, Y => 
                           M_0_23_port);
   XOR0_i_0_24 : XNOR2_7 port map( A => A(24), B => X_Logic0_port, Y => 
                           M_0_24_port);
   XOR0_i_0_25 : XNOR2_6 port map( A => A(25), B => X_Logic0_port, Y => 
                           M_0_25_port);
   XOR0_i_0_26 : XNOR2_5 port map( A => A(26), B => X_Logic0_port, Y => 
                           M_0_26_port);
   XOR0_i_0_27 : XNOR2_4 port map( A => A(27), B => X_Logic0_port, Y => 
                           M_0_27_port);
   XOR0_i_0_28 : XNOR2_3 port map( A => A(28), B => X_Logic0_port, Y => 
                           M_0_28_port);
   XOR0_i_0_29 : XNOR2_2 port map( A => A(29), B => X_Logic0_port, Y => 
                           M_0_29_port);
   XOR0_i_0_30 : XNOR2_1 port map( A => A(30), B => X_Logic0_port, Y => 
                           M_0_30_port);
   XOR0_i_0_31 : XNOR2_0 port map( A => A(31), B => X_Logic0_port, Y => 
                           M_0_31_port);
   AND_i_1_0 : AND2_30 port map( A => M_0_0_port, B => M_0_1_port, Y => 
                           M_1_0_port);
   AND_i_1_1 : AND2_29 port map( A => M_0_2_port, B => M_0_3_port, Y => 
                           M_1_1_port);
   AND_i_1_2 : AND2_28 port map( A => M_0_4_port, B => M_0_5_port, Y => 
                           M_1_2_port);
   AND_i_1_3 : AND2_27 port map( A => M_0_6_port, B => M_0_7_port, Y => 
                           M_1_3_port);
   AND_i_1_4 : AND2_26 port map( A => M_0_8_port, B => M_0_9_port, Y => 
                           M_1_4_port);
   AND_i_1_5 : AND2_25 port map( A => M_0_10_port, B => M_0_11_port, Y => 
                           M_1_5_port);
   AND_i_1_6 : AND2_24 port map( A => M_0_12_port, B => M_0_13_port, Y => 
                           M_1_6_port);
   AND_i_1_7 : AND2_23 port map( A => M_0_14_port, B => M_0_15_port, Y => 
                           M_1_7_port);
   AND_i_1_8 : AND2_22 port map( A => M_0_16_port, B => M_0_17_port, Y => 
                           M_1_8_port);
   AND_i_1_9 : AND2_21 port map( A => M_0_18_port, B => M_0_19_port, Y => 
                           M_1_9_port);
   AND_i_1_10 : AND2_20 port map( A => M_0_20_port, B => M_0_21_port, Y => 
                           M_1_10_port);
   AND_i_1_11 : AND2_19 port map( A => M_0_22_port, B => M_0_23_port, Y => 
                           M_1_11_port);
   AND_i_1_12 : AND2_18 port map( A => M_0_24_port, B => M_0_25_port, Y => 
                           M_1_12_port);
   AND_i_1_13 : AND2_17 port map( A => M_0_26_port, B => M_0_27_port, Y => 
                           M_1_13_port);
   AND_i_1_14 : AND2_16 port map( A => M_0_28_port, B => M_0_29_port, Y => 
                           M_1_14_port);
   AND_i_1_15 : AND2_15 port map( A => M_0_30_port, B => M_0_31_port, Y => 
                           M_1_15_port);
   AND_i_2_0 : AND2_14 port map( A => M_1_0_port, B => M_1_1_port, Y => 
                           M_2_0_port);
   AND_i_2_1 : AND2_13 port map( A => M_1_2_port, B => M_1_3_port, Y => 
                           M_2_1_port);
   AND_i_2_2 : AND2_12 port map( A => M_1_4_port, B => M_1_5_port, Y => 
                           M_2_2_port);
   AND_i_2_3 : AND2_11 port map( A => M_1_6_port, B => M_1_7_port, Y => 
                           M_2_3_port);
   AND_i_2_4 : AND2_10 port map( A => M_1_8_port, B => M_1_9_port, Y => 
                           M_2_4_port);
   AND_i_2_5 : AND2_9 port map( A => M_1_10_port, B => M_1_11_port, Y => 
                           M_2_5_port);
   AND_i_2_6 : AND2_8 port map( A => M_1_12_port, B => M_1_13_port, Y => 
                           M_2_6_port);
   AND_i_2_7 : AND2_7 port map( A => M_1_14_port, B => M_1_15_port, Y => 
                           M_2_7_port);
   AND_i_3_0 : AND2_6 port map( A => M_2_0_port, B => M_2_1_port, Y => 
                           M_3_0_port);
   AND_i_3_1 : AND2_5 port map( A => M_2_2_port, B => M_2_3_port, Y => 
                           M_3_1_port);
   AND_i_3_2 : AND2_4 port map( A => M_2_4_port, B => M_2_5_port, Y => 
                           M_3_2_port);
   AND_i_3_3 : AND2_3 port map( A => M_2_6_port, B => M_2_7_port, Y => 
                           M_3_3_port);
   AND_i_4_0 : AND2_2 port map( A => M_3_0_port, B => M_3_1_port, Y => 
                           M_4_0_port);
   AND_i_4_1 : AND2_1 port map( A => M_3_2_port, B => M_3_3_port, Y => 
                           M_4_1_port);
   AND_i_5_0 : AND2_0 port map( A => M_4_0_port, B => M_4_1_port, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity COMPARATOR_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic_vector (3 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end COMPARATOR_N32;

architecture SYN_BEHAVIORAL of COMPARATOR_N32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal X_Logic0_port, Y_0_port, N46, N48, N49, N50, N51, n17, n18, n1, n2, 
      n3, n4, n5, n6, n7, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, 
      n_1267 : std_logic;

begin
   Y <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, Y_0_port );
   
   X_Logic0_port <= '0';
   n17 <= '1';
   n18 <= '0';
   r91 : COMPARATOR_N32_DW01_cmp6_0_DW01_cmp6_4 port map( A(31) => A(31), A(30)
                           => A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), TC => n17, LT => N48, GT => 
                           N50, EQ => n_1261, LE => n_1262, GE => n_1263, NE =>
                           n_1264);
   r90 : COMPARATOR_N32_DW01_cmp6_1_DW01_cmp6_5 port map( A(31) => A(31), A(30)
                           => A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), TC => n18, LT => N49, GT => 
                           N51, EQ => N46, LE => n_1265, GE => n_1266, NE => 
                           n_1267);
   U4 : MUX2_X1 port map( A => n1, B => n2, S => S(3), Z => Y_0_port);
   U5 : NOR3_X1 port map( A1 => n3, A2 => S(2), A3 => S(1), ZN => n2);
   U6 : MUX2_X1 port map( A => n4, B => n5, S => S(2), Z => n1);
   U7 : XOR2_X1 port map( A => S(1), B => n6, Z => n5);
   U8 : MUX2_X1 port map( A => N50, B => N51, S => S(0), Z => n6);
   U9 : MUX2_X1 port map( A => n7, B => n3, S => S(1), Z => n4);
   U10 : MUX2_X1 port map( A => N48, B => N49, S => S(0), Z => n3);
   U11 : XOR2_X1 port map( A => N46, B => S(0), Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LOGIC_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic_vector (1 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end LOGIC_N32;

architecture SYN_BEHAVIORAL of LOGIC_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164 : std_logic;

begin
   
   U2 : OR2_X1 port map( A1 => n8, A2 => S(0), ZN => n1);
   U3 : AND2_X4 port map( A1 => S(0), A2 => n8, ZN => n6);
   U4 : INV_X4 port map( A => n1, ZN => n2);
   U5 : INV_X2 port map( A => S(1), ZN => n8);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n4, A => n5, ZN => Y(9));
   U7 : OAI21_X1 port map( B1 => n6, B2 => n7, A => B(9), ZN => n5);
   U8 : MUX2_X1 port map( A => n8, B => n2, S => n4, Z => n7);
   U9 : INV_X1 port map( A => A(9), ZN => n4);
   U10 : AOI21_X1 port map( B1 => n2, B2 => n9, A => n6, ZN => n3);
   U11 : INV_X1 port map( A => B(9), ZN => n9);
   U12 : OAI21_X1 port map( B1 => n10, B2 => n11, A => n12, ZN => Y(8));
   U13 : OAI21_X1 port map( B1 => n6, B2 => n13, A => B(8), ZN => n12);
   U14 : MUX2_X1 port map( A => n8, B => n2, S => n11, Z => n13);
   U15 : INV_X1 port map( A => A(8), ZN => n11);
   U16 : AOI21_X1 port map( B1 => n2, B2 => n14, A => n6, ZN => n10);
   U17 : INV_X1 port map( A => B(8), ZN => n14);
   U18 : OAI21_X1 port map( B1 => n15, B2 => n16, A => n17, ZN => Y(7));
   U19 : OAI21_X1 port map( B1 => n6, B2 => n18, A => B(7), ZN => n17);
   U20 : MUX2_X1 port map( A => n8, B => n2, S => n16, Z => n18);
   U21 : INV_X1 port map( A => A(7), ZN => n16);
   U22 : AOI21_X1 port map( B1 => n2, B2 => n19, A => n6, ZN => n15);
   U23 : INV_X1 port map( A => B(7), ZN => n19);
   U24 : OAI21_X1 port map( B1 => n20, B2 => n21, A => n22, ZN => Y(6));
   U25 : OAI21_X1 port map( B1 => n6, B2 => n23, A => B(6), ZN => n22);
   U26 : MUX2_X1 port map( A => n8, B => n2, S => n21, Z => n23);
   U27 : INV_X1 port map( A => A(6), ZN => n21);
   U28 : AOI21_X1 port map( B1 => n2, B2 => n24, A => n6, ZN => n20);
   U29 : INV_X1 port map( A => B(6), ZN => n24);
   U30 : OAI21_X1 port map( B1 => n25, B2 => n26, A => n27, ZN => Y(5));
   U31 : OAI21_X1 port map( B1 => n6, B2 => n28, A => B(5), ZN => n27);
   U32 : MUX2_X1 port map( A => n8, B => n2, S => n26, Z => n28);
   U33 : INV_X1 port map( A => A(5), ZN => n26);
   U34 : AOI21_X1 port map( B1 => n2, B2 => n29, A => n6, ZN => n25);
   U35 : INV_X1 port map( A => B(5), ZN => n29);
   U36 : OAI21_X1 port map( B1 => n30, B2 => n31, A => n32, ZN => Y(4));
   U37 : OAI21_X1 port map( B1 => n6, B2 => n33, A => B(4), ZN => n32);
   U38 : MUX2_X1 port map( A => n8, B => n2, S => n31, Z => n33);
   U39 : INV_X1 port map( A => A(4), ZN => n31);
   U40 : AOI21_X1 port map( B1 => n2, B2 => n34, A => n6, ZN => n30);
   U41 : INV_X1 port map( A => B(4), ZN => n34);
   U42 : OAI21_X1 port map( B1 => n35, B2 => n36, A => n37, ZN => Y(3));
   U43 : OAI21_X1 port map( B1 => n6, B2 => n38, A => B(3), ZN => n37);
   U44 : MUX2_X1 port map( A => n8, B => n2, S => n36, Z => n38);
   U45 : INV_X1 port map( A => A(3), ZN => n36);
   U46 : AOI21_X1 port map( B1 => n2, B2 => n39, A => n6, ZN => n35);
   U47 : INV_X1 port map( A => B(3), ZN => n39);
   U48 : OAI21_X1 port map( B1 => n40, B2 => n41, A => n42, ZN => Y(31));
   U49 : OAI21_X1 port map( B1 => n6, B2 => n43, A => B(31), ZN => n42);
   U50 : MUX2_X1 port map( A => n8, B => n2, S => n41, Z => n43);
   U51 : INV_X1 port map( A => A(31), ZN => n41);
   U52 : AOI21_X1 port map( B1 => n2, B2 => n44, A => n6, ZN => n40);
   U53 : INV_X1 port map( A => B(31), ZN => n44);
   U54 : OAI21_X1 port map( B1 => n45, B2 => n46, A => n47, ZN => Y(30));
   U55 : OAI21_X1 port map( B1 => n6, B2 => n48, A => B(30), ZN => n47);
   U56 : MUX2_X1 port map( A => n8, B => n2, S => n46, Z => n48);
   U57 : INV_X1 port map( A => A(30), ZN => n46);
   U58 : AOI21_X1 port map( B1 => n2, B2 => n49, A => n6, ZN => n45);
   U59 : INV_X1 port map( A => B(30), ZN => n49);
   U60 : OAI21_X1 port map( B1 => n50, B2 => n51, A => n52, ZN => Y(2));
   U61 : OAI21_X1 port map( B1 => n6, B2 => n53, A => B(2), ZN => n52);
   U62 : MUX2_X1 port map( A => n8, B => n2, S => n51, Z => n53);
   U63 : INV_X1 port map( A => A(2), ZN => n51);
   U64 : AOI21_X1 port map( B1 => n2, B2 => n54, A => n6, ZN => n50);
   U65 : INV_X1 port map( A => B(2), ZN => n54);
   U66 : OAI21_X1 port map( B1 => n55, B2 => n56, A => n57, ZN => Y(29));
   U67 : OAI21_X1 port map( B1 => n6, B2 => n58, A => B(29), ZN => n57);
   U68 : MUX2_X1 port map( A => n8, B => n2, S => n56, Z => n58);
   U69 : INV_X1 port map( A => A(29), ZN => n56);
   U70 : AOI21_X1 port map( B1 => n2, B2 => n59, A => n6, ZN => n55);
   U71 : INV_X1 port map( A => B(29), ZN => n59);
   U72 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => Y(28));
   U73 : OAI21_X1 port map( B1 => n6, B2 => n63, A => B(28), ZN => n62);
   U74 : MUX2_X1 port map( A => n8, B => n2, S => n61, Z => n63);
   U75 : INV_X1 port map( A => A(28), ZN => n61);
   U76 : AOI21_X1 port map( B1 => n2, B2 => n64, A => n6, ZN => n60);
   U77 : INV_X1 port map( A => B(28), ZN => n64);
   U78 : OAI21_X1 port map( B1 => n65, B2 => n66, A => n67, ZN => Y(27));
   U79 : OAI21_X1 port map( B1 => n6, B2 => n68, A => B(27), ZN => n67);
   U80 : MUX2_X1 port map( A => n8, B => n2, S => n66, Z => n68);
   U81 : INV_X1 port map( A => A(27), ZN => n66);
   U82 : AOI21_X1 port map( B1 => n2, B2 => n69, A => n6, ZN => n65);
   U83 : INV_X1 port map( A => B(27), ZN => n69);
   U84 : OAI21_X1 port map( B1 => n70, B2 => n71, A => n72, ZN => Y(26));
   U85 : OAI21_X1 port map( B1 => n6, B2 => n73, A => B(26), ZN => n72);
   U86 : MUX2_X1 port map( A => n8, B => n2, S => n71, Z => n73);
   U87 : INV_X1 port map( A => A(26), ZN => n71);
   U88 : AOI21_X1 port map( B1 => n2, B2 => n74, A => n6, ZN => n70);
   U89 : INV_X1 port map( A => B(26), ZN => n74);
   U90 : OAI21_X1 port map( B1 => n75, B2 => n76, A => n77, ZN => Y(25));
   U91 : OAI21_X1 port map( B1 => n6, B2 => n78, A => B(25), ZN => n77);
   U92 : MUX2_X1 port map( A => n8, B => n2, S => n76, Z => n78);
   U93 : INV_X1 port map( A => A(25), ZN => n76);
   U94 : AOI21_X1 port map( B1 => n2, B2 => n79, A => n6, ZN => n75);
   U95 : INV_X1 port map( A => B(25), ZN => n79);
   U96 : OAI21_X1 port map( B1 => n80, B2 => n81, A => n82, ZN => Y(24));
   U97 : OAI21_X1 port map( B1 => n6, B2 => n83, A => B(24), ZN => n82);
   U98 : MUX2_X1 port map( A => n8, B => n2, S => n81, Z => n83);
   U99 : INV_X1 port map( A => A(24), ZN => n81);
   U100 : AOI21_X1 port map( B1 => n2, B2 => n84, A => n6, ZN => n80);
   U101 : INV_X1 port map( A => B(24), ZN => n84);
   U102 : OAI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => Y(23));
   U103 : OAI21_X1 port map( B1 => n6, B2 => n88, A => B(23), ZN => n87);
   U104 : MUX2_X1 port map( A => n8, B => n2, S => n86, Z => n88);
   U105 : INV_X1 port map( A => A(23), ZN => n86);
   U106 : AOI21_X1 port map( B1 => n2, B2 => n89, A => n6, ZN => n85);
   U107 : INV_X1 port map( A => B(23), ZN => n89);
   U108 : OAI21_X1 port map( B1 => n90, B2 => n91, A => n92, ZN => Y(22));
   U109 : OAI21_X1 port map( B1 => n6, B2 => n93, A => B(22), ZN => n92);
   U110 : MUX2_X1 port map( A => n8, B => n2, S => n91, Z => n93);
   U111 : INV_X1 port map( A => A(22), ZN => n91);
   U112 : AOI21_X1 port map( B1 => n2, B2 => n94, A => n6, ZN => n90);
   U113 : INV_X1 port map( A => B(22), ZN => n94);
   U114 : OAI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => Y(21));
   U115 : OAI21_X1 port map( B1 => n6, B2 => n98, A => B(21), ZN => n97);
   U116 : MUX2_X1 port map( A => n8, B => n2, S => n96, Z => n98);
   U117 : INV_X1 port map( A => A(21), ZN => n96);
   U118 : AOI21_X1 port map( B1 => n2, B2 => n99, A => n6, ZN => n95);
   U119 : INV_X1 port map( A => B(21), ZN => n99);
   U120 : OAI21_X1 port map( B1 => n100, B2 => n101, A => n102, ZN => Y(20));
   U121 : OAI21_X1 port map( B1 => n6, B2 => n103, A => B(20), ZN => n102);
   U122 : MUX2_X1 port map( A => n8, B => n2, S => n101, Z => n103);
   U123 : INV_X1 port map( A => A(20), ZN => n101);
   U124 : AOI21_X1 port map( B1 => n2, B2 => n104, A => n6, ZN => n100);
   U125 : INV_X1 port map( A => B(20), ZN => n104);
   U126 : OAI21_X1 port map( B1 => n105, B2 => n106, A => n107, ZN => Y(1));
   U127 : OAI21_X1 port map( B1 => n6, B2 => n108, A => B(1), ZN => n107);
   U128 : MUX2_X1 port map( A => n8, B => n2, S => n106, Z => n108);
   U129 : INV_X1 port map( A => A(1), ZN => n106);
   U130 : AOI21_X1 port map( B1 => n2, B2 => n109, A => n6, ZN => n105);
   U131 : INV_X1 port map( A => B(1), ZN => n109);
   U132 : OAI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => Y(19));
   U133 : OAI21_X1 port map( B1 => n6, B2 => n113, A => B(19), ZN => n112);
   U134 : MUX2_X1 port map( A => n8, B => n2, S => n111, Z => n113);
   U135 : INV_X1 port map( A => A(19), ZN => n111);
   U136 : AOI21_X1 port map( B1 => n2, B2 => n114, A => n6, ZN => n110);
   U137 : INV_X1 port map( A => B(19), ZN => n114);
   U138 : OAI21_X1 port map( B1 => n115, B2 => n116, A => n117, ZN => Y(18));
   U139 : OAI21_X1 port map( B1 => n6, B2 => n118, A => B(18), ZN => n117);
   U140 : MUX2_X1 port map( A => n8, B => n2, S => n116, Z => n118);
   U141 : INV_X1 port map( A => A(18), ZN => n116);
   U142 : AOI21_X1 port map( B1 => n2, B2 => n119, A => n6, ZN => n115);
   U143 : INV_X1 port map( A => B(18), ZN => n119);
   U144 : OAI21_X1 port map( B1 => n120, B2 => n121, A => n122, ZN => Y(17));
   U145 : OAI21_X1 port map( B1 => n6, B2 => n123, A => B(17), ZN => n122);
   U146 : MUX2_X1 port map( A => n8, B => n2, S => n121, Z => n123);
   U147 : INV_X1 port map( A => A(17), ZN => n121);
   U148 : AOI21_X1 port map( B1 => n2, B2 => n124, A => n6, ZN => n120);
   U149 : INV_X1 port map( A => B(17), ZN => n124);
   U150 : OAI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => Y(16));
   U151 : OAI21_X1 port map( B1 => n6, B2 => n128, A => B(16), ZN => n127);
   U152 : MUX2_X1 port map( A => n8, B => n2, S => n126, Z => n128);
   U153 : INV_X1 port map( A => A(16), ZN => n126);
   U154 : AOI21_X1 port map( B1 => n2, B2 => n129, A => n6, ZN => n125);
   U155 : INV_X1 port map( A => B(16), ZN => n129);
   U156 : OAI21_X1 port map( B1 => n130, B2 => n131, A => n132, ZN => Y(15));
   U157 : OAI21_X1 port map( B1 => n6, B2 => n133, A => B(15), ZN => n132);
   U158 : MUX2_X1 port map( A => n8, B => n2, S => n131, Z => n133);
   U159 : INV_X1 port map( A => A(15), ZN => n131);
   U160 : AOI21_X1 port map( B1 => n2, B2 => n134, A => n6, ZN => n130);
   U161 : INV_X1 port map( A => B(15), ZN => n134);
   U162 : OAI21_X1 port map( B1 => n135, B2 => n136, A => n137, ZN => Y(14));
   U163 : OAI21_X1 port map( B1 => n6, B2 => n138, A => B(14), ZN => n137);
   U164 : MUX2_X1 port map( A => n8, B => n2, S => n136, Z => n138);
   U165 : INV_X1 port map( A => A(14), ZN => n136);
   U166 : AOI21_X1 port map( B1 => n2, B2 => n139, A => n6, ZN => n135);
   U167 : INV_X1 port map( A => B(14), ZN => n139);
   U168 : OAI21_X1 port map( B1 => n140, B2 => n141, A => n142, ZN => Y(13));
   U169 : OAI21_X1 port map( B1 => n6, B2 => n143, A => B(13), ZN => n142);
   U170 : MUX2_X1 port map( A => n8, B => n2, S => n141, Z => n143);
   U171 : INV_X1 port map( A => A(13), ZN => n141);
   U172 : AOI21_X1 port map( B1 => n2, B2 => n144, A => n6, ZN => n140);
   U173 : INV_X1 port map( A => B(13), ZN => n144);
   U174 : OAI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => Y(12));
   U175 : OAI21_X1 port map( B1 => n6, B2 => n148, A => B(12), ZN => n147);
   U176 : MUX2_X1 port map( A => n8, B => n2, S => n146, Z => n148);
   U177 : INV_X1 port map( A => A(12), ZN => n146);
   U178 : AOI21_X1 port map( B1 => n2, B2 => n149, A => n6, ZN => n145);
   U179 : INV_X1 port map( A => B(12), ZN => n149);
   U180 : OAI21_X1 port map( B1 => n150, B2 => n151, A => n152, ZN => Y(11));
   U181 : OAI21_X1 port map( B1 => n6, B2 => n153, A => B(11), ZN => n152);
   U182 : MUX2_X1 port map( A => n8, B => n2, S => n151, Z => n153);
   U183 : INV_X1 port map( A => A(11), ZN => n151);
   U184 : AOI21_X1 port map( B1 => n2, B2 => n154, A => n6, ZN => n150);
   U185 : INV_X1 port map( A => B(11), ZN => n154);
   U186 : OAI21_X1 port map( B1 => n155, B2 => n156, A => n157, ZN => Y(10));
   U187 : OAI21_X1 port map( B1 => n6, B2 => n158, A => B(10), ZN => n157);
   U188 : MUX2_X1 port map( A => n8, B => n2, S => n156, Z => n158);
   U189 : INV_X1 port map( A => A(10), ZN => n156);
   U190 : AOI21_X1 port map( B1 => n2, B2 => n159, A => n6, ZN => n155);
   U191 : INV_X1 port map( A => B(10), ZN => n159);
   U192 : OAI21_X1 port map( B1 => n160, B2 => n161, A => n162, ZN => Y(0));
   U193 : OAI21_X1 port map( B1 => n6, B2 => n163, A => B(0), ZN => n162);
   U194 : MUX2_X1 port map( A => n8, B => n2, S => n161, Z => n163);
   U195 : INV_X1 port map( A => A(0), ZN => n161);
   U196 : AOI21_X1 port map( B1 => n2, B2 => n164, A => n6, ZN => n160);
   U197 : INV_X1 port map( A => B(0), ZN => n164);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BARREL_SHIFTER_RIGHT_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end BARREL_SHIFTER_RIGHT_N32;

architecture SYN_STRUCTURAL of BARREL_SHIFTER_RIGHT_N32 is

   component MUX21_L_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_32
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_33
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_34
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_35
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_36
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_37
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_38
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_39
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_40
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_41
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_42
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_43
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_44
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_45
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_46
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_47
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_48
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_49
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_50
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_51
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_52
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_53
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_54
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_55
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_56
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_57
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_58
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_59
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_60
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_61
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_62
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_63
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_64
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_65
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_66
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_67
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_68
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_69
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_70
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_71
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_72
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_73
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_74
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_75
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_76
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_77
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_78
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_79
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_80
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_81
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_82
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_83
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_84
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_85
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_86
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_87
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_88
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_89
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_90
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_91
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_92
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_93
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_94
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_95
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_96
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_97
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_98
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_99
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_100
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_101
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_102
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_103
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_104
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_105
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_106
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_107
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_108
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_109
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_110
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_111
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_112
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_113
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_114
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_115
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_116
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_117
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_118
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_119
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_120
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_121
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_122
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_123
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_124
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_125
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_126
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_127
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_128
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_129
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_130
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_131
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_132
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_133
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_134
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_135
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_136
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_137
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_138
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_139
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_140
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_141
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_142
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_143
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_144
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_145
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_146
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_147
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_148
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_149
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_150
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_151
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_152
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_153
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_154
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_155
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_156
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_157
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_158
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_159
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal TMP_4_31_port, TMP_4_30_port, TMP_4_29_port, TMP_4_28_port, 
      TMP_4_27_port, TMP_4_26_port, TMP_4_25_port, TMP_4_24_port, TMP_4_23_port
      , TMP_4_22_port, TMP_4_21_port, TMP_4_20_port, TMP_4_19_port, 
      TMP_4_18_port, TMP_4_17_port, TMP_4_16_port, TMP_4_15_port, TMP_4_14_port
      , TMP_4_13_port, TMP_4_12_port, TMP_4_11_port, TMP_4_10_port, 
      TMP_4_9_port, TMP_4_8_port, TMP_4_7_port, TMP_4_6_port, TMP_4_5_port, 
      TMP_4_4_port, TMP_4_3_port, TMP_4_2_port, TMP_4_1_port, TMP_4_0_port, 
      TMP_3_31_port, TMP_3_30_port, TMP_3_29_port, TMP_3_28_port, TMP_3_27_port
      , TMP_3_26_port, TMP_3_25_port, TMP_3_24_port, TMP_3_23_port, 
      TMP_3_22_port, TMP_3_21_port, TMP_3_20_port, TMP_3_19_port, TMP_3_18_port
      , TMP_3_17_port, TMP_3_16_port, TMP_3_15_port, TMP_3_14_port, 
      TMP_3_13_port, TMP_3_12_port, TMP_3_11_port, TMP_3_10_port, TMP_3_9_port,
      TMP_3_8_port, TMP_3_7_port, TMP_3_6_port, TMP_3_5_port, TMP_3_4_port, 
      TMP_3_3_port, TMP_3_2_port, TMP_3_1_port, TMP_3_0_port, TMP_2_31_port, 
      TMP_2_30_port, TMP_2_29_port, TMP_2_28_port, TMP_2_27_port, TMP_2_26_port
      , TMP_2_25_port, TMP_2_24_port, TMP_2_23_port, TMP_2_22_port, 
      TMP_2_21_port, TMP_2_20_port, TMP_2_19_port, TMP_2_18_port, TMP_2_17_port
      , TMP_2_16_port, TMP_2_15_port, TMP_2_14_port, TMP_2_13_port, 
      TMP_2_12_port, TMP_2_11_port, TMP_2_10_port, TMP_2_9_port, TMP_2_8_port, 
      TMP_2_7_port, TMP_2_6_port, TMP_2_5_port, TMP_2_4_port, TMP_2_3_port, 
      TMP_2_2_port, TMP_2_1_port, TMP_2_0_port, TMP_1_31_port, TMP_1_30_port, 
      TMP_1_29_port, TMP_1_28_port, TMP_1_27_port, TMP_1_26_port, TMP_1_25_port
      , TMP_1_24_port, TMP_1_23_port, TMP_1_22_port, TMP_1_21_port, 
      TMP_1_20_port, TMP_1_19_port, TMP_1_18_port, TMP_1_17_port, TMP_1_16_port
      , TMP_1_15_port, TMP_1_14_port, TMP_1_13_port, TMP_1_12_port, 
      TMP_1_11_port, TMP_1_10_port, TMP_1_9_port, TMP_1_8_port, TMP_1_7_port, 
      TMP_1_6_port, TMP_1_5_port, TMP_1_4_port, TMP_1_3_port, TMP_1_2_port, 
      TMP_1_1_port, TMP_1_0_port : std_logic;

begin
   
   MUX21_K_0_0 : MUX21_L_159 port map( A => A(0), B => A(1), S => B(0), Y => 
                           TMP_1_0_port);
   MUX21_K_0_1 : MUX21_L_158 port map( A => A(1), B => A(2), S => B(0), Y => 
                           TMP_1_1_port);
   MUX21_K_0_2 : MUX21_L_157 port map( A => A(2), B => A(3), S => B(0), Y => 
                           TMP_1_2_port);
   MUX21_K_0_3 : MUX21_L_156 port map( A => A(3), B => A(4), S => B(0), Y => 
                           TMP_1_3_port);
   MUX21_K_0_4 : MUX21_L_155 port map( A => A(4), B => A(5), S => B(0), Y => 
                           TMP_1_4_port);
   MUX21_K_0_5 : MUX21_L_154 port map( A => A(5), B => A(6), S => B(0), Y => 
                           TMP_1_5_port);
   MUX21_K_0_6 : MUX21_L_153 port map( A => A(6), B => A(7), S => B(0), Y => 
                           TMP_1_6_port);
   MUX21_K_0_7 : MUX21_L_152 port map( A => A(7), B => A(8), S => B(0), Y => 
                           TMP_1_7_port);
   MUX21_K_0_8 : MUX21_L_151 port map( A => A(8), B => A(9), S => B(0), Y => 
                           TMP_1_8_port);
   MUX21_K_0_9 : MUX21_L_150 port map( A => A(9), B => A(10), S => B(0), Y => 
                           TMP_1_9_port);
   MUX21_K_0_10 : MUX21_L_149 port map( A => A(10), B => A(11), S => B(0), Y =>
                           TMP_1_10_port);
   MUX21_K_0_11 : MUX21_L_148 port map( A => A(11), B => A(12), S => B(0), Y =>
                           TMP_1_11_port);
   MUX21_K_0_12 : MUX21_L_147 port map( A => A(12), B => A(13), S => B(0), Y =>
                           TMP_1_12_port);
   MUX21_K_0_13 : MUX21_L_146 port map( A => A(13), B => A(14), S => B(0), Y =>
                           TMP_1_13_port);
   MUX21_K_0_14 : MUX21_L_145 port map( A => A(14), B => A(15), S => B(0), Y =>
                           TMP_1_14_port);
   MUX21_K_0_15 : MUX21_L_144 port map( A => A(15), B => A(16), S => B(0), Y =>
                           TMP_1_15_port);
   MUX21_K_0_16 : MUX21_L_143 port map( A => A(16), B => A(17), S => B(0), Y =>
                           TMP_1_16_port);
   MUX21_K_0_17 : MUX21_L_142 port map( A => A(17), B => A(18), S => B(0), Y =>
                           TMP_1_17_port);
   MUX21_K_0_18 : MUX21_L_141 port map( A => A(18), B => A(19), S => B(0), Y =>
                           TMP_1_18_port);
   MUX21_K_0_19 : MUX21_L_140 port map( A => A(19), B => A(20), S => B(0), Y =>
                           TMP_1_19_port);
   MUX21_K_0_20 : MUX21_L_139 port map( A => A(20), B => A(21), S => B(0), Y =>
                           TMP_1_20_port);
   MUX21_K_0_21 : MUX21_L_138 port map( A => A(21), B => A(22), S => B(0), Y =>
                           TMP_1_21_port);
   MUX21_K_0_22 : MUX21_L_137 port map( A => A(22), B => A(23), S => B(0), Y =>
                           TMP_1_22_port);
   MUX21_K_0_23 : MUX21_L_136 port map( A => A(23), B => A(24), S => B(0), Y =>
                           TMP_1_23_port);
   MUX21_K_0_24 : MUX21_L_135 port map( A => A(24), B => A(25), S => B(0), Y =>
                           TMP_1_24_port);
   MUX21_K_0_25 : MUX21_L_134 port map( A => A(25), B => A(26), S => B(0), Y =>
                           TMP_1_25_port);
   MUX21_K_0_26 : MUX21_L_133 port map( A => A(26), B => A(27), S => B(0), Y =>
                           TMP_1_26_port);
   MUX21_K_0_27 : MUX21_L_132 port map( A => A(27), B => A(28), S => B(0), Y =>
                           TMP_1_27_port);
   MUX21_K_0_28 : MUX21_L_131 port map( A => A(28), B => A(29), S => B(0), Y =>
                           TMP_1_28_port);
   MUX21_K_0_29 : MUX21_L_130 port map( A => A(29), B => A(30), S => B(0), Y =>
                           TMP_1_29_port);
   MUX21_K_0_30 : MUX21_L_129 port map( A => A(30), B => A(31), S => B(0), Y =>
                           TMP_1_30_port);
   MUX21_J_0_0 : MUX21_L_128 port map( A => A(31), B => S, S => B(0), Y => 
                           TMP_1_31_port);
   MUX21_K_1_0 : MUX21_L_127 port map( A => TMP_1_0_port, B => TMP_1_2_port, S 
                           => B(1), Y => TMP_2_0_port);
   MUX21_K_1_1 : MUX21_L_126 port map( A => TMP_1_1_port, B => TMP_1_3_port, S 
                           => B(1), Y => TMP_2_1_port);
   MUX21_K_1_2 : MUX21_L_125 port map( A => TMP_1_2_port, B => TMP_1_4_port, S 
                           => B(1), Y => TMP_2_2_port);
   MUX21_K_1_3 : MUX21_L_124 port map( A => TMP_1_3_port, B => TMP_1_5_port, S 
                           => B(1), Y => TMP_2_3_port);
   MUX21_K_1_4 : MUX21_L_123 port map( A => TMP_1_4_port, B => TMP_1_6_port, S 
                           => B(1), Y => TMP_2_4_port);
   MUX21_K_1_5 : MUX21_L_122 port map( A => TMP_1_5_port, B => TMP_1_7_port, S 
                           => B(1), Y => TMP_2_5_port);
   MUX21_K_1_6 : MUX21_L_121 port map( A => TMP_1_6_port, B => TMP_1_8_port, S 
                           => B(1), Y => TMP_2_6_port);
   MUX21_K_1_7 : MUX21_L_120 port map( A => TMP_1_7_port, B => TMP_1_9_port, S 
                           => B(1), Y => TMP_2_7_port);
   MUX21_K_1_8 : MUX21_L_119 port map( A => TMP_1_8_port, B => TMP_1_10_port, S
                           => B(1), Y => TMP_2_8_port);
   MUX21_K_1_9 : MUX21_L_118 port map( A => TMP_1_9_port, B => TMP_1_11_port, S
                           => B(1), Y => TMP_2_9_port);
   MUX21_K_1_10 : MUX21_L_117 port map( A => TMP_1_10_port, B => TMP_1_12_port,
                           S => B(1), Y => TMP_2_10_port);
   MUX21_K_1_11 : MUX21_L_116 port map( A => TMP_1_11_port, B => TMP_1_13_port,
                           S => B(1), Y => TMP_2_11_port);
   MUX21_K_1_12 : MUX21_L_115 port map( A => TMP_1_12_port, B => TMP_1_14_port,
                           S => B(1), Y => TMP_2_12_port);
   MUX21_K_1_13 : MUX21_L_114 port map( A => TMP_1_13_port, B => TMP_1_15_port,
                           S => B(1), Y => TMP_2_13_port);
   MUX21_K_1_14 : MUX21_L_113 port map( A => TMP_1_14_port, B => TMP_1_16_port,
                           S => B(1), Y => TMP_2_14_port);
   MUX21_K_1_15 : MUX21_L_112 port map( A => TMP_1_15_port, B => TMP_1_17_port,
                           S => B(1), Y => TMP_2_15_port);
   MUX21_K_1_16 : MUX21_L_111 port map( A => TMP_1_16_port, B => TMP_1_18_port,
                           S => B(1), Y => TMP_2_16_port);
   MUX21_K_1_17 : MUX21_L_110 port map( A => TMP_1_17_port, B => TMP_1_19_port,
                           S => B(1), Y => TMP_2_17_port);
   MUX21_K_1_18 : MUX21_L_109 port map( A => TMP_1_18_port, B => TMP_1_20_port,
                           S => B(1), Y => TMP_2_18_port);
   MUX21_K_1_19 : MUX21_L_108 port map( A => TMP_1_19_port, B => TMP_1_21_port,
                           S => B(1), Y => TMP_2_19_port);
   MUX21_K_1_20 : MUX21_L_107 port map( A => TMP_1_20_port, B => TMP_1_22_port,
                           S => B(1), Y => TMP_2_20_port);
   MUX21_K_1_21 : MUX21_L_106 port map( A => TMP_1_21_port, B => TMP_1_23_port,
                           S => B(1), Y => TMP_2_21_port);
   MUX21_K_1_22 : MUX21_L_105 port map( A => TMP_1_22_port, B => TMP_1_24_port,
                           S => B(1), Y => TMP_2_22_port);
   MUX21_K_1_23 : MUX21_L_104 port map( A => TMP_1_23_port, B => TMP_1_25_port,
                           S => B(1), Y => TMP_2_23_port);
   MUX21_K_1_24 : MUX21_L_103 port map( A => TMP_1_24_port, B => TMP_1_26_port,
                           S => B(1), Y => TMP_2_24_port);
   MUX21_K_1_25 : MUX21_L_102 port map( A => TMP_1_25_port, B => TMP_1_27_port,
                           S => B(1), Y => TMP_2_25_port);
   MUX21_K_1_26 : MUX21_L_101 port map( A => TMP_1_26_port, B => TMP_1_28_port,
                           S => B(1), Y => TMP_2_26_port);
   MUX21_K_1_27 : MUX21_L_100 port map( A => TMP_1_27_port, B => TMP_1_29_port,
                           S => B(1), Y => TMP_2_27_port);
   MUX21_K_1_28 : MUX21_L_99 port map( A => TMP_1_28_port, B => TMP_1_30_port, 
                           S => B(1), Y => TMP_2_28_port);
   MUX21_K_1_29 : MUX21_L_98 port map( A => TMP_1_29_port, B => TMP_1_31_port, 
                           S => B(1), Y => TMP_2_29_port);
   MUX21_J_1_0 : MUX21_L_97 port map( A => TMP_1_30_port, B => S, S => B(1), Y 
                           => TMP_2_30_port);
   MUX21_J_1_1 : MUX21_L_96 port map( A => TMP_1_31_port, B => S, S => B(1), Y 
                           => TMP_2_31_port);
   MUX21_K_2_0 : MUX21_L_95 port map( A => TMP_2_0_port, B => TMP_2_4_port, S 
                           => B(2), Y => TMP_3_0_port);
   MUX21_K_2_1 : MUX21_L_94 port map( A => TMP_2_1_port, B => TMP_2_5_port, S 
                           => B(2), Y => TMP_3_1_port);
   MUX21_K_2_2 : MUX21_L_93 port map( A => TMP_2_2_port, B => TMP_2_6_port, S 
                           => B(2), Y => TMP_3_2_port);
   MUX21_K_2_3 : MUX21_L_92 port map( A => TMP_2_3_port, B => TMP_2_7_port, S 
                           => B(2), Y => TMP_3_3_port);
   MUX21_K_2_4 : MUX21_L_91 port map( A => TMP_2_4_port, B => TMP_2_8_port, S 
                           => B(2), Y => TMP_3_4_port);
   MUX21_K_2_5 : MUX21_L_90 port map( A => TMP_2_5_port, B => TMP_2_9_port, S 
                           => B(2), Y => TMP_3_5_port);
   MUX21_K_2_6 : MUX21_L_89 port map( A => TMP_2_6_port, B => TMP_2_10_port, S 
                           => B(2), Y => TMP_3_6_port);
   MUX21_K_2_7 : MUX21_L_88 port map( A => TMP_2_7_port, B => TMP_2_11_port, S 
                           => B(2), Y => TMP_3_7_port);
   MUX21_K_2_8 : MUX21_L_87 port map( A => TMP_2_8_port, B => TMP_2_12_port, S 
                           => B(2), Y => TMP_3_8_port);
   MUX21_K_2_9 : MUX21_L_86 port map( A => TMP_2_9_port, B => TMP_2_13_port, S 
                           => B(2), Y => TMP_3_9_port);
   MUX21_K_2_10 : MUX21_L_85 port map( A => TMP_2_10_port, B => TMP_2_14_port, 
                           S => B(2), Y => TMP_3_10_port);
   MUX21_K_2_11 : MUX21_L_84 port map( A => TMP_2_11_port, B => TMP_2_15_port, 
                           S => B(2), Y => TMP_3_11_port);
   MUX21_K_2_12 : MUX21_L_83 port map( A => TMP_2_12_port, B => TMP_2_16_port, 
                           S => B(2), Y => TMP_3_12_port);
   MUX21_K_2_13 : MUX21_L_82 port map( A => TMP_2_13_port, B => TMP_2_17_port, 
                           S => B(2), Y => TMP_3_13_port);
   MUX21_K_2_14 : MUX21_L_81 port map( A => TMP_2_14_port, B => TMP_2_18_port, 
                           S => B(2), Y => TMP_3_14_port);
   MUX21_K_2_15 : MUX21_L_80 port map( A => TMP_2_15_port, B => TMP_2_19_port, 
                           S => B(2), Y => TMP_3_15_port);
   MUX21_K_2_16 : MUX21_L_79 port map( A => TMP_2_16_port, B => TMP_2_20_port, 
                           S => B(2), Y => TMP_3_16_port);
   MUX21_K_2_17 : MUX21_L_78 port map( A => TMP_2_17_port, B => TMP_2_21_port, 
                           S => B(2), Y => TMP_3_17_port);
   MUX21_K_2_18 : MUX21_L_77 port map( A => TMP_2_18_port, B => TMP_2_22_port, 
                           S => B(2), Y => TMP_3_18_port);
   MUX21_K_2_19 : MUX21_L_76 port map( A => TMP_2_19_port, B => TMP_2_23_port, 
                           S => B(2), Y => TMP_3_19_port);
   MUX21_K_2_20 : MUX21_L_75 port map( A => TMP_2_20_port, B => TMP_2_24_port, 
                           S => B(2), Y => TMP_3_20_port);
   MUX21_K_2_21 : MUX21_L_74 port map( A => TMP_2_21_port, B => TMP_2_25_port, 
                           S => B(2), Y => TMP_3_21_port);
   MUX21_K_2_22 : MUX21_L_73 port map( A => TMP_2_22_port, B => TMP_2_26_port, 
                           S => B(2), Y => TMP_3_22_port);
   MUX21_K_2_23 : MUX21_L_72 port map( A => TMP_2_23_port, B => TMP_2_27_port, 
                           S => B(2), Y => TMP_3_23_port);
   MUX21_K_2_24 : MUX21_L_71 port map( A => TMP_2_24_port, B => TMP_2_28_port, 
                           S => B(2), Y => TMP_3_24_port);
   MUX21_K_2_25 : MUX21_L_70 port map( A => TMP_2_25_port, B => TMP_2_29_port, 
                           S => B(2), Y => TMP_3_25_port);
   MUX21_K_2_26 : MUX21_L_69 port map( A => TMP_2_26_port, B => TMP_2_30_port, 
                           S => B(2), Y => TMP_3_26_port);
   MUX21_K_2_27 : MUX21_L_68 port map( A => TMP_2_27_port, B => TMP_2_31_port, 
                           S => B(2), Y => TMP_3_27_port);
   MUX21_J_2_0 : MUX21_L_67 port map( A => TMP_2_28_port, B => S, S => B(2), Y 
                           => TMP_3_28_port);
   MUX21_J_2_1 : MUX21_L_66 port map( A => TMP_2_29_port, B => S, S => B(2), Y 
                           => TMP_3_29_port);
   MUX21_J_2_2 : MUX21_L_65 port map( A => TMP_2_30_port, B => S, S => B(2), Y 
                           => TMP_3_30_port);
   MUX21_J_2_3 : MUX21_L_64 port map( A => TMP_2_31_port, B => S, S => B(2), Y 
                           => TMP_3_31_port);
   MUX21_K_3_0 : MUX21_L_63 port map( A => TMP_3_0_port, B => TMP_3_8_port, S 
                           => B(3), Y => TMP_4_0_port);
   MUX21_K_3_1 : MUX21_L_62 port map( A => TMP_3_1_port, B => TMP_3_9_port, S 
                           => B(3), Y => TMP_4_1_port);
   MUX21_K_3_2 : MUX21_L_61 port map( A => TMP_3_2_port, B => TMP_3_10_port, S 
                           => B(3), Y => TMP_4_2_port);
   MUX21_K_3_3 : MUX21_L_60 port map( A => TMP_3_3_port, B => TMP_3_11_port, S 
                           => B(3), Y => TMP_4_3_port);
   MUX21_K_3_4 : MUX21_L_59 port map( A => TMP_3_4_port, B => TMP_3_12_port, S 
                           => B(3), Y => TMP_4_4_port);
   MUX21_K_3_5 : MUX21_L_58 port map( A => TMP_3_5_port, B => TMP_3_13_port, S 
                           => B(3), Y => TMP_4_5_port);
   MUX21_K_3_6 : MUX21_L_57 port map( A => TMP_3_6_port, B => TMP_3_14_port, S 
                           => B(3), Y => TMP_4_6_port);
   MUX21_K_3_7 : MUX21_L_56 port map( A => TMP_3_7_port, B => TMP_3_15_port, S 
                           => B(3), Y => TMP_4_7_port);
   MUX21_K_3_8 : MUX21_L_55 port map( A => TMP_3_8_port, B => TMP_3_16_port, S 
                           => B(3), Y => TMP_4_8_port);
   MUX21_K_3_9 : MUX21_L_54 port map( A => TMP_3_9_port, B => TMP_3_17_port, S 
                           => B(3), Y => TMP_4_9_port);
   MUX21_K_3_10 : MUX21_L_53 port map( A => TMP_3_10_port, B => TMP_3_18_port, 
                           S => B(3), Y => TMP_4_10_port);
   MUX21_K_3_11 : MUX21_L_52 port map( A => TMP_3_11_port, B => TMP_3_19_port, 
                           S => B(3), Y => TMP_4_11_port);
   MUX21_K_3_12 : MUX21_L_51 port map( A => TMP_3_12_port, B => TMP_3_20_port, 
                           S => B(3), Y => TMP_4_12_port);
   MUX21_K_3_13 : MUX21_L_50 port map( A => TMP_3_13_port, B => TMP_3_21_port, 
                           S => B(3), Y => TMP_4_13_port);
   MUX21_K_3_14 : MUX21_L_49 port map( A => TMP_3_14_port, B => TMP_3_22_port, 
                           S => B(3), Y => TMP_4_14_port);
   MUX21_K_3_15 : MUX21_L_48 port map( A => TMP_3_15_port, B => TMP_3_23_port, 
                           S => B(3), Y => TMP_4_15_port);
   MUX21_K_3_16 : MUX21_L_47 port map( A => TMP_3_16_port, B => TMP_3_24_port, 
                           S => B(3), Y => TMP_4_16_port);
   MUX21_K_3_17 : MUX21_L_46 port map( A => TMP_3_17_port, B => TMP_3_25_port, 
                           S => B(3), Y => TMP_4_17_port);
   MUX21_K_3_18 : MUX21_L_45 port map( A => TMP_3_18_port, B => TMP_3_26_port, 
                           S => B(3), Y => TMP_4_18_port);
   MUX21_K_3_19 : MUX21_L_44 port map( A => TMP_3_19_port, B => TMP_3_27_port, 
                           S => B(3), Y => TMP_4_19_port);
   MUX21_K_3_20 : MUX21_L_43 port map( A => TMP_3_20_port, B => TMP_3_28_port, 
                           S => B(3), Y => TMP_4_20_port);
   MUX21_K_3_21 : MUX21_L_42 port map( A => TMP_3_21_port, B => TMP_3_29_port, 
                           S => B(3), Y => TMP_4_21_port);
   MUX21_K_3_22 : MUX21_L_41 port map( A => TMP_3_22_port, B => TMP_3_30_port, 
                           S => B(3), Y => TMP_4_22_port);
   MUX21_K_3_23 : MUX21_L_40 port map( A => TMP_3_23_port, B => TMP_3_31_port, 
                           S => B(3), Y => TMP_4_23_port);
   MUX21_J_3_0 : MUX21_L_39 port map( A => TMP_3_24_port, B => S, S => B(3), Y 
                           => TMP_4_24_port);
   MUX21_J_3_1 : MUX21_L_38 port map( A => TMP_3_25_port, B => S, S => B(3), Y 
                           => TMP_4_25_port);
   MUX21_J_3_2 : MUX21_L_37 port map( A => TMP_3_26_port, B => S, S => B(3), Y 
                           => TMP_4_26_port);
   MUX21_J_3_3 : MUX21_L_36 port map( A => TMP_3_27_port, B => S, S => B(3), Y 
                           => TMP_4_27_port);
   MUX21_J_3_4 : MUX21_L_35 port map( A => TMP_3_28_port, B => S, S => B(3), Y 
                           => TMP_4_28_port);
   MUX21_J_3_5 : MUX21_L_34 port map( A => TMP_3_29_port, B => S, S => B(3), Y 
                           => TMP_4_29_port);
   MUX21_J_3_6 : MUX21_L_33 port map( A => TMP_3_30_port, B => S, S => B(3), Y 
                           => TMP_4_30_port);
   MUX21_J_3_7 : MUX21_L_32 port map( A => TMP_3_31_port, B => S, S => B(3), Y 
                           => TMP_4_31_port);
   MUX21_K_4_0 : MUX21_L_31 port map( A => TMP_4_0_port, B => TMP_4_16_port, S 
                           => B(4), Y => Y(0));
   MUX21_K_4_1 : MUX21_L_30 port map( A => TMP_4_1_port, B => TMP_4_17_port, S 
                           => B(4), Y => Y(1));
   MUX21_K_4_2 : MUX21_L_29 port map( A => TMP_4_2_port, B => TMP_4_18_port, S 
                           => B(4), Y => Y(2));
   MUX21_K_4_3 : MUX21_L_28 port map( A => TMP_4_3_port, B => TMP_4_19_port, S 
                           => B(4), Y => Y(3));
   MUX21_K_4_4 : MUX21_L_27 port map( A => TMP_4_4_port, B => TMP_4_20_port, S 
                           => B(4), Y => Y(4));
   MUX21_K_4_5 : MUX21_L_26 port map( A => TMP_4_5_port, B => TMP_4_21_port, S 
                           => B(4), Y => Y(5));
   MUX21_K_4_6 : MUX21_L_25 port map( A => TMP_4_6_port, B => TMP_4_22_port, S 
                           => B(4), Y => Y(6));
   MUX21_K_4_7 : MUX21_L_24 port map( A => TMP_4_7_port, B => TMP_4_23_port, S 
                           => B(4), Y => Y(7));
   MUX21_K_4_8 : MUX21_L_23 port map( A => TMP_4_8_port, B => TMP_4_24_port, S 
                           => B(4), Y => Y(8));
   MUX21_K_4_9 : MUX21_L_22 port map( A => TMP_4_9_port, B => TMP_4_25_port, S 
                           => B(4), Y => Y(9));
   MUX21_K_4_10 : MUX21_L_21 port map( A => TMP_4_10_port, B => TMP_4_26_port, 
                           S => B(4), Y => Y(10));
   MUX21_K_4_11 : MUX21_L_20 port map( A => TMP_4_11_port, B => TMP_4_27_port, 
                           S => B(4), Y => Y(11));
   MUX21_K_4_12 : MUX21_L_19 port map( A => TMP_4_12_port, B => TMP_4_28_port, 
                           S => B(4), Y => Y(12));
   MUX21_K_4_13 : MUX21_L_18 port map( A => TMP_4_13_port, B => TMP_4_29_port, 
                           S => B(4), Y => Y(13));
   MUX21_K_4_14 : MUX21_L_17 port map( A => TMP_4_14_port, B => TMP_4_30_port, 
                           S => B(4), Y => Y(14));
   MUX21_K_4_15 : MUX21_L_16 port map( A => TMP_4_15_port, B => TMP_4_31_port, 
                           S => B(4), Y => Y(15));
   MUX21_J_4_0 : MUX21_L_15 port map( A => TMP_4_16_port, B => S, S => B(4), Y 
                           => Y(16));
   MUX21_J_4_1 : MUX21_L_14 port map( A => TMP_4_17_port, B => S, S => B(4), Y 
                           => Y(17));
   MUX21_J_4_2 : MUX21_L_13 port map( A => TMP_4_18_port, B => S, S => B(4), Y 
                           => Y(18));
   MUX21_J_4_3 : MUX21_L_12 port map( A => TMP_4_19_port, B => S, S => B(4), Y 
                           => Y(19));
   MUX21_J_4_4 : MUX21_L_11 port map( A => TMP_4_20_port, B => S, S => B(4), Y 
                           => Y(20));
   MUX21_J_4_5 : MUX21_L_10 port map( A => TMP_4_21_port, B => S, S => B(4), Y 
                           => Y(21));
   MUX21_J_4_6 : MUX21_L_9 port map( A => TMP_4_22_port, B => S, S => B(4), Y 
                           => Y(22));
   MUX21_J_4_7 : MUX21_L_8 port map( A => TMP_4_23_port, B => S, S => B(4), Y 
                           => Y(23));
   MUX21_J_4_8 : MUX21_L_7 port map( A => TMP_4_24_port, B => S, S => B(4), Y 
                           => Y(24));
   MUX21_J_4_9 : MUX21_L_6 port map( A => TMP_4_25_port, B => S, S => B(4), Y 
                           => Y(25));
   MUX21_J_4_10 : MUX21_L_5 port map( A => TMP_4_26_port, B => S, S => B(4), Y 
                           => Y(26));
   MUX21_J_4_11 : MUX21_L_4 port map( A => TMP_4_27_port, B => S, S => B(4), Y 
                           => Y(27));
   MUX21_J_4_12 : MUX21_L_3 port map( A => TMP_4_28_port, B => S, S => B(4), Y 
                           => Y(28));
   MUX21_J_4_13 : MUX21_L_2 port map( A => TMP_4_29_port, B => S, S => B(4), Y 
                           => Y(29));
   MUX21_J_4_14 : MUX21_L_1 port map( A => TMP_4_30_port, B => S, S => B(4), Y 
                           => Y(30));
   MUX21_J_4_15 : MUX21_L_0 port map( A => TMP_4_31_port, B => S, S => B(4), Y 
                           => Y(31));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BARREL_SHIFTER_LEFT_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
         (31 downto 0));

end BARREL_SHIFTER_LEFT_N32;

architecture SYN_STRUCTURAL of BARREL_SHIFTER_LEFT_N32 is

   component MUX21_L_160
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_161
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_162
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_163
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_164
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_165
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_166
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_167
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_168
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_169
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_170
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_171
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_172
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_173
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_174
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_175
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_176
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_177
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_178
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_179
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_180
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_181
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_182
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_183
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_184
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_185
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_186
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_187
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_188
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_189
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_190
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_191
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_192
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_193
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_194
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_195
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_196
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_197
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_198
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_199
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_200
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_201
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_202
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_203
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_204
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_205
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_206
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_207
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_208
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_209
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_210
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_211
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_212
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_213
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_214
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_215
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_216
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_217
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_218
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_219
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_220
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_221
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_222
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_223
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_224
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_225
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_226
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_227
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_228
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_229
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_230
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_231
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_232
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_233
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_234
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_235
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_236
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_237
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_238
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_239
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_240
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_241
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_242
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_243
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_244
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_245
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_246
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_247
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_248
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_249
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_250
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_251
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_252
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_253
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_254
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_255
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_256
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_257
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_258
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_259
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_260
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_261
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_262
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_263
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_264
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_265
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_266
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_267
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_268
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_269
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_270
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_271
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_272
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_273
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_274
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_275
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_276
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_277
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_278
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_279
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_280
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_281
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_282
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_283
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_284
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_285
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_286
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_287
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_288
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_289
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_290
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_291
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_292
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_293
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_294
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_295
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_296
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_297
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_298
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_299
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_300
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_301
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_302
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_303
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_304
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_305
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_306
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_307
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_308
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_309
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_310
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_311
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_312
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_313
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_314
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_315
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_316
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_317
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_318
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_L_319
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, TMP_4_31_port, TMP_4_30_port, TMP_4_29_port, 
      TMP_4_28_port, TMP_4_27_port, TMP_4_26_port, TMP_4_25_port, TMP_4_24_port
      , TMP_4_23_port, TMP_4_22_port, TMP_4_21_port, TMP_4_20_port, 
      TMP_4_19_port, TMP_4_18_port, TMP_4_17_port, TMP_4_16_port, TMP_4_15_port
      , TMP_4_14_port, TMP_4_13_port, TMP_4_12_port, TMP_4_11_port, 
      TMP_4_10_port, TMP_4_9_port, TMP_4_8_port, TMP_4_7_port, TMP_4_6_port, 
      TMP_4_5_port, TMP_4_4_port, TMP_4_3_port, TMP_4_2_port, TMP_4_1_port, 
      TMP_4_0_port, TMP_3_31_port, TMP_3_30_port, TMP_3_29_port, TMP_3_28_port,
      TMP_3_27_port, TMP_3_26_port, TMP_3_25_port, TMP_3_24_port, TMP_3_23_port
      , TMP_3_22_port, TMP_3_21_port, TMP_3_20_port, TMP_3_19_port, 
      TMP_3_18_port, TMP_3_17_port, TMP_3_16_port, TMP_3_15_port, TMP_3_14_port
      , TMP_3_13_port, TMP_3_12_port, TMP_3_11_port, TMP_3_10_port, 
      TMP_3_9_port, TMP_3_8_port, TMP_3_7_port, TMP_3_6_port, TMP_3_5_port, 
      TMP_3_4_port, TMP_3_3_port, TMP_3_2_port, TMP_3_1_port, TMP_3_0_port, 
      TMP_2_31_port, TMP_2_30_port, TMP_2_29_port, TMP_2_28_port, TMP_2_27_port
      , TMP_2_26_port, TMP_2_25_port, TMP_2_24_port, TMP_2_23_port, 
      TMP_2_22_port, TMP_2_21_port, TMP_2_20_port, TMP_2_19_port, TMP_2_18_port
      , TMP_2_17_port, TMP_2_16_port, TMP_2_15_port, TMP_2_14_port, 
      TMP_2_13_port, TMP_2_12_port, TMP_2_11_port, TMP_2_10_port, TMP_2_9_port,
      TMP_2_8_port, TMP_2_7_port, TMP_2_6_port, TMP_2_5_port, TMP_2_4_port, 
      TMP_2_3_port, TMP_2_2_port, TMP_2_1_port, TMP_2_0_port, TMP_1_31_port, 
      TMP_1_30_port, TMP_1_29_port, TMP_1_28_port, TMP_1_27_port, TMP_1_26_port
      , TMP_1_25_port, TMP_1_24_port, TMP_1_23_port, TMP_1_22_port, 
      TMP_1_21_port, TMP_1_20_port, TMP_1_19_port, TMP_1_18_port, TMP_1_17_port
      , TMP_1_16_port, TMP_1_15_port, TMP_1_14_port, TMP_1_13_port, 
      TMP_1_12_port, TMP_1_11_port, TMP_1_10_port, TMP_1_9_port, TMP_1_8_port, 
      TMP_1_7_port, TMP_1_6_port, TMP_1_5_port, TMP_1_4_port, TMP_1_3_port, 
      TMP_1_2_port, TMP_1_1_port, TMP_1_0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   MUX21_J_0_0 : MUX21_L_319 port map( A => A(0), B => X_Logic0_port, S => B(0)
                           , Y => TMP_1_0_port);
   MUX21_K_0_0 : MUX21_L_318 port map( A => A(1), B => A(0), S => B(0), Y => 
                           TMP_1_1_port);
   MUX21_K_0_1 : MUX21_L_317 port map( A => A(2), B => A(1), S => B(0), Y => 
                           TMP_1_2_port);
   MUX21_K_0_2 : MUX21_L_316 port map( A => A(3), B => A(2), S => B(0), Y => 
                           TMP_1_3_port);
   MUX21_K_0_3 : MUX21_L_315 port map( A => A(4), B => A(3), S => B(0), Y => 
                           TMP_1_4_port);
   MUX21_K_0_4 : MUX21_L_314 port map( A => A(5), B => A(4), S => B(0), Y => 
                           TMP_1_5_port);
   MUX21_K_0_5 : MUX21_L_313 port map( A => A(6), B => A(5), S => B(0), Y => 
                           TMP_1_6_port);
   MUX21_K_0_6 : MUX21_L_312 port map( A => A(7), B => A(6), S => B(0), Y => 
                           TMP_1_7_port);
   MUX21_K_0_7 : MUX21_L_311 port map( A => A(8), B => A(7), S => B(0), Y => 
                           TMP_1_8_port);
   MUX21_K_0_8 : MUX21_L_310 port map( A => A(9), B => A(8), S => B(0), Y => 
                           TMP_1_9_port);
   MUX21_K_0_9 : MUX21_L_309 port map( A => A(10), B => A(9), S => B(0), Y => 
                           TMP_1_10_port);
   MUX21_K_0_10 : MUX21_L_308 port map( A => A(11), B => A(10), S => B(0), Y =>
                           TMP_1_11_port);
   MUX21_K_0_11 : MUX21_L_307 port map( A => A(12), B => A(11), S => B(0), Y =>
                           TMP_1_12_port);
   MUX21_K_0_12 : MUX21_L_306 port map( A => A(13), B => A(12), S => B(0), Y =>
                           TMP_1_13_port);
   MUX21_K_0_13 : MUX21_L_305 port map( A => A(14), B => A(13), S => B(0), Y =>
                           TMP_1_14_port);
   MUX21_K_0_14 : MUX21_L_304 port map( A => A(15), B => A(14), S => B(0), Y =>
                           TMP_1_15_port);
   MUX21_K_0_15 : MUX21_L_303 port map( A => A(16), B => A(15), S => B(0), Y =>
                           TMP_1_16_port);
   MUX21_K_0_16 : MUX21_L_302 port map( A => A(17), B => A(16), S => B(0), Y =>
                           TMP_1_17_port);
   MUX21_K_0_17 : MUX21_L_301 port map( A => A(18), B => A(17), S => B(0), Y =>
                           TMP_1_18_port);
   MUX21_K_0_18 : MUX21_L_300 port map( A => A(19), B => A(18), S => B(0), Y =>
                           TMP_1_19_port);
   MUX21_K_0_19 : MUX21_L_299 port map( A => A(20), B => A(19), S => B(0), Y =>
                           TMP_1_20_port);
   MUX21_K_0_20 : MUX21_L_298 port map( A => A(21), B => A(20), S => B(0), Y =>
                           TMP_1_21_port);
   MUX21_K_0_21 : MUX21_L_297 port map( A => A(22), B => A(21), S => B(0), Y =>
                           TMP_1_22_port);
   MUX21_K_0_22 : MUX21_L_296 port map( A => A(23), B => A(22), S => B(0), Y =>
                           TMP_1_23_port);
   MUX21_K_0_23 : MUX21_L_295 port map( A => A(24), B => A(23), S => B(0), Y =>
                           TMP_1_24_port);
   MUX21_K_0_24 : MUX21_L_294 port map( A => A(25), B => A(24), S => B(0), Y =>
                           TMP_1_25_port);
   MUX21_K_0_25 : MUX21_L_293 port map( A => A(26), B => A(25), S => B(0), Y =>
                           TMP_1_26_port);
   MUX21_K_0_26 : MUX21_L_292 port map( A => A(27), B => A(26), S => B(0), Y =>
                           TMP_1_27_port);
   MUX21_K_0_27 : MUX21_L_291 port map( A => A(28), B => A(27), S => B(0), Y =>
                           TMP_1_28_port);
   MUX21_K_0_28 : MUX21_L_290 port map( A => A(29), B => A(28), S => B(0), Y =>
                           TMP_1_29_port);
   MUX21_K_0_29 : MUX21_L_289 port map( A => A(30), B => A(29), S => B(0), Y =>
                           TMP_1_30_port);
   MUX21_K_0_30 : MUX21_L_288 port map( A => A(31), B => A(30), S => B(0), Y =>
                           TMP_1_31_port);
   MUX21_J_1_0 : MUX21_L_287 port map( A => TMP_1_0_port, B => X_Logic0_port, S
                           => B(1), Y => TMP_2_0_port);
   MUX21_J_1_1 : MUX21_L_286 port map( A => TMP_1_1_port, B => X_Logic0_port, S
                           => B(1), Y => TMP_2_1_port);
   MUX21_K_1_0 : MUX21_L_285 port map( A => TMP_1_2_port, B => TMP_1_0_port, S 
                           => B(1), Y => TMP_2_2_port);
   MUX21_K_1_1 : MUX21_L_284 port map( A => TMP_1_3_port, B => TMP_1_1_port, S 
                           => B(1), Y => TMP_2_3_port);
   MUX21_K_1_2 : MUX21_L_283 port map( A => TMP_1_4_port, B => TMP_1_2_port, S 
                           => B(1), Y => TMP_2_4_port);
   MUX21_K_1_3 : MUX21_L_282 port map( A => TMP_1_5_port, B => TMP_1_3_port, S 
                           => B(1), Y => TMP_2_5_port);
   MUX21_K_1_4 : MUX21_L_281 port map( A => TMP_1_6_port, B => TMP_1_4_port, S 
                           => B(1), Y => TMP_2_6_port);
   MUX21_K_1_5 : MUX21_L_280 port map( A => TMP_1_7_port, B => TMP_1_5_port, S 
                           => B(1), Y => TMP_2_7_port);
   MUX21_K_1_6 : MUX21_L_279 port map( A => TMP_1_8_port, B => TMP_1_6_port, S 
                           => B(1), Y => TMP_2_8_port);
   MUX21_K_1_7 : MUX21_L_278 port map( A => TMP_1_9_port, B => TMP_1_7_port, S 
                           => B(1), Y => TMP_2_9_port);
   MUX21_K_1_8 : MUX21_L_277 port map( A => TMP_1_10_port, B => TMP_1_8_port, S
                           => B(1), Y => TMP_2_10_port);
   MUX21_K_1_9 : MUX21_L_276 port map( A => TMP_1_11_port, B => TMP_1_9_port, S
                           => B(1), Y => TMP_2_11_port);
   MUX21_K_1_10 : MUX21_L_275 port map( A => TMP_1_12_port, B => TMP_1_10_port,
                           S => B(1), Y => TMP_2_12_port);
   MUX21_K_1_11 : MUX21_L_274 port map( A => TMP_1_13_port, B => TMP_1_11_port,
                           S => B(1), Y => TMP_2_13_port);
   MUX21_K_1_12 : MUX21_L_273 port map( A => TMP_1_14_port, B => TMP_1_12_port,
                           S => B(1), Y => TMP_2_14_port);
   MUX21_K_1_13 : MUX21_L_272 port map( A => TMP_1_15_port, B => TMP_1_13_port,
                           S => B(1), Y => TMP_2_15_port);
   MUX21_K_1_14 : MUX21_L_271 port map( A => TMP_1_16_port, B => TMP_1_14_port,
                           S => B(1), Y => TMP_2_16_port);
   MUX21_K_1_15 : MUX21_L_270 port map( A => TMP_1_17_port, B => TMP_1_15_port,
                           S => B(1), Y => TMP_2_17_port);
   MUX21_K_1_16 : MUX21_L_269 port map( A => TMP_1_18_port, B => TMP_1_16_port,
                           S => B(1), Y => TMP_2_18_port);
   MUX21_K_1_17 : MUX21_L_268 port map( A => TMP_1_19_port, B => TMP_1_17_port,
                           S => B(1), Y => TMP_2_19_port);
   MUX21_K_1_18 : MUX21_L_267 port map( A => TMP_1_20_port, B => TMP_1_18_port,
                           S => B(1), Y => TMP_2_20_port);
   MUX21_K_1_19 : MUX21_L_266 port map( A => TMP_1_21_port, B => TMP_1_19_port,
                           S => B(1), Y => TMP_2_21_port);
   MUX21_K_1_20 : MUX21_L_265 port map( A => TMP_1_22_port, B => TMP_1_20_port,
                           S => B(1), Y => TMP_2_22_port);
   MUX21_K_1_21 : MUX21_L_264 port map( A => TMP_1_23_port, B => TMP_1_21_port,
                           S => B(1), Y => TMP_2_23_port);
   MUX21_K_1_22 : MUX21_L_263 port map( A => TMP_1_24_port, B => TMP_1_22_port,
                           S => B(1), Y => TMP_2_24_port);
   MUX21_K_1_23 : MUX21_L_262 port map( A => TMP_1_25_port, B => TMP_1_23_port,
                           S => B(1), Y => TMP_2_25_port);
   MUX21_K_1_24 : MUX21_L_261 port map( A => TMP_1_26_port, B => TMP_1_24_port,
                           S => B(1), Y => TMP_2_26_port);
   MUX21_K_1_25 : MUX21_L_260 port map( A => TMP_1_27_port, B => TMP_1_25_port,
                           S => B(1), Y => TMP_2_27_port);
   MUX21_K_1_26 : MUX21_L_259 port map( A => TMP_1_28_port, B => TMP_1_26_port,
                           S => B(1), Y => TMP_2_28_port);
   MUX21_K_1_27 : MUX21_L_258 port map( A => TMP_1_29_port, B => TMP_1_27_port,
                           S => B(1), Y => TMP_2_29_port);
   MUX21_K_1_28 : MUX21_L_257 port map( A => TMP_1_30_port, B => TMP_1_28_port,
                           S => B(1), Y => TMP_2_30_port);
   MUX21_K_1_29 : MUX21_L_256 port map( A => TMP_1_31_port, B => TMP_1_29_port,
                           S => B(1), Y => TMP_2_31_port);
   MUX21_J_2_0 : MUX21_L_255 port map( A => TMP_2_0_port, B => X_Logic0_port, S
                           => B(2), Y => TMP_3_0_port);
   MUX21_J_2_1 : MUX21_L_254 port map( A => TMP_2_1_port, B => X_Logic0_port, S
                           => B(2), Y => TMP_3_1_port);
   MUX21_J_2_2 : MUX21_L_253 port map( A => TMP_2_2_port, B => X_Logic0_port, S
                           => B(2), Y => TMP_3_2_port);
   MUX21_J_2_3 : MUX21_L_252 port map( A => TMP_2_3_port, B => X_Logic0_port, S
                           => B(2), Y => TMP_3_3_port);
   MUX21_K_2_0 : MUX21_L_251 port map( A => TMP_2_4_port, B => TMP_2_0_port, S 
                           => B(2), Y => TMP_3_4_port);
   MUX21_K_2_1 : MUX21_L_250 port map( A => TMP_2_5_port, B => TMP_2_1_port, S 
                           => B(2), Y => TMP_3_5_port);
   MUX21_K_2_2 : MUX21_L_249 port map( A => TMP_2_6_port, B => TMP_2_2_port, S 
                           => B(2), Y => TMP_3_6_port);
   MUX21_K_2_3 : MUX21_L_248 port map( A => TMP_2_7_port, B => TMP_2_3_port, S 
                           => B(2), Y => TMP_3_7_port);
   MUX21_K_2_4 : MUX21_L_247 port map( A => TMP_2_8_port, B => TMP_2_4_port, S 
                           => B(2), Y => TMP_3_8_port);
   MUX21_K_2_5 : MUX21_L_246 port map( A => TMP_2_9_port, B => TMP_2_5_port, S 
                           => B(2), Y => TMP_3_9_port);
   MUX21_K_2_6 : MUX21_L_245 port map( A => TMP_2_10_port, B => TMP_2_6_port, S
                           => B(2), Y => TMP_3_10_port);
   MUX21_K_2_7 : MUX21_L_244 port map( A => TMP_2_11_port, B => TMP_2_7_port, S
                           => B(2), Y => TMP_3_11_port);
   MUX21_K_2_8 : MUX21_L_243 port map( A => TMP_2_12_port, B => TMP_2_8_port, S
                           => B(2), Y => TMP_3_12_port);
   MUX21_K_2_9 : MUX21_L_242 port map( A => TMP_2_13_port, B => TMP_2_9_port, S
                           => B(2), Y => TMP_3_13_port);
   MUX21_K_2_10 : MUX21_L_241 port map( A => TMP_2_14_port, B => TMP_2_10_port,
                           S => B(2), Y => TMP_3_14_port);
   MUX21_K_2_11 : MUX21_L_240 port map( A => TMP_2_15_port, B => TMP_2_11_port,
                           S => B(2), Y => TMP_3_15_port);
   MUX21_K_2_12 : MUX21_L_239 port map( A => TMP_2_16_port, B => TMP_2_12_port,
                           S => B(2), Y => TMP_3_16_port);
   MUX21_K_2_13 : MUX21_L_238 port map( A => TMP_2_17_port, B => TMP_2_13_port,
                           S => B(2), Y => TMP_3_17_port);
   MUX21_K_2_14 : MUX21_L_237 port map( A => TMP_2_18_port, B => TMP_2_14_port,
                           S => B(2), Y => TMP_3_18_port);
   MUX21_K_2_15 : MUX21_L_236 port map( A => TMP_2_19_port, B => TMP_2_15_port,
                           S => B(2), Y => TMP_3_19_port);
   MUX21_K_2_16 : MUX21_L_235 port map( A => TMP_2_20_port, B => TMP_2_16_port,
                           S => B(2), Y => TMP_3_20_port);
   MUX21_K_2_17 : MUX21_L_234 port map( A => TMP_2_21_port, B => TMP_2_17_port,
                           S => B(2), Y => TMP_3_21_port);
   MUX21_K_2_18 : MUX21_L_233 port map( A => TMP_2_22_port, B => TMP_2_18_port,
                           S => B(2), Y => TMP_3_22_port);
   MUX21_K_2_19 : MUX21_L_232 port map( A => TMP_2_23_port, B => TMP_2_19_port,
                           S => B(2), Y => TMP_3_23_port);
   MUX21_K_2_20 : MUX21_L_231 port map( A => TMP_2_24_port, B => TMP_2_20_port,
                           S => B(2), Y => TMP_3_24_port);
   MUX21_K_2_21 : MUX21_L_230 port map( A => TMP_2_25_port, B => TMP_2_21_port,
                           S => B(2), Y => TMP_3_25_port);
   MUX21_K_2_22 : MUX21_L_229 port map( A => TMP_2_26_port, B => TMP_2_22_port,
                           S => B(2), Y => TMP_3_26_port);
   MUX21_K_2_23 : MUX21_L_228 port map( A => TMP_2_27_port, B => TMP_2_23_port,
                           S => B(2), Y => TMP_3_27_port);
   MUX21_K_2_24 : MUX21_L_227 port map( A => TMP_2_28_port, B => TMP_2_24_port,
                           S => B(2), Y => TMP_3_28_port);
   MUX21_K_2_25 : MUX21_L_226 port map( A => TMP_2_29_port, B => TMP_2_25_port,
                           S => B(2), Y => TMP_3_29_port);
   MUX21_K_2_26 : MUX21_L_225 port map( A => TMP_2_30_port, B => TMP_2_26_port,
                           S => B(2), Y => TMP_3_30_port);
   MUX21_K_2_27 : MUX21_L_224 port map( A => TMP_2_31_port, B => TMP_2_27_port,
                           S => B(2), Y => TMP_3_31_port);
   MUX21_J_3_0 : MUX21_L_223 port map( A => TMP_3_0_port, B => X_Logic0_port, S
                           => B(3), Y => TMP_4_0_port);
   MUX21_J_3_1 : MUX21_L_222 port map( A => TMP_3_1_port, B => X_Logic0_port, S
                           => B(3), Y => TMP_4_1_port);
   MUX21_J_3_2 : MUX21_L_221 port map( A => TMP_3_2_port, B => X_Logic0_port, S
                           => B(3), Y => TMP_4_2_port);
   MUX21_J_3_3 : MUX21_L_220 port map( A => TMP_3_3_port, B => X_Logic0_port, S
                           => B(3), Y => TMP_4_3_port);
   MUX21_J_3_4 : MUX21_L_219 port map( A => TMP_3_4_port, B => X_Logic0_port, S
                           => B(3), Y => TMP_4_4_port);
   MUX21_J_3_5 : MUX21_L_218 port map( A => TMP_3_5_port, B => X_Logic0_port, S
                           => B(3), Y => TMP_4_5_port);
   MUX21_J_3_6 : MUX21_L_217 port map( A => TMP_3_6_port, B => X_Logic0_port, S
                           => B(3), Y => TMP_4_6_port);
   MUX21_J_3_7 : MUX21_L_216 port map( A => TMP_3_7_port, B => X_Logic0_port, S
                           => B(3), Y => TMP_4_7_port);
   MUX21_K_3_0 : MUX21_L_215 port map( A => TMP_3_8_port, B => TMP_3_0_port, S 
                           => B(3), Y => TMP_4_8_port);
   MUX21_K_3_1 : MUX21_L_214 port map( A => TMP_3_9_port, B => TMP_3_1_port, S 
                           => B(3), Y => TMP_4_9_port);
   MUX21_K_3_2 : MUX21_L_213 port map( A => TMP_3_10_port, B => TMP_3_2_port, S
                           => B(3), Y => TMP_4_10_port);
   MUX21_K_3_3 : MUX21_L_212 port map( A => TMP_3_11_port, B => TMP_3_3_port, S
                           => B(3), Y => TMP_4_11_port);
   MUX21_K_3_4 : MUX21_L_211 port map( A => TMP_3_12_port, B => TMP_3_4_port, S
                           => B(3), Y => TMP_4_12_port);
   MUX21_K_3_5 : MUX21_L_210 port map( A => TMP_3_13_port, B => TMP_3_5_port, S
                           => B(3), Y => TMP_4_13_port);
   MUX21_K_3_6 : MUX21_L_209 port map( A => TMP_3_14_port, B => TMP_3_6_port, S
                           => B(3), Y => TMP_4_14_port);
   MUX21_K_3_7 : MUX21_L_208 port map( A => TMP_3_15_port, B => TMP_3_7_port, S
                           => B(3), Y => TMP_4_15_port);
   MUX21_K_3_8 : MUX21_L_207 port map( A => TMP_3_16_port, B => TMP_3_8_port, S
                           => B(3), Y => TMP_4_16_port);
   MUX21_K_3_9 : MUX21_L_206 port map( A => TMP_3_17_port, B => TMP_3_9_port, S
                           => B(3), Y => TMP_4_17_port);
   MUX21_K_3_10 : MUX21_L_205 port map( A => TMP_3_18_port, B => TMP_3_10_port,
                           S => B(3), Y => TMP_4_18_port);
   MUX21_K_3_11 : MUX21_L_204 port map( A => TMP_3_19_port, B => TMP_3_11_port,
                           S => B(3), Y => TMP_4_19_port);
   MUX21_K_3_12 : MUX21_L_203 port map( A => TMP_3_20_port, B => TMP_3_12_port,
                           S => B(3), Y => TMP_4_20_port);
   MUX21_K_3_13 : MUX21_L_202 port map( A => TMP_3_21_port, B => TMP_3_13_port,
                           S => B(3), Y => TMP_4_21_port);
   MUX21_K_3_14 : MUX21_L_201 port map( A => TMP_3_22_port, B => TMP_3_14_port,
                           S => B(3), Y => TMP_4_22_port);
   MUX21_K_3_15 : MUX21_L_200 port map( A => TMP_3_23_port, B => TMP_3_15_port,
                           S => B(3), Y => TMP_4_23_port);
   MUX21_K_3_16 : MUX21_L_199 port map( A => TMP_3_24_port, B => TMP_3_16_port,
                           S => B(3), Y => TMP_4_24_port);
   MUX21_K_3_17 : MUX21_L_198 port map( A => TMP_3_25_port, B => TMP_3_17_port,
                           S => B(3), Y => TMP_4_25_port);
   MUX21_K_3_18 : MUX21_L_197 port map( A => TMP_3_26_port, B => TMP_3_18_port,
                           S => B(3), Y => TMP_4_26_port);
   MUX21_K_3_19 : MUX21_L_196 port map( A => TMP_3_27_port, B => TMP_3_19_port,
                           S => B(3), Y => TMP_4_27_port);
   MUX21_K_3_20 : MUX21_L_195 port map( A => TMP_3_28_port, B => TMP_3_20_port,
                           S => B(3), Y => TMP_4_28_port);
   MUX21_K_3_21 : MUX21_L_194 port map( A => TMP_3_29_port, B => TMP_3_21_port,
                           S => B(3), Y => TMP_4_29_port);
   MUX21_K_3_22 : MUX21_L_193 port map( A => TMP_3_30_port, B => TMP_3_22_port,
                           S => B(3), Y => TMP_4_30_port);
   MUX21_K_3_23 : MUX21_L_192 port map( A => TMP_3_31_port, B => TMP_3_23_port,
                           S => B(3), Y => TMP_4_31_port);
   MUX21_J_4_0 : MUX21_L_191 port map( A => TMP_4_0_port, B => X_Logic0_port, S
                           => B(4), Y => Y(0));
   MUX21_J_4_1 : MUX21_L_190 port map( A => TMP_4_1_port, B => X_Logic0_port, S
                           => B(4), Y => Y(1));
   MUX21_J_4_2 : MUX21_L_189 port map( A => TMP_4_2_port, B => X_Logic0_port, S
                           => B(4), Y => Y(2));
   MUX21_J_4_3 : MUX21_L_188 port map( A => TMP_4_3_port, B => X_Logic0_port, S
                           => B(4), Y => Y(3));
   MUX21_J_4_4 : MUX21_L_187 port map( A => TMP_4_4_port, B => X_Logic0_port, S
                           => B(4), Y => Y(4));
   MUX21_J_4_5 : MUX21_L_186 port map( A => TMP_4_5_port, B => X_Logic0_port, S
                           => B(4), Y => Y(5));
   MUX21_J_4_6 : MUX21_L_185 port map( A => TMP_4_6_port, B => X_Logic0_port, S
                           => B(4), Y => Y(6));
   MUX21_J_4_7 : MUX21_L_184 port map( A => TMP_4_7_port, B => X_Logic0_port, S
                           => B(4), Y => Y(7));
   MUX21_J_4_8 : MUX21_L_183 port map( A => TMP_4_8_port, B => X_Logic0_port, S
                           => B(4), Y => Y(8));
   MUX21_J_4_9 : MUX21_L_182 port map( A => TMP_4_9_port, B => X_Logic0_port, S
                           => B(4), Y => Y(9));
   MUX21_J_4_10 : MUX21_L_181 port map( A => TMP_4_10_port, B => X_Logic0_port,
                           S => B(4), Y => Y(10));
   MUX21_J_4_11 : MUX21_L_180 port map( A => TMP_4_11_port, B => X_Logic0_port,
                           S => B(4), Y => Y(11));
   MUX21_J_4_12 : MUX21_L_179 port map( A => TMP_4_12_port, B => X_Logic0_port,
                           S => B(4), Y => Y(12));
   MUX21_J_4_13 : MUX21_L_178 port map( A => TMP_4_13_port, B => X_Logic0_port,
                           S => B(4), Y => Y(13));
   MUX21_J_4_14 : MUX21_L_177 port map( A => TMP_4_14_port, B => X_Logic0_port,
                           S => B(4), Y => Y(14));
   MUX21_J_4_15 : MUX21_L_176 port map( A => TMP_4_15_port, B => X_Logic0_port,
                           S => B(4), Y => Y(15));
   MUX21_K_4_0 : MUX21_L_175 port map( A => TMP_4_16_port, B => TMP_4_0_port, S
                           => B(4), Y => Y(16));
   MUX21_K_4_1 : MUX21_L_174 port map( A => TMP_4_17_port, B => TMP_4_1_port, S
                           => B(4), Y => Y(17));
   MUX21_K_4_2 : MUX21_L_173 port map( A => TMP_4_18_port, B => TMP_4_2_port, S
                           => B(4), Y => Y(18));
   MUX21_K_4_3 : MUX21_L_172 port map( A => TMP_4_19_port, B => TMP_4_3_port, S
                           => B(4), Y => Y(19));
   MUX21_K_4_4 : MUX21_L_171 port map( A => TMP_4_20_port, B => TMP_4_4_port, S
                           => B(4), Y => Y(20));
   MUX21_K_4_5 : MUX21_L_170 port map( A => TMP_4_21_port, B => TMP_4_5_port, S
                           => B(4), Y => Y(21));
   MUX21_K_4_6 : MUX21_L_169 port map( A => TMP_4_22_port, B => TMP_4_6_port, S
                           => B(4), Y => Y(22));
   MUX21_K_4_7 : MUX21_L_168 port map( A => TMP_4_23_port, B => TMP_4_7_port, S
                           => B(4), Y => Y(23));
   MUX21_K_4_8 : MUX21_L_167 port map( A => TMP_4_24_port, B => TMP_4_8_port, S
                           => B(4), Y => Y(24));
   MUX21_K_4_9 : MUX21_L_166 port map( A => TMP_4_25_port, B => TMP_4_9_port, S
                           => B(4), Y => Y(25));
   MUX21_K_4_10 : MUX21_L_165 port map( A => TMP_4_26_port, B => TMP_4_10_port,
                           S => B(4), Y => Y(26));
   MUX21_K_4_11 : MUX21_L_164 port map( A => TMP_4_27_port, B => TMP_4_11_port,
                           S => B(4), Y => Y(27));
   MUX21_K_4_12 : MUX21_L_163 port map( A => TMP_4_28_port, B => TMP_4_12_port,
                           S => B(4), Y => Y(28));
   MUX21_K_4_13 : MUX21_L_162 port map( A => TMP_4_29_port, B => TMP_4_13_port,
                           S => B(4), Y => Y(29));
   MUX21_K_4_14 : MUX21_L_161 port map( A => TMP_4_30_port, B => TMP_4_14_port,
                           S => B(4), Y => Y(30));
   MUX21_K_4_15 : MUX21_L_160 port map( A => TMP_4_31_port, B => TMP_4_15_port,
                           S => B(4), Y => Y(31));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BOOTH_MULTIPLIER_N32 is

   port( A, B : in std_logic_vector (15 downto 0);  P : out std_logic_vector 
         (31 downto 0));

end BOOTH_MULTIPLIER_N32;

architecture SYN_STRUCTURAL of BOOTH_MULTIPLIER_N32 is

   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component MUX81_N32_0
      port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component RCA_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component MUX81_N32_1
      port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component RCA_N32_2
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component MUX81_N32_2
      port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX81_N32_3
      port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  S : in
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component BOOTH_ENCODER_N16
      port( B : in std_logic_vector (15 downto 0);  Bo : out std_logic_vector 
            (23 downto 0));
   end component;
   
   signal X_Logic0_port, Bo_signal_11_port, Bo_signal_10_port, Bo_signal_9_port
      , Bo_signal_8_port, Bo_signal_7_port, Bo_signal_6_port, Bo_signal_5_port,
      Bo_signal_4_port, Bo_signal_3_port, Bo_signal_2_port, Bo_signal_1_port, 
      Bo_signal_0_port, aMatrix_15_0_port, aMatrix_13_0_port, aMatrix_11_0_port
      , aMatrix_9_31_port, aMatrix_9_19_port, aMatrix_9_18_port, 
      aMatrix_9_17_port, aMatrix_9_16_port, aMatrix_9_15_port, 
      aMatrix_9_14_port, aMatrix_9_13_port, aMatrix_9_12_port, 
      aMatrix_9_11_port, aMatrix_9_10_port, aMatrix_9_9_port, aMatrix_9_8_port,
      aMatrix_9_7_port, aMatrix_9_6_port, aMatrix_9_5_port, aMatrix_9_0_port, 
      aMatrix_7_0_port, aMatrix_5_0_port, aMatrix_3_0_port, 
      aEncMatrix_3_31_port, aEncMatrix_3_30_port, aEncMatrix_3_29_port, 
      aEncMatrix_3_28_port, aEncMatrix_3_27_port, aEncMatrix_3_26_port, 
      aEncMatrix_3_25_port, aEncMatrix_3_24_port, aEncMatrix_3_23_port, 
      aEncMatrix_3_22_port, aEncMatrix_3_21_port, aEncMatrix_3_20_port, 
      aEncMatrix_3_19_port, aEncMatrix_3_18_port, aEncMatrix_3_17_port, 
      aEncMatrix_3_16_port, aEncMatrix_3_15_port, aEncMatrix_3_14_port, 
      aEncMatrix_3_13_port, aEncMatrix_3_12_port, aEncMatrix_3_11_port, 
      aEncMatrix_3_10_port, aEncMatrix_3_9_port, aEncMatrix_3_8_port, 
      aEncMatrix_3_7_port, aEncMatrix_3_6_port, aEncMatrix_3_5_port, 
      aEncMatrix_3_4_port, aEncMatrix_3_3_port, aEncMatrix_3_2_port, 
      aEncMatrix_3_1_port, aEncMatrix_3_0_port, aEncMatrix_2_31_port, 
      aEncMatrix_2_30_port, aEncMatrix_2_29_port, aEncMatrix_2_28_port, 
      aEncMatrix_2_27_port, aEncMatrix_2_26_port, aEncMatrix_2_25_port, 
      aEncMatrix_2_24_port, aEncMatrix_2_23_port, aEncMatrix_2_22_port, 
      aEncMatrix_2_21_port, aEncMatrix_2_20_port, aEncMatrix_2_19_port, 
      aEncMatrix_2_18_port, aEncMatrix_2_17_port, aEncMatrix_2_16_port, 
      aEncMatrix_2_15_port, aEncMatrix_2_14_port, aEncMatrix_2_13_port, 
      aEncMatrix_2_12_port, aEncMatrix_2_11_port, aEncMatrix_2_10_port, 
      aEncMatrix_2_9_port, aEncMatrix_2_8_port, aEncMatrix_2_7_port, 
      aEncMatrix_2_6_port, aEncMatrix_2_5_port, aEncMatrix_2_4_port, 
      aEncMatrix_2_3_port, aEncMatrix_2_2_port, aEncMatrix_2_1_port, 
      aEncMatrix_2_0_port, aEncMatrix_1_31_port, aEncMatrix_1_30_port, 
      aEncMatrix_1_29_port, aEncMatrix_1_28_port, aEncMatrix_1_27_port, 
      aEncMatrix_1_26_port, aEncMatrix_1_25_port, aEncMatrix_1_24_port, 
      aEncMatrix_1_23_port, aEncMatrix_1_22_port, aEncMatrix_1_21_port, 
      aEncMatrix_1_20_port, aEncMatrix_1_19_port, aEncMatrix_1_18_port, 
      aEncMatrix_1_17_port, aEncMatrix_1_16_port, aEncMatrix_1_15_port, 
      aEncMatrix_1_14_port, aEncMatrix_1_13_port, aEncMatrix_1_12_port, 
      aEncMatrix_1_11_port, aEncMatrix_1_10_port, aEncMatrix_1_9_port, 
      aEncMatrix_1_8_port, aEncMatrix_1_7_port, aEncMatrix_1_6_port, 
      aEncMatrix_1_5_port, aEncMatrix_1_4_port, aEncMatrix_1_3_port, 
      aEncMatrix_1_2_port, aEncMatrix_1_1_port, aEncMatrix_1_0_port, 
      aEncMatrix_0_31_port, aEncMatrix_0_30_port, aEncMatrix_0_29_port, 
      aEncMatrix_0_28_port, aEncMatrix_0_27_port, aEncMatrix_0_26_port, 
      aEncMatrix_0_25_port, aEncMatrix_0_24_port, aEncMatrix_0_23_port, 
      aEncMatrix_0_22_port, aEncMatrix_0_21_port, aEncMatrix_0_20_port, 
      aEncMatrix_0_19_port, aEncMatrix_0_18_port, aEncMatrix_0_17_port, 
      aEncMatrix_0_16_port, aEncMatrix_0_15_port, aEncMatrix_0_14_port, 
      aEncMatrix_0_13_port, aEncMatrix_0_12_port, aEncMatrix_0_11_port, 
      aEncMatrix_0_10_port, aEncMatrix_0_9_port, aEncMatrix_0_8_port, 
      aEncMatrix_0_7_port, aEncMatrix_0_6_port, aEncMatrix_0_5_port, 
      aEncMatrix_0_4_port, aEncMatrix_0_3_port, aEncMatrix_0_2_port, 
      aEncMatrix_0_1_port, aEncMatrix_0_0_port, pSumMatrix_1_31_port, 
      pSumMatrix_1_30_port, pSumMatrix_1_29_port, pSumMatrix_1_28_port, 
      pSumMatrix_1_27_port, pSumMatrix_1_26_port, pSumMatrix_1_25_port, 
      pSumMatrix_1_24_port, pSumMatrix_1_23_port, pSumMatrix_1_22_port, 
      pSumMatrix_1_21_port, pSumMatrix_1_20_port, pSumMatrix_1_19_port, 
      pSumMatrix_1_18_port, pSumMatrix_1_17_port, pSumMatrix_1_16_port, 
      pSumMatrix_1_15_port, pSumMatrix_1_14_port, pSumMatrix_1_13_port, 
      pSumMatrix_1_12_port, pSumMatrix_1_11_port, pSumMatrix_1_10_port, 
      pSumMatrix_1_9_port, pSumMatrix_1_8_port, pSumMatrix_1_7_port, 
      pSumMatrix_1_6_port, pSumMatrix_1_5_port, pSumMatrix_1_4_port, 
      pSumMatrix_1_3_port, pSumMatrix_1_2_port, pSumMatrix_1_1_port, 
      pSumMatrix_1_0_port, pSumMatrix_0_31_port, pSumMatrix_0_30_port, 
      pSumMatrix_0_29_port, pSumMatrix_0_28_port, pSumMatrix_0_27_port, 
      pSumMatrix_0_26_port, pSumMatrix_0_25_port, pSumMatrix_0_24_port, 
      pSumMatrix_0_23_port, pSumMatrix_0_22_port, pSumMatrix_0_21_port, 
      pSumMatrix_0_20_port, pSumMatrix_0_19_port, pSumMatrix_0_18_port, 
      pSumMatrix_0_17_port, pSumMatrix_0_16_port, pSumMatrix_0_15_port, 
      pSumMatrix_0_14_port, pSumMatrix_0_13_port, pSumMatrix_0_12_port, 
      pSumMatrix_0_11_port, pSumMatrix_0_10_port, pSumMatrix_0_9_port, 
      pSumMatrix_0_8_port, pSumMatrix_0_7_port, pSumMatrix_0_6_port, 
      pSumMatrix_0_5_port, pSumMatrix_0_4_port, pSumMatrix_0_3_port, 
      pSumMatrix_0_2_port, pSumMatrix_0_1_port, pSumMatrix_0_0_port, n1, n2, n3
      , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275,
      n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282 : std_logic;

begin
   
   X_Logic0_port <= '0';
   B_INSTANCE : BOOTH_ENCODER_N16 port map( B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           Bo(23) => n_1268, Bo(22) => n_1269, Bo(21) => n_1270
                           , Bo(20) => n_1271, Bo(19) => n_1272, Bo(18) => 
                           n_1273, Bo(17) => n_1274, Bo(16) => n_1275, Bo(15) 
                           => n_1276, Bo(14) => n_1277, Bo(13) => n_1278, 
                           Bo(12) => n_1279, Bo(11) => Bo_signal_11_port, 
                           Bo(10) => Bo_signal_10_port, Bo(9) => 
                           Bo_signal_9_port, Bo(8) => Bo_signal_8_port, Bo(7) 
                           => Bo_signal_7_port, Bo(6) => Bo_signal_6_port, 
                           Bo(5) => Bo_signal_5_port, Bo(4) => Bo_signal_4_port
                           , Bo(3) => Bo_signal_3_port, Bo(2) => 
                           Bo_signal_2_port, Bo(1) => Bo_signal_1_port, Bo(0) 
                           => Bo_signal_0_port);
   FIRST_MUX : MUX81_N32_3 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => A(15), B(30) => A(15), B(29)
                           => A(15), B(28) => A(15), B(27) => A(15), B(26) => 
                           A(15), B(25) => A(15), B(24) => A(15), B(23) => 
                           A(15), B(22) => A(15), B(21) => A(15), B(20) => 
                           A(15), B(19) => A(15), B(18) => A(15), B(17) => 
                           A(15), B(16) => A(15), B(15) => A(15), B(14) => 
                           A(14), B(13) => A(13), B(12) => A(12), B(11) => 
                           A(11), B(10) => A(10), B(9) => A(9), B(8) => A(8), 
                           B(7) => A(7), B(6) => A(6), B(5) => A(5), B(4) => 
                           A(4), B(3) => A(3), B(2) => A(2), B(1) => A(1), B(0)
                           => A(0), C(31) => aMatrix_9_31_port, C(30) => 
                           aMatrix_9_31_port, C(29) => aMatrix_9_31_port, C(28)
                           => aMatrix_9_31_port, C(27) => aMatrix_9_31_port, 
                           C(26) => aMatrix_9_31_port, C(25) => 
                           aMatrix_9_31_port, C(24) => aMatrix_9_31_port, C(23)
                           => aMatrix_9_31_port, C(22) => aMatrix_9_31_port, 
                           C(21) => aMatrix_9_31_port, C(20) => 
                           aMatrix_9_31_port, C(19) => aMatrix_9_31_port, C(18)
                           => aMatrix_9_31_port, C(17) => aMatrix_9_31_port, 
                           C(16) => aMatrix_9_31_port, C(15) => 
                           aMatrix_9_19_port, C(14) => aMatrix_9_18_port, C(13)
                           => aMatrix_9_17_port, C(12) => aMatrix_9_16_port, 
                           C(11) => aMatrix_9_15_port, C(10) => 
                           aMatrix_9_14_port, C(9) => aMatrix_9_13_port, C(8) 
                           => aMatrix_9_12_port, C(7) => aMatrix_9_11_port, 
                           C(6) => aMatrix_9_10_port, C(5) => aMatrix_9_9_port,
                           C(4) => aMatrix_9_8_port, C(3) => aMatrix_9_7_port, 
                           C(2) => aMatrix_9_6_port, C(1) => aMatrix_9_5_port, 
                           C(0) => A(0), D(31) => A(15), D(30) => A(15), D(29) 
                           => A(15), D(28) => A(15), D(27) => A(15), D(26) => 
                           A(15), D(25) => A(15), D(24) => A(15), D(23) => 
                           A(15), D(22) => A(15), D(21) => A(15), D(20) => 
                           A(15), D(19) => A(15), D(18) => A(15), D(17) => 
                           A(15), D(16) => A(15), D(15) => A(14), D(14) => 
                           A(13), D(13) => A(12), D(12) => A(11), D(11) => 
                           A(10), D(10) => A(9), D(9) => A(8), D(8) => A(7), 
                           D(7) => A(6), D(6) => A(5), D(5) => A(4), D(4) => 
                           A(3), D(3) => A(2), D(2) => A(1), D(1) => A(0), D(0)
                           => X_Logic0_port, E(31) => aMatrix_9_31_port, E(30) 
                           => aMatrix_9_31_port, E(29) => aMatrix_9_31_port, 
                           E(28) => aMatrix_9_31_port, E(27) => 
                           aMatrix_9_31_port, E(26) => aMatrix_9_31_port, E(25)
                           => aMatrix_9_31_port, E(24) => aMatrix_9_31_port, 
                           E(23) => aMatrix_9_31_port, E(22) => 
                           aMatrix_9_31_port, E(21) => aMatrix_9_31_port, E(20)
                           => aMatrix_9_31_port, E(19) => aMatrix_9_31_port, 
                           E(18) => aMatrix_9_31_port, E(17) => 
                           aMatrix_9_31_port, E(16) => aMatrix_9_19_port, E(15)
                           => aMatrix_9_18_port, E(14) => aMatrix_9_17_port, 
                           E(13) => aMatrix_9_16_port, E(12) => 
                           aMatrix_9_15_port, E(11) => aMatrix_9_14_port, E(10)
                           => aMatrix_9_13_port, E(9) => aMatrix_9_12_port, 
                           E(8) => aMatrix_9_11_port, E(7) => aMatrix_9_10_port
                           , E(6) => aMatrix_9_9_port, E(5) => aMatrix_9_8_port
                           , E(4) => aMatrix_9_7_port, E(3) => aMatrix_9_6_port
                           , E(2) => aMatrix_9_5_port, E(1) => A(0), E(0) => 
                           aMatrix_3_0_port, F(31) => X_Logic0_port, F(30) => 
                           X_Logic0_port, F(29) => X_Logic0_port, F(28) => 
                           X_Logic0_port, F(27) => X_Logic0_port, F(26) => 
                           X_Logic0_port, F(25) => X_Logic0_port, F(24) => 
                           X_Logic0_port, F(23) => X_Logic0_port, F(22) => 
                           X_Logic0_port, F(21) => X_Logic0_port, F(20) => 
                           X_Logic0_port, F(19) => X_Logic0_port, F(18) => 
                           X_Logic0_port, F(17) => X_Logic0_port, F(16) => 
                           X_Logic0_port, F(15) => X_Logic0_port, F(14) => 
                           X_Logic0_port, F(13) => X_Logic0_port, F(12) => 
                           X_Logic0_port, F(11) => X_Logic0_port, F(10) => 
                           X_Logic0_port, F(9) => X_Logic0_port, F(8) => 
                           X_Logic0_port, F(7) => X_Logic0_port, F(6) => 
                           X_Logic0_port, F(5) => X_Logic0_port, F(4) => 
                           X_Logic0_port, F(3) => X_Logic0_port, F(2) => 
                           X_Logic0_port, F(1) => X_Logic0_port, F(0) => 
                           X_Logic0_port, G(31) => X_Logic0_port, G(30) => 
                           X_Logic0_port, G(29) => X_Logic0_port, G(28) => 
                           X_Logic0_port, G(27) => X_Logic0_port, G(26) => 
                           X_Logic0_port, G(25) => X_Logic0_port, G(24) => 
                           X_Logic0_port, G(23) => X_Logic0_port, G(22) => 
                           X_Logic0_port, G(21) => X_Logic0_port, G(20) => 
                           X_Logic0_port, G(19) => X_Logic0_port, G(18) => 
                           X_Logic0_port, G(17) => X_Logic0_port, G(16) => 
                           X_Logic0_port, G(15) => X_Logic0_port, G(14) => 
                           X_Logic0_port, G(13) => X_Logic0_port, G(12) => 
                           X_Logic0_port, G(11) => X_Logic0_port, G(10) => 
                           X_Logic0_port, G(9) => X_Logic0_port, G(8) => 
                           X_Logic0_port, G(7) => X_Logic0_port, G(6) => 
                           X_Logic0_port, G(5) => X_Logic0_port, G(4) => 
                           X_Logic0_port, G(3) => X_Logic0_port, G(2) => 
                           X_Logic0_port, G(1) => X_Logic0_port, G(0) => 
                           X_Logic0_port, H(31) => X_Logic0_port, H(30) => 
                           X_Logic0_port, H(29) => X_Logic0_port, H(28) => 
                           X_Logic0_port, H(27) => X_Logic0_port, H(26) => 
                           X_Logic0_port, H(25) => X_Logic0_port, H(24) => 
                           X_Logic0_port, H(23) => X_Logic0_port, H(22) => 
                           X_Logic0_port, H(21) => X_Logic0_port, H(20) => 
                           X_Logic0_port, H(19) => X_Logic0_port, H(18) => 
                           X_Logic0_port, H(17) => X_Logic0_port, H(16) => 
                           X_Logic0_port, H(15) => X_Logic0_port, H(14) => 
                           X_Logic0_port, H(13) => X_Logic0_port, H(12) => 
                           X_Logic0_port, H(11) => X_Logic0_port, H(10) => 
                           X_Logic0_port, H(9) => X_Logic0_port, H(8) => 
                           X_Logic0_port, H(7) => X_Logic0_port, H(6) => 
                           X_Logic0_port, H(5) => X_Logic0_port, H(4) => 
                           X_Logic0_port, H(3) => X_Logic0_port, H(2) => 
                           X_Logic0_port, H(1) => X_Logic0_port, H(0) => 
                           X_Logic0_port, S(2) => Bo_signal_2_port, S(1) => 
                           Bo_signal_1_port, S(0) => Bo_signal_0_port, Y(31) =>
                           aEncMatrix_0_31_port, Y(30) => aEncMatrix_0_30_port,
                           Y(29) => aEncMatrix_0_29_port, Y(28) => 
                           aEncMatrix_0_28_port, Y(27) => aEncMatrix_0_27_port,
                           Y(26) => aEncMatrix_0_26_port, Y(25) => 
                           aEncMatrix_0_25_port, Y(24) => aEncMatrix_0_24_port,
                           Y(23) => aEncMatrix_0_23_port, Y(22) => 
                           aEncMatrix_0_22_port, Y(21) => aEncMatrix_0_21_port,
                           Y(20) => aEncMatrix_0_20_port, Y(19) => 
                           aEncMatrix_0_19_port, Y(18) => aEncMatrix_0_18_port,
                           Y(17) => aEncMatrix_0_17_port, Y(16) => 
                           aEncMatrix_0_16_port, Y(15) => aEncMatrix_0_15_port,
                           Y(14) => aEncMatrix_0_14_port, Y(13) => 
                           aEncMatrix_0_13_port, Y(12) => aEncMatrix_0_12_port,
                           Y(11) => aEncMatrix_0_11_port, Y(10) => 
                           aEncMatrix_0_10_port, Y(9) => aEncMatrix_0_9_port, 
                           Y(8) => aEncMatrix_0_8_port, Y(7) => 
                           aEncMatrix_0_7_port, Y(6) => aEncMatrix_0_6_port, 
                           Y(5) => aEncMatrix_0_5_port, Y(4) => 
                           aEncMatrix_0_4_port, Y(3) => aEncMatrix_0_3_port, 
                           Y(2) => aEncMatrix_0_2_port, Y(1) => 
                           aEncMatrix_0_1_port, Y(0) => aEncMatrix_0_0_port);
   MUXES_1 : MUX81_N32_2 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => A(15), B(30) => A(15), B(29)
                           => A(15), B(28) => A(15), B(27) => A(15), B(26) => 
                           A(15), B(25) => A(15), B(24) => A(15), B(23) => 
                           A(15), B(22) => A(15), B(21) => A(15), B(20) => 
                           A(15), B(19) => A(15), B(18) => A(15), B(17) => 
                           A(15), B(16) => A(14), B(15) => A(13), B(14) => 
                           A(12), B(13) => A(11), B(12) => A(10), B(11) => A(9)
                           , B(10) => A(8), B(9) => A(7), B(8) => A(6), B(7) =>
                           A(5), B(6) => A(4), B(5) => A(3), B(4) => A(2), B(3)
                           => A(1), B(2) => A(0), B(1) => X_Logic0_port, B(0) 
                           => X_Logic0_port, C(31) => aMatrix_9_31_port, C(30) 
                           => aMatrix_9_31_port, C(29) => aMatrix_9_31_port, 
                           C(28) => aMatrix_9_31_port, C(27) => 
                           aMatrix_9_31_port, C(26) => aMatrix_9_31_port, C(25)
                           => aMatrix_9_31_port, C(24) => aMatrix_9_31_port, 
                           C(23) => aMatrix_9_31_port, C(22) => 
                           aMatrix_9_31_port, C(21) => aMatrix_9_31_port, C(20)
                           => aMatrix_9_31_port, C(19) => aMatrix_9_31_port, 
                           C(18) => aMatrix_9_31_port, C(17) => 
                           aMatrix_9_19_port, C(16) => aMatrix_9_18_port, C(15)
                           => aMatrix_9_17_port, C(14) => aMatrix_9_16_port, 
                           C(13) => aMatrix_9_15_port, C(12) => 
                           aMatrix_9_14_port, C(11) => aMatrix_9_13_port, C(10)
                           => aMatrix_9_12_port, C(9) => aMatrix_9_11_port, 
                           C(8) => aMatrix_9_10_port, C(7) => aMatrix_9_9_port,
                           C(6) => aMatrix_9_8_port, C(5) => aMatrix_9_7_port, 
                           C(4) => aMatrix_9_6_port, C(3) => aMatrix_9_5_port, 
                           C(2) => A(0), C(1) => n20, C(0) => aMatrix_5_0_port,
                           D(31) => A(15), D(30) => A(15), D(29) => A(15), 
                           D(28) => A(15), D(27) => A(15), D(26) => A(15), 
                           D(25) => A(15), D(24) => A(15), D(23) => A(15), 
                           D(22) => A(15), D(21) => A(15), D(20) => A(15), 
                           D(19) => A(15), D(18) => A(15), D(17) => A(14), 
                           D(16) => A(13), D(15) => A(12), D(14) => A(11), 
                           D(13) => A(10), D(12) => A(9), D(11) => A(8), D(10) 
                           => A(7), D(9) => A(6), D(8) => A(5), D(7) => A(4), 
                           D(6) => A(3), D(5) => A(2), D(4) => A(1), D(3) => 
                           A(0), D(2) => X_Logic0_port, D(1) => X_Logic0_port, 
                           D(0) => X_Logic0_port, E(31) => aMatrix_9_31_port, 
                           E(30) => aMatrix_9_31_port, E(29) => 
                           aMatrix_9_31_port, E(28) => aMatrix_9_31_port, E(27)
                           => aMatrix_9_31_port, E(26) => aMatrix_9_31_port, 
                           E(25) => aMatrix_9_31_port, E(24) => 
                           aMatrix_9_31_port, E(23) => aMatrix_9_31_port, E(22)
                           => aMatrix_9_31_port, E(21) => aMatrix_9_31_port, 
                           E(20) => aMatrix_9_31_port, E(19) => 
                           aMatrix_9_31_port, E(18) => aMatrix_9_19_port, E(17)
                           => aMatrix_9_18_port, E(16) => aMatrix_9_17_port, 
                           E(15) => aMatrix_9_16_port, E(14) => 
                           aMatrix_9_15_port, E(13) => aMatrix_9_14_port, E(12)
                           => aMatrix_9_13_port, E(11) => aMatrix_9_12_port, 
                           E(10) => aMatrix_9_11_port, E(9) => 
                           aMatrix_9_10_port, E(8) => aMatrix_9_9_port, E(7) =>
                           aMatrix_9_8_port, E(6) => aMatrix_9_7_port, E(5) => 
                           aMatrix_9_6_port, E(4) => aMatrix_9_5_port, E(3) => 
                           A(0), E(2) => n20, E(1) => n20, E(0) => 
                           aMatrix_7_0_port, F(31) => X_Logic0_port, F(30) => 
                           X_Logic0_port, F(29) => X_Logic0_port, F(28) => 
                           X_Logic0_port, F(27) => X_Logic0_port, F(26) => 
                           X_Logic0_port, F(25) => X_Logic0_port, F(24) => 
                           X_Logic0_port, F(23) => X_Logic0_port, F(22) => 
                           X_Logic0_port, F(21) => X_Logic0_port, F(20) => 
                           X_Logic0_port, F(19) => X_Logic0_port, F(18) => 
                           X_Logic0_port, F(17) => X_Logic0_port, F(16) => 
                           X_Logic0_port, F(15) => X_Logic0_port, F(14) => 
                           X_Logic0_port, F(13) => X_Logic0_port, F(12) => 
                           X_Logic0_port, F(11) => X_Logic0_port, F(10) => 
                           X_Logic0_port, F(9) => X_Logic0_port, F(8) => 
                           X_Logic0_port, F(7) => X_Logic0_port, F(6) => 
                           X_Logic0_port, F(5) => X_Logic0_port, F(4) => 
                           X_Logic0_port, F(3) => X_Logic0_port, F(2) => 
                           X_Logic0_port, F(1) => X_Logic0_port, F(0) => 
                           X_Logic0_port, G(31) => X_Logic0_port, G(30) => 
                           X_Logic0_port, G(29) => X_Logic0_port, G(28) => 
                           X_Logic0_port, G(27) => X_Logic0_port, G(26) => 
                           X_Logic0_port, G(25) => X_Logic0_port, G(24) => 
                           X_Logic0_port, G(23) => X_Logic0_port, G(22) => 
                           X_Logic0_port, G(21) => X_Logic0_port, G(20) => 
                           X_Logic0_port, G(19) => X_Logic0_port, G(18) => 
                           X_Logic0_port, G(17) => X_Logic0_port, G(16) => 
                           X_Logic0_port, G(15) => X_Logic0_port, G(14) => 
                           X_Logic0_port, G(13) => X_Logic0_port, G(12) => 
                           X_Logic0_port, G(11) => X_Logic0_port, G(10) => 
                           X_Logic0_port, G(9) => X_Logic0_port, G(8) => 
                           X_Logic0_port, G(7) => X_Logic0_port, G(6) => 
                           X_Logic0_port, G(5) => X_Logic0_port, G(4) => 
                           X_Logic0_port, G(3) => X_Logic0_port, G(2) => 
                           X_Logic0_port, G(1) => X_Logic0_port, G(0) => 
                           X_Logic0_port, H(31) => X_Logic0_port, H(30) => 
                           X_Logic0_port, H(29) => X_Logic0_port, H(28) => 
                           X_Logic0_port, H(27) => X_Logic0_port, H(26) => 
                           X_Logic0_port, H(25) => X_Logic0_port, H(24) => 
                           X_Logic0_port, H(23) => X_Logic0_port, H(22) => 
                           X_Logic0_port, H(21) => X_Logic0_port, H(20) => 
                           X_Logic0_port, H(19) => X_Logic0_port, H(18) => 
                           X_Logic0_port, H(17) => X_Logic0_port, H(16) => 
                           X_Logic0_port, H(15) => X_Logic0_port, H(14) => 
                           X_Logic0_port, H(13) => X_Logic0_port, H(12) => 
                           X_Logic0_port, H(11) => X_Logic0_port, H(10) => 
                           X_Logic0_port, H(9) => X_Logic0_port, H(8) => 
                           X_Logic0_port, H(7) => X_Logic0_port, H(6) => 
                           X_Logic0_port, H(5) => X_Logic0_port, H(4) => 
                           X_Logic0_port, H(3) => X_Logic0_port, H(2) => 
                           X_Logic0_port, H(1) => X_Logic0_port, H(0) => 
                           X_Logic0_port, S(2) => Bo_signal_5_port, S(1) => 
                           Bo_signal_4_port, S(0) => Bo_signal_3_port, Y(31) =>
                           aEncMatrix_1_31_port, Y(30) => aEncMatrix_1_30_port,
                           Y(29) => aEncMatrix_1_29_port, Y(28) => 
                           aEncMatrix_1_28_port, Y(27) => aEncMatrix_1_27_port,
                           Y(26) => aEncMatrix_1_26_port, Y(25) => 
                           aEncMatrix_1_25_port, Y(24) => aEncMatrix_1_24_port,
                           Y(23) => aEncMatrix_1_23_port, Y(22) => 
                           aEncMatrix_1_22_port, Y(21) => aEncMatrix_1_21_port,
                           Y(20) => aEncMatrix_1_20_port, Y(19) => 
                           aEncMatrix_1_19_port, Y(18) => aEncMatrix_1_18_port,
                           Y(17) => aEncMatrix_1_17_port, Y(16) => 
                           aEncMatrix_1_16_port, Y(15) => aEncMatrix_1_15_port,
                           Y(14) => aEncMatrix_1_14_port, Y(13) => 
                           aEncMatrix_1_13_port, Y(12) => aEncMatrix_1_12_port,
                           Y(11) => aEncMatrix_1_11_port, Y(10) => 
                           aEncMatrix_1_10_port, Y(9) => aEncMatrix_1_9_port, 
                           Y(8) => aEncMatrix_1_8_port, Y(7) => 
                           aEncMatrix_1_7_port, Y(6) => aEncMatrix_1_6_port, 
                           Y(5) => aEncMatrix_1_5_port, Y(4) => 
                           aEncMatrix_1_4_port, Y(3) => aEncMatrix_1_3_port, 
                           Y(2) => aEncMatrix_1_2_port, Y(1) => 
                           aEncMatrix_1_1_port, Y(0) => aEncMatrix_1_0_port);
   FIRST_RCA_1 : RCA_N32_2 port map( A(31) => aEncMatrix_1_31_port, A(30) => 
                           aEncMatrix_1_30_port, A(29) => aEncMatrix_1_29_port,
                           A(28) => aEncMatrix_1_28_port, A(27) => 
                           aEncMatrix_1_27_port, A(26) => aEncMatrix_1_26_port,
                           A(25) => aEncMatrix_1_25_port, A(24) => 
                           aEncMatrix_1_24_port, A(23) => aEncMatrix_1_23_port,
                           A(22) => aEncMatrix_1_22_port, A(21) => 
                           aEncMatrix_1_21_port, A(20) => aEncMatrix_1_20_port,
                           A(19) => aEncMatrix_1_19_port, A(18) => 
                           aEncMatrix_1_18_port, A(17) => aEncMatrix_1_17_port,
                           A(16) => aEncMatrix_1_16_port, A(15) => 
                           aEncMatrix_1_15_port, A(14) => aEncMatrix_1_14_port,
                           A(13) => aEncMatrix_1_13_port, A(12) => 
                           aEncMatrix_1_12_port, A(11) => aEncMatrix_1_11_port,
                           A(10) => aEncMatrix_1_10_port, A(9) => 
                           aEncMatrix_1_9_port, A(8) => aEncMatrix_1_8_port, 
                           A(7) => aEncMatrix_1_7_port, A(6) => 
                           aEncMatrix_1_6_port, A(5) => aEncMatrix_1_5_port, 
                           A(4) => aEncMatrix_1_4_port, A(3) => 
                           aEncMatrix_1_3_port, A(2) => aEncMatrix_1_2_port, 
                           A(1) => aEncMatrix_1_1_port, A(0) => 
                           aEncMatrix_1_0_port, B(31) => aEncMatrix_0_31_port, 
                           B(30) => aEncMatrix_0_30_port, B(29) => 
                           aEncMatrix_0_29_port, B(28) => aEncMatrix_0_28_port,
                           B(27) => aEncMatrix_0_27_port, B(26) => 
                           aEncMatrix_0_26_port, B(25) => aEncMatrix_0_25_port,
                           B(24) => aEncMatrix_0_24_port, B(23) => 
                           aEncMatrix_0_23_port, B(22) => aEncMatrix_0_22_port,
                           B(21) => aEncMatrix_0_21_port, B(20) => 
                           aEncMatrix_0_20_port, B(19) => aEncMatrix_0_19_port,
                           B(18) => aEncMatrix_0_18_port, B(17) => 
                           aEncMatrix_0_17_port, B(16) => aEncMatrix_0_16_port,
                           B(15) => aEncMatrix_0_15_port, B(14) => 
                           aEncMatrix_0_14_port, B(13) => aEncMatrix_0_13_port,
                           B(12) => aEncMatrix_0_12_port, B(11) => 
                           aEncMatrix_0_11_port, B(10) => aEncMatrix_0_10_port,
                           B(9) => aEncMatrix_0_9_port, B(8) => 
                           aEncMatrix_0_8_port, B(7) => aEncMatrix_0_7_port, 
                           B(6) => aEncMatrix_0_6_port, B(5) => 
                           aEncMatrix_0_5_port, B(4) => aEncMatrix_0_4_port, 
                           B(3) => aEncMatrix_0_3_port, B(2) => 
                           aEncMatrix_0_2_port, B(1) => aEncMatrix_0_1_port, 
                           B(0) => aEncMatrix_0_0_port, Ci => X_Logic0_port, 
                           S(31) => pSumMatrix_0_31_port, S(30) => 
                           pSumMatrix_0_30_port, S(29) => pSumMatrix_0_29_port,
                           S(28) => pSumMatrix_0_28_port, S(27) => 
                           pSumMatrix_0_27_port, S(26) => pSumMatrix_0_26_port,
                           S(25) => pSumMatrix_0_25_port, S(24) => 
                           pSumMatrix_0_24_port, S(23) => pSumMatrix_0_23_port,
                           S(22) => pSumMatrix_0_22_port, S(21) => 
                           pSumMatrix_0_21_port, S(20) => pSumMatrix_0_20_port,
                           S(19) => pSumMatrix_0_19_port, S(18) => 
                           pSumMatrix_0_18_port, S(17) => pSumMatrix_0_17_port,
                           S(16) => pSumMatrix_0_16_port, S(15) => 
                           pSumMatrix_0_15_port, S(14) => pSumMatrix_0_14_port,
                           S(13) => pSumMatrix_0_13_port, S(12) => 
                           pSumMatrix_0_12_port, S(11) => pSumMatrix_0_11_port,
                           S(10) => pSumMatrix_0_10_port, S(9) => 
                           pSumMatrix_0_9_port, S(8) => pSumMatrix_0_8_port, 
                           S(7) => pSumMatrix_0_7_port, S(6) => 
                           pSumMatrix_0_6_port, S(5) => pSumMatrix_0_5_port, 
                           S(4) => pSumMatrix_0_4_port, S(3) => 
                           pSumMatrix_0_3_port, S(2) => pSumMatrix_0_2_port, 
                           S(1) => pSumMatrix_0_1_port, S(0) => 
                           pSumMatrix_0_0_port, Co => n_1280);
   MUXES_2 : MUX81_N32_1 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => A(15), B(30) => A(15), B(29)
                           => A(15), B(28) => A(15), B(27) => A(15), B(26) => 
                           A(15), B(25) => A(15), B(24) => A(15), B(23) => 
                           A(15), B(22) => A(15), B(21) => A(15), B(20) => 
                           A(15), B(19) => A(15), B(18) => A(14), B(17) => 
                           A(13), B(16) => A(12), B(15) => A(11), B(14) => 
                           A(10), B(13) => A(9), B(12) => A(8), B(11) => A(7), 
                           B(10) => A(6), B(9) => A(5), B(8) => A(4), B(7) => 
                           A(3), B(6) => A(2), B(5) => A(1), B(4) => A(0), B(3)
                           => X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(31) => 
                           aMatrix_9_31_port, C(30) => aMatrix_9_31_port, C(29)
                           => aMatrix_9_31_port, C(28) => aMatrix_9_31_port, 
                           C(27) => aMatrix_9_31_port, C(26) => 
                           aMatrix_9_31_port, C(25) => aMatrix_9_31_port, C(24)
                           => aMatrix_9_31_port, C(23) => aMatrix_9_31_port, 
                           C(22) => aMatrix_9_31_port, C(21) => 
                           aMatrix_9_31_port, C(20) => aMatrix_9_31_port, C(19)
                           => aMatrix_9_19_port, C(18) => aMatrix_9_18_port, 
                           C(17) => aMatrix_9_17_port, C(16) => 
                           aMatrix_9_16_port, C(15) => aMatrix_9_15_port, C(14)
                           => aMatrix_9_14_port, C(13) => aMatrix_9_13_port, 
                           C(12) => aMatrix_9_12_port, C(11) => 
                           aMatrix_9_11_port, C(10) => aMatrix_9_10_port, C(9) 
                           => aMatrix_9_9_port, C(8) => aMatrix_9_8_port, C(7) 
                           => aMatrix_9_7_port, C(6) => aMatrix_9_6_port, C(5) 
                           => aMatrix_9_5_port, C(4) => A(0), C(3) => n20, C(2)
                           => n20, C(1) => n20, C(0) => aMatrix_9_0_port, D(31)
                           => A(15), D(30) => A(15), D(29) => A(15), D(28) => 
                           A(15), D(27) => A(15), D(26) => A(15), D(25) => 
                           A(15), D(24) => A(15), D(23) => A(15), D(22) => 
                           A(15), D(21) => A(15), D(20) => A(15), D(19) => 
                           A(14), D(18) => A(13), D(17) => A(12), D(16) => 
                           A(11), D(15) => A(10), D(14) => A(9), D(13) => A(8),
                           D(12) => A(7), D(11) => A(6), D(10) => A(5), D(9) =>
                           A(4), D(8) => A(3), D(7) => A(2), D(6) => A(1), D(5)
                           => A(0), D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, E(31) => 
                           aMatrix_9_31_port, E(30) => aMatrix_9_31_port, E(29)
                           => aMatrix_9_31_port, E(28) => aMatrix_9_31_port, 
                           E(27) => aMatrix_9_31_port, E(26) => 
                           aMatrix_9_31_port, E(25) => aMatrix_9_31_port, E(24)
                           => aMatrix_9_31_port, E(23) => aMatrix_9_31_port, 
                           E(22) => aMatrix_9_31_port, E(21) => 
                           aMatrix_9_31_port, E(20) => aMatrix_9_19_port, E(19)
                           => aMatrix_9_18_port, E(18) => aMatrix_9_17_port, 
                           E(17) => aMatrix_9_16_port, E(16) => 
                           aMatrix_9_15_port, E(15) => aMatrix_9_14_port, E(14)
                           => aMatrix_9_13_port, E(13) => aMatrix_9_12_port, 
                           E(12) => aMatrix_9_11_port, E(11) => 
                           aMatrix_9_10_port, E(10) => aMatrix_9_9_port, E(9) 
                           => aMatrix_9_8_port, E(8) => aMatrix_9_7_port, E(7) 
                           => aMatrix_9_6_port, E(6) => aMatrix_9_5_port, E(5) 
                           => A(0), E(4) => n20, E(3) => n20, E(2) => n20, E(1)
                           => n20, E(0) => aMatrix_11_0_port, F(31) => 
                           X_Logic0_port, F(30) => X_Logic0_port, F(29) => 
                           X_Logic0_port, F(28) => X_Logic0_port, F(27) => 
                           X_Logic0_port, F(26) => X_Logic0_port, F(25) => 
                           X_Logic0_port, F(24) => X_Logic0_port, F(23) => 
                           X_Logic0_port, F(22) => X_Logic0_port, F(21) => 
                           X_Logic0_port, F(20) => X_Logic0_port, F(19) => 
                           X_Logic0_port, F(18) => X_Logic0_port, F(17) => 
                           X_Logic0_port, F(16) => X_Logic0_port, F(15) => 
                           X_Logic0_port, F(14) => X_Logic0_port, F(13) => 
                           X_Logic0_port, F(12) => X_Logic0_port, F(11) => 
                           X_Logic0_port, F(10) => X_Logic0_port, F(9) => 
                           X_Logic0_port, F(8) => X_Logic0_port, F(7) => 
                           X_Logic0_port, F(6) => X_Logic0_port, F(5) => 
                           X_Logic0_port, F(4) => X_Logic0_port, F(3) => 
                           X_Logic0_port, F(2) => X_Logic0_port, F(1) => 
                           X_Logic0_port, F(0) => X_Logic0_port, G(31) => 
                           X_Logic0_port, G(30) => X_Logic0_port, G(29) => 
                           X_Logic0_port, G(28) => X_Logic0_port, G(27) => 
                           X_Logic0_port, G(26) => X_Logic0_port, G(25) => 
                           X_Logic0_port, G(24) => X_Logic0_port, G(23) => 
                           X_Logic0_port, G(22) => X_Logic0_port, G(21) => 
                           X_Logic0_port, G(20) => X_Logic0_port, G(19) => 
                           X_Logic0_port, G(18) => X_Logic0_port, G(17) => 
                           X_Logic0_port, G(16) => X_Logic0_port, G(15) => 
                           X_Logic0_port, G(14) => X_Logic0_port, G(13) => 
                           X_Logic0_port, G(12) => X_Logic0_port, G(11) => 
                           X_Logic0_port, G(10) => X_Logic0_port, G(9) => 
                           X_Logic0_port, G(8) => X_Logic0_port, G(7) => 
                           X_Logic0_port, G(6) => X_Logic0_port, G(5) => 
                           X_Logic0_port, G(4) => X_Logic0_port, G(3) => 
                           X_Logic0_port, G(2) => X_Logic0_port, G(1) => 
                           X_Logic0_port, G(0) => X_Logic0_port, H(31) => 
                           X_Logic0_port, H(30) => X_Logic0_port, H(29) => 
                           X_Logic0_port, H(28) => X_Logic0_port, H(27) => 
                           X_Logic0_port, H(26) => X_Logic0_port, H(25) => 
                           X_Logic0_port, H(24) => X_Logic0_port, H(23) => 
                           X_Logic0_port, H(22) => X_Logic0_port, H(21) => 
                           X_Logic0_port, H(20) => X_Logic0_port, H(19) => 
                           X_Logic0_port, H(18) => X_Logic0_port, H(17) => 
                           X_Logic0_port, H(16) => X_Logic0_port, H(15) => 
                           X_Logic0_port, H(14) => X_Logic0_port, H(13) => 
                           X_Logic0_port, H(12) => X_Logic0_port, H(11) => 
                           X_Logic0_port, H(10) => X_Logic0_port, H(9) => 
                           X_Logic0_port, H(8) => X_Logic0_port, H(7) => 
                           X_Logic0_port, H(6) => X_Logic0_port, H(5) => 
                           X_Logic0_port, H(4) => X_Logic0_port, H(3) => 
                           X_Logic0_port, H(2) => X_Logic0_port, H(1) => 
                           X_Logic0_port, H(0) => X_Logic0_port, S(2) => 
                           Bo_signal_8_port, S(1) => Bo_signal_7_port, S(0) => 
                           Bo_signal_6_port, Y(31) => aEncMatrix_2_31_port, 
                           Y(30) => aEncMatrix_2_30_port, Y(29) => 
                           aEncMatrix_2_29_port, Y(28) => aEncMatrix_2_28_port,
                           Y(27) => aEncMatrix_2_27_port, Y(26) => 
                           aEncMatrix_2_26_port, Y(25) => aEncMatrix_2_25_port,
                           Y(24) => aEncMatrix_2_24_port, Y(23) => 
                           aEncMatrix_2_23_port, Y(22) => aEncMatrix_2_22_port,
                           Y(21) => aEncMatrix_2_21_port, Y(20) => 
                           aEncMatrix_2_20_port, Y(19) => aEncMatrix_2_19_port,
                           Y(18) => aEncMatrix_2_18_port, Y(17) => 
                           aEncMatrix_2_17_port, Y(16) => aEncMatrix_2_16_port,
                           Y(15) => aEncMatrix_2_15_port, Y(14) => 
                           aEncMatrix_2_14_port, Y(13) => aEncMatrix_2_13_port,
                           Y(12) => aEncMatrix_2_12_port, Y(11) => 
                           aEncMatrix_2_11_port, Y(10) => aEncMatrix_2_10_port,
                           Y(9) => aEncMatrix_2_9_port, Y(8) => 
                           aEncMatrix_2_8_port, Y(7) => aEncMatrix_2_7_port, 
                           Y(6) => aEncMatrix_2_6_port, Y(5) => 
                           aEncMatrix_2_5_port, Y(4) => aEncMatrix_2_4_port, 
                           Y(3) => aEncMatrix_2_3_port, Y(2) => 
                           aEncMatrix_2_2_port, Y(1) => aEncMatrix_2_1_port, 
                           Y(0) => aEncMatrix_2_0_port);
   RCAS_2 : RCA_N32_1 port map( A(31) => aEncMatrix_2_31_port, A(30) => 
                           aEncMatrix_2_30_port, A(29) => aEncMatrix_2_29_port,
                           A(28) => aEncMatrix_2_28_port, A(27) => 
                           aEncMatrix_2_27_port, A(26) => aEncMatrix_2_26_port,
                           A(25) => aEncMatrix_2_25_port, A(24) => 
                           aEncMatrix_2_24_port, A(23) => aEncMatrix_2_23_port,
                           A(22) => aEncMatrix_2_22_port, A(21) => 
                           aEncMatrix_2_21_port, A(20) => aEncMatrix_2_20_port,
                           A(19) => aEncMatrix_2_19_port, A(18) => 
                           aEncMatrix_2_18_port, A(17) => aEncMatrix_2_17_port,
                           A(16) => aEncMatrix_2_16_port, A(15) => 
                           aEncMatrix_2_15_port, A(14) => aEncMatrix_2_14_port,
                           A(13) => aEncMatrix_2_13_port, A(12) => 
                           aEncMatrix_2_12_port, A(11) => aEncMatrix_2_11_port,
                           A(10) => aEncMatrix_2_10_port, A(9) => 
                           aEncMatrix_2_9_port, A(8) => aEncMatrix_2_8_port, 
                           A(7) => aEncMatrix_2_7_port, A(6) => 
                           aEncMatrix_2_6_port, A(5) => aEncMatrix_2_5_port, 
                           A(4) => aEncMatrix_2_4_port, A(3) => 
                           aEncMatrix_2_3_port, A(2) => aEncMatrix_2_2_port, 
                           A(1) => aEncMatrix_2_1_port, A(0) => 
                           aEncMatrix_2_0_port, B(31) => pSumMatrix_0_31_port, 
                           B(30) => pSumMatrix_0_30_port, B(29) => 
                           pSumMatrix_0_29_port, B(28) => pSumMatrix_0_28_port,
                           B(27) => pSumMatrix_0_27_port, B(26) => 
                           pSumMatrix_0_26_port, B(25) => pSumMatrix_0_25_port,
                           B(24) => pSumMatrix_0_24_port, B(23) => 
                           pSumMatrix_0_23_port, B(22) => pSumMatrix_0_22_port,
                           B(21) => pSumMatrix_0_21_port, B(20) => 
                           pSumMatrix_0_20_port, B(19) => pSumMatrix_0_19_port,
                           B(18) => pSumMatrix_0_18_port, B(17) => 
                           pSumMatrix_0_17_port, B(16) => pSumMatrix_0_16_port,
                           B(15) => pSumMatrix_0_15_port, B(14) => 
                           pSumMatrix_0_14_port, B(13) => pSumMatrix_0_13_port,
                           B(12) => pSumMatrix_0_12_port, B(11) => 
                           pSumMatrix_0_11_port, B(10) => pSumMatrix_0_10_port,
                           B(9) => pSumMatrix_0_9_port, B(8) => 
                           pSumMatrix_0_8_port, B(7) => pSumMatrix_0_7_port, 
                           B(6) => pSumMatrix_0_6_port, B(5) => 
                           pSumMatrix_0_5_port, B(4) => pSumMatrix_0_4_port, 
                           B(3) => pSumMatrix_0_3_port, B(2) => 
                           pSumMatrix_0_2_port, B(1) => pSumMatrix_0_1_port, 
                           B(0) => pSumMatrix_0_0_port, Ci => X_Logic0_port, 
                           S(31) => pSumMatrix_1_31_port, S(30) => 
                           pSumMatrix_1_30_port, S(29) => pSumMatrix_1_29_port,
                           S(28) => pSumMatrix_1_28_port, S(27) => 
                           pSumMatrix_1_27_port, S(26) => pSumMatrix_1_26_port,
                           S(25) => pSumMatrix_1_25_port, S(24) => 
                           pSumMatrix_1_24_port, S(23) => pSumMatrix_1_23_port,
                           S(22) => pSumMatrix_1_22_port, S(21) => 
                           pSumMatrix_1_21_port, S(20) => pSumMatrix_1_20_port,
                           S(19) => pSumMatrix_1_19_port, S(18) => 
                           pSumMatrix_1_18_port, S(17) => pSumMatrix_1_17_port,
                           S(16) => pSumMatrix_1_16_port, S(15) => 
                           pSumMatrix_1_15_port, S(14) => pSumMatrix_1_14_port,
                           S(13) => pSumMatrix_1_13_port, S(12) => 
                           pSumMatrix_1_12_port, S(11) => pSumMatrix_1_11_port,
                           S(10) => pSumMatrix_1_10_port, S(9) => 
                           pSumMatrix_1_9_port, S(8) => pSumMatrix_1_8_port, 
                           S(7) => pSumMatrix_1_7_port, S(6) => 
                           pSumMatrix_1_6_port, S(5) => pSumMatrix_1_5_port, 
                           S(4) => pSumMatrix_1_4_port, S(3) => 
                           pSumMatrix_1_3_port, S(2) => pSumMatrix_1_2_port, 
                           S(1) => pSumMatrix_1_1_port, S(0) => 
                           pSumMatrix_1_0_port, Co => n_1281);
   MUXES_3 : MUX81_N32_0 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => A(15), B(30) => A(15), B(29)
                           => A(15), B(28) => A(15), B(27) => A(15), B(26) => 
                           A(15), B(25) => A(15), B(24) => A(15), B(23) => 
                           A(15), B(22) => A(15), B(21) => A(15), B(20) => 
                           A(14), B(19) => A(13), B(18) => A(12), B(17) => 
                           A(11), B(16) => A(10), B(15) => A(9), B(14) => A(8),
                           B(13) => A(7), B(12) => A(6), B(11) => A(5), B(10) 
                           => A(4), B(9) => A(3), B(8) => A(2), B(7) => A(1), 
                           B(6) => A(0), B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, C(31) => aMatrix_9_31_port, C(30) => 
                           aMatrix_9_31_port, C(29) => aMatrix_9_31_port, C(28)
                           => aMatrix_9_31_port, C(27) => aMatrix_9_31_port, 
                           C(26) => aMatrix_9_31_port, C(25) => 
                           aMatrix_9_31_port, C(24) => aMatrix_9_31_port, C(23)
                           => aMatrix_9_31_port, C(22) => aMatrix_9_31_port, 
                           C(21) => aMatrix_9_19_port, C(20) => 
                           aMatrix_9_18_port, C(19) => aMatrix_9_17_port, C(18)
                           => aMatrix_9_16_port, C(17) => aMatrix_9_15_port, 
                           C(16) => aMatrix_9_14_port, C(15) => 
                           aMatrix_9_13_port, C(14) => aMatrix_9_12_port, C(13)
                           => aMatrix_9_11_port, C(12) => aMatrix_9_10_port, 
                           C(11) => aMatrix_9_9_port, C(10) => aMatrix_9_8_port
                           , C(9) => aMatrix_9_7_port, C(8) => aMatrix_9_6_port
                           , C(7) => aMatrix_9_5_port, C(6) => A(0), C(5) => 
                           n20, C(4) => n20, C(3) => n20, C(2) => n20, C(1) => 
                           n20, C(0) => aMatrix_13_0_port, D(31) => A(15), 
                           D(30) => A(15), D(29) => A(15), D(28) => A(15), 
                           D(27) => A(15), D(26) => A(15), D(25) => A(15), 
                           D(24) => A(15), D(23) => A(15), D(22) => A(15), 
                           D(21) => A(14), D(20) => A(13), D(19) => A(12), 
                           D(18) => A(11), D(17) => A(10), D(16) => A(9), D(15)
                           => A(8), D(14) => A(7), D(13) => A(6), D(12) => A(5)
                           , D(11) => A(4), D(10) => A(3), D(9) => A(2), D(8) 
                           => A(1), D(7) => A(0), D(6) => X_Logic0_port, D(5) 
                           => X_Logic0_port, D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, E(31) => 
                           aMatrix_9_31_port, E(30) => aMatrix_9_31_port, E(29)
                           => aMatrix_9_31_port, E(28) => aMatrix_9_31_port, 
                           E(27) => aMatrix_9_31_port, E(26) => 
                           aMatrix_9_31_port, E(25) => aMatrix_9_31_port, E(24)
                           => aMatrix_9_31_port, E(23) => aMatrix_9_31_port, 
                           E(22) => aMatrix_9_19_port, E(21) => 
                           aMatrix_9_18_port, E(20) => aMatrix_9_17_port, E(19)
                           => aMatrix_9_16_port, E(18) => aMatrix_9_15_port, 
                           E(17) => aMatrix_9_14_port, E(16) => 
                           aMatrix_9_13_port, E(15) => aMatrix_9_12_port, E(14)
                           => aMatrix_9_11_port, E(13) => aMatrix_9_10_port, 
                           E(12) => aMatrix_9_9_port, E(11) => aMatrix_9_8_port
                           , E(10) => aMatrix_9_7_port, E(9) => 
                           aMatrix_9_6_port, E(8) => aMatrix_9_5_port, E(7) => 
                           A(0), E(6) => n20, E(5) => n20, E(4) => n20, E(3) =>
                           n20, E(2) => n20, E(1) => n20, E(0) => 
                           aMatrix_15_0_port, F(31) => X_Logic0_port, F(30) => 
                           X_Logic0_port, F(29) => X_Logic0_port, F(28) => 
                           X_Logic0_port, F(27) => X_Logic0_port, F(26) => 
                           X_Logic0_port, F(25) => X_Logic0_port, F(24) => 
                           X_Logic0_port, F(23) => X_Logic0_port, F(22) => 
                           X_Logic0_port, F(21) => X_Logic0_port, F(20) => 
                           X_Logic0_port, F(19) => X_Logic0_port, F(18) => 
                           X_Logic0_port, F(17) => X_Logic0_port, F(16) => 
                           X_Logic0_port, F(15) => X_Logic0_port, F(14) => 
                           X_Logic0_port, F(13) => X_Logic0_port, F(12) => 
                           X_Logic0_port, F(11) => X_Logic0_port, F(10) => 
                           X_Logic0_port, F(9) => X_Logic0_port, F(8) => 
                           X_Logic0_port, F(7) => X_Logic0_port, F(6) => 
                           X_Logic0_port, F(5) => X_Logic0_port, F(4) => 
                           X_Logic0_port, F(3) => X_Logic0_port, F(2) => 
                           X_Logic0_port, F(1) => X_Logic0_port, F(0) => 
                           X_Logic0_port, G(31) => X_Logic0_port, G(30) => 
                           X_Logic0_port, G(29) => X_Logic0_port, G(28) => 
                           X_Logic0_port, G(27) => X_Logic0_port, G(26) => 
                           X_Logic0_port, G(25) => X_Logic0_port, G(24) => 
                           X_Logic0_port, G(23) => X_Logic0_port, G(22) => 
                           X_Logic0_port, G(21) => X_Logic0_port, G(20) => 
                           X_Logic0_port, G(19) => X_Logic0_port, G(18) => 
                           X_Logic0_port, G(17) => X_Logic0_port, G(16) => 
                           X_Logic0_port, G(15) => X_Logic0_port, G(14) => 
                           X_Logic0_port, G(13) => X_Logic0_port, G(12) => 
                           X_Logic0_port, G(11) => X_Logic0_port, G(10) => 
                           X_Logic0_port, G(9) => X_Logic0_port, G(8) => 
                           X_Logic0_port, G(7) => X_Logic0_port, G(6) => 
                           X_Logic0_port, G(5) => X_Logic0_port, G(4) => 
                           X_Logic0_port, G(3) => X_Logic0_port, G(2) => 
                           X_Logic0_port, G(1) => X_Logic0_port, G(0) => 
                           X_Logic0_port, H(31) => X_Logic0_port, H(30) => 
                           X_Logic0_port, H(29) => X_Logic0_port, H(28) => 
                           X_Logic0_port, H(27) => X_Logic0_port, H(26) => 
                           X_Logic0_port, H(25) => X_Logic0_port, H(24) => 
                           X_Logic0_port, H(23) => X_Logic0_port, H(22) => 
                           X_Logic0_port, H(21) => X_Logic0_port, H(20) => 
                           X_Logic0_port, H(19) => X_Logic0_port, H(18) => 
                           X_Logic0_port, H(17) => X_Logic0_port, H(16) => 
                           X_Logic0_port, H(15) => X_Logic0_port, H(14) => 
                           X_Logic0_port, H(13) => X_Logic0_port, H(12) => 
                           X_Logic0_port, H(11) => X_Logic0_port, H(10) => 
                           X_Logic0_port, H(9) => X_Logic0_port, H(8) => 
                           X_Logic0_port, H(7) => X_Logic0_port, H(6) => 
                           X_Logic0_port, H(5) => X_Logic0_port, H(4) => 
                           X_Logic0_port, H(3) => X_Logic0_port, H(2) => 
                           X_Logic0_port, H(1) => X_Logic0_port, H(0) => 
                           X_Logic0_port, S(2) => Bo_signal_11_port, S(1) => 
                           Bo_signal_10_port, S(0) => Bo_signal_9_port, Y(31) 
                           => aEncMatrix_3_31_port, Y(30) => 
                           aEncMatrix_3_30_port, Y(29) => aEncMatrix_3_29_port,
                           Y(28) => aEncMatrix_3_28_port, Y(27) => 
                           aEncMatrix_3_27_port, Y(26) => aEncMatrix_3_26_port,
                           Y(25) => aEncMatrix_3_25_port, Y(24) => 
                           aEncMatrix_3_24_port, Y(23) => aEncMatrix_3_23_port,
                           Y(22) => aEncMatrix_3_22_port, Y(21) => 
                           aEncMatrix_3_21_port, Y(20) => aEncMatrix_3_20_port,
                           Y(19) => aEncMatrix_3_19_port, Y(18) => 
                           aEncMatrix_3_18_port, Y(17) => aEncMatrix_3_17_port,
                           Y(16) => aEncMatrix_3_16_port, Y(15) => 
                           aEncMatrix_3_15_port, Y(14) => aEncMatrix_3_14_port,
                           Y(13) => aEncMatrix_3_13_port, Y(12) => 
                           aEncMatrix_3_12_port, Y(11) => aEncMatrix_3_11_port,
                           Y(10) => aEncMatrix_3_10_port, Y(9) => 
                           aEncMatrix_3_9_port, Y(8) => aEncMatrix_3_8_port, 
                           Y(7) => aEncMatrix_3_7_port, Y(6) => 
                           aEncMatrix_3_6_port, Y(5) => aEncMatrix_3_5_port, 
                           Y(4) => aEncMatrix_3_4_port, Y(3) => 
                           aEncMatrix_3_3_port, Y(2) => aEncMatrix_3_2_port, 
                           Y(1) => aEncMatrix_3_1_port, Y(0) => 
                           aEncMatrix_3_0_port);
   RCAS_3 : RCA_N32_0 port map( A(31) => aEncMatrix_3_31_port, A(30) => 
                           aEncMatrix_3_30_port, A(29) => aEncMatrix_3_29_port,
                           A(28) => aEncMatrix_3_28_port, A(27) => 
                           aEncMatrix_3_27_port, A(26) => aEncMatrix_3_26_port,
                           A(25) => aEncMatrix_3_25_port, A(24) => 
                           aEncMatrix_3_24_port, A(23) => aEncMatrix_3_23_port,
                           A(22) => aEncMatrix_3_22_port, A(21) => 
                           aEncMatrix_3_21_port, A(20) => aEncMatrix_3_20_port,
                           A(19) => aEncMatrix_3_19_port, A(18) => 
                           aEncMatrix_3_18_port, A(17) => aEncMatrix_3_17_port,
                           A(16) => aEncMatrix_3_16_port, A(15) => 
                           aEncMatrix_3_15_port, A(14) => aEncMatrix_3_14_port,
                           A(13) => aEncMatrix_3_13_port, A(12) => 
                           aEncMatrix_3_12_port, A(11) => aEncMatrix_3_11_port,
                           A(10) => aEncMatrix_3_10_port, A(9) => 
                           aEncMatrix_3_9_port, A(8) => aEncMatrix_3_8_port, 
                           A(7) => aEncMatrix_3_7_port, A(6) => 
                           aEncMatrix_3_6_port, A(5) => aEncMatrix_3_5_port, 
                           A(4) => aEncMatrix_3_4_port, A(3) => 
                           aEncMatrix_3_3_port, A(2) => aEncMatrix_3_2_port, 
                           A(1) => aEncMatrix_3_1_port, A(0) => 
                           aEncMatrix_3_0_port, B(31) => pSumMatrix_1_31_port, 
                           B(30) => pSumMatrix_1_30_port, B(29) => 
                           pSumMatrix_1_29_port, B(28) => pSumMatrix_1_28_port,
                           B(27) => pSumMatrix_1_27_port, B(26) => 
                           pSumMatrix_1_26_port, B(25) => pSumMatrix_1_25_port,
                           B(24) => pSumMatrix_1_24_port, B(23) => 
                           pSumMatrix_1_23_port, B(22) => pSumMatrix_1_22_port,
                           B(21) => pSumMatrix_1_21_port, B(20) => 
                           pSumMatrix_1_20_port, B(19) => pSumMatrix_1_19_port,
                           B(18) => pSumMatrix_1_18_port, B(17) => 
                           pSumMatrix_1_17_port, B(16) => pSumMatrix_1_16_port,
                           B(15) => pSumMatrix_1_15_port, B(14) => 
                           pSumMatrix_1_14_port, B(13) => pSumMatrix_1_13_port,
                           B(12) => pSumMatrix_1_12_port, B(11) => 
                           pSumMatrix_1_11_port, B(10) => pSumMatrix_1_10_port,
                           B(9) => pSumMatrix_1_9_port, B(8) => 
                           pSumMatrix_1_8_port, B(7) => pSumMatrix_1_7_port, 
                           B(6) => pSumMatrix_1_6_port, B(5) => 
                           pSumMatrix_1_5_port, B(4) => pSumMatrix_1_4_port, 
                           B(3) => pSumMatrix_1_3_port, B(2) => 
                           pSumMatrix_1_2_port, B(1) => pSumMatrix_1_1_port, 
                           B(0) => pSumMatrix_1_0_port, Ci => X_Logic0_port, 
                           S(31) => P(31), S(30) => P(30), S(29) => P(29), 
                           S(28) => P(28), S(27) => P(27), S(26) => P(26), 
                           S(25) => P(25), S(24) => P(24), S(23) => P(23), 
                           S(22) => P(22), S(21) => P(21), S(20) => P(20), 
                           S(19) => P(19), S(18) => P(18), S(17) => P(17), 
                           S(16) => P(16), S(15) => P(15), S(14) => P(14), 
                           S(13) => P(13), S(12) => P(12), S(11) => P(11), 
                           S(10) => P(10), S(9) => P(9), S(8) => P(8), S(7) => 
                           P(7), S(6) => P(6), S(5) => P(5), S(4) => P(4), S(3)
                           => P(3), S(2) => P(2), S(1) => P(1), S(0) => P(0), 
                           Co => n_1282);
   U3 : INV_X8 port map( A => n4, ZN => aMatrix_9_31_port);
   U4 : XOR2_X1 port map( A => n1, B => A(4), Z => aMatrix_9_8_port);
   U5 : OR2_X1 port map( A1 => n2, A2 => A(3), ZN => n1);
   U6 : XOR2_X1 port map( A => n2, B => A(3), Z => aMatrix_9_7_port);
   U7 : XNOR2_X1 port map( A => A(2), B => n3, ZN => aMatrix_9_6_port);
   U8 : NOR2_X1 port map( A1 => A(0), A2 => A(1), ZN => n3);
   U9 : XOR2_X1 port map( A => A(1), B => A(0), Z => aMatrix_9_5_port);
   U10 : OAI21_X1 port map( B1 => n5, B2 => n6, A => n4, ZN => 
                           aMatrix_9_19_port);
   U11 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => n4);
   U12 : INV_X1 port map( A => A(15), ZN => n6);
   U13 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => n5);
   U14 : INV_X1 port map( A => A(14), ZN => n8);
   U15 : MUX2_X1 port map( A => n9, B => n7, S => A(14), Z => aMatrix_9_18_port
                           );
   U16 : NOR2_X1 port map( A1 => n10, A2 => A(13), ZN => n7);
   U17 : OR2_X1 port map( A1 => A(13), A2 => n10, ZN => n9);
   U18 : XOR2_X1 port map( A => n10, B => A(13), Z => aMatrix_9_17_port);
   U19 : OR3_X1 port map( A1 => A(11), A2 => A(12), A3 => n11, ZN => n10);
   U20 : XOR2_X1 port map( A => n12, B => A(12), Z => aMatrix_9_16_port);
   U21 : OR2_X1 port map( A1 => n11, A2 => A(11), ZN => n12);
   U22 : XOR2_X1 port map( A => n11, B => A(11), Z => aMatrix_9_15_port);
   U23 : OR2_X1 port map( A1 => n13, A2 => A(10), ZN => n11);
   U24 : XOR2_X1 port map( A => n13, B => A(10), Z => aMatrix_9_14_port);
   U25 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U26 : INV_X1 port map( A => A(9), ZN => n15);
   U27 : XNOR2_X1 port map( A => n14, B => A(9), ZN => aMatrix_9_13_port);
   U28 : NOR3_X1 port map( A1 => A(7), A2 => A(8), A3 => n16, ZN => n14);
   U29 : XOR2_X1 port map( A => n17, B => A(8), Z => aMatrix_9_12_port);
   U30 : OR2_X1 port map( A1 => n16, A2 => A(7), ZN => n17);
   U31 : XOR2_X1 port map( A => n16, B => A(7), Z => aMatrix_9_11_port);
   U32 : OR3_X1 port map( A1 => A(5), A2 => A(6), A3 => n18, ZN => n16);
   U33 : XOR2_X1 port map( A => n19, B => A(6), Z => aMatrix_9_10_port);
   U34 : OR2_X1 port map( A1 => n18, A2 => A(5), ZN => n19);
   U35 : XOR2_X1 port map( A => n18, B => A(5), Z => aMatrix_9_9_port);
   U36 : OR3_X1 port map( A1 => A(3), A2 => A(4), A3 => n2, ZN => n18);
   U37 : OR3_X1 port map( A1 => A(1), A2 => A(2), A3 => A(0), ZN => n2);
   n20 <= '0';
   aMatrix_3_0_port <= '0';
   aMatrix_5_0_port <= '0';
   aMatrix_7_0_port <= '0';
   aMatrix_9_0_port <= '0';
   aMatrix_11_0_port <= '0';
   aMatrix_13_0_port <= '0';
   aMatrix_15_0_port <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity P4_ADDER_N32_NB8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end P4_ADDER_N32_NB8;

architecture SYN_STRUCTURAL of P4_ADDER_N32_NB8 is

   component SUM_GENERATOR_N32_NB8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_N32_NB8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  Co :
            out std_logic_vector (7 downto 0));
   end component;
   
   signal CarriesOut_6_port, CarriesOut_5_port, CarriesOut_4_port, 
      CarriesOut_3_port, CarriesOut_2_port, CarriesOut_1_port, 
      CarriesOut_0_port : std_logic;

begin
   
   CARRY_GENERATOR_INSTANCE : CARRY_GENERATOR_N32_NB8 port map( A(31) => A(31),
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci => Ci, Co(7) =>
                           Co, Co(6) => CarriesOut_6_port, Co(5) => 
                           CarriesOut_5_port, Co(4) => CarriesOut_4_port, Co(3)
                           => CarriesOut_3_port, Co(2) => CarriesOut_2_port, 
                           Co(1) => CarriesOut_1_port, Co(0) => 
                           CarriesOut_0_port);
   SUM_GENERATOR_INSTANCE : SUM_GENERATOR_N32_NB8 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci(7) => 
                           CarriesOut_6_port, Ci(6) => CarriesOut_5_port, Ci(5)
                           => CarriesOut_4_port, Ci(4) => CarriesOut_3_port, 
                           Ci(3) => CarriesOut_2_port, Ci(2) => 
                           CarriesOut_1_port, Ci(1) => CarriesOut_0_port, Ci(0)
                           => Ci, S(31) => S(31), S(30) => S(30), S(29) => 
                           S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFD_31 is

   port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);

end FFD_31;

architecture SYN_BEHAVIORAL of FFD_31 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n4, n1, n_1283 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n4, CK => CLK, Q => Q_port, QN => n_1283);
   U3 : AND2_X1 port map( A1 => n1, A2 => RST, ZN => n4);
   U4 : MUX2_X1 port map( A => Q_port, B => D, S => EN, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LD_224 is

   port( RST, EN, D : in std_logic;  Q : out std_logic);

end LD_224;

architecture SYN_BEHAVIORAL of LD_224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2, N3, n1 : std_logic;

begin
   
   Q_reg : DLH_X1 port map( G => N2, D => N3, Q => Q);
   U3 : AND2_X1 port map( A1 => RST, A2 => D, ZN => N3);
   U4 : NAND2_X1 port map( A1 => n1, A2 => RST, ZN => N2);
   U5 : INV_X1 port map( A => EN, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FU_N5 is

   port( RS1, RS2, RD_MEM, RD_WB : in std_logic_vector (4 downto 0);  RF_WE_MEM
         , RF_WE_WB : in std_logic;  FORWARD_A, FORWARD_B : out 
         std_logic_vector (1 downto 0));

end FU_N5;

architecture SYN_BEHAVIORAL of FU_N5 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27 : std_logic;

begin
   
   U2 : INV_X1 port map( A => n1, ZN => FORWARD_A(0));
   U3 : INV_X1 port map( A => n2, ZN => FORWARD_B(0));
   U4 : NOR4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => 
                           FORWARD_B(1));
   U5 : XOR2_X1 port map( A => RS2(3), B => RD_WB(3), Z => n6);
   U6 : XOR2_X1 port map( A => RS2(1), B => RD_WB(1), Z => n5);
   U7 : XOR2_X1 port map( A => RS2(4), B => RD_WB(4), Z => n4);
   U8 : NAND4_X1 port map( A1 => n7, A2 => n8, A3 => RF_WE_WB, A4 => n2, ZN => 
                           n3);
   U9 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n2)
                           ;
   U10 : NOR3_X1 port map( A1 => n13, A2 => n14, A3 => n15, ZN => n12);
   U11 : XOR2_X1 port map( A => RS2(1), B => RD_MEM(1), Z => n15);
   U12 : XOR2_X1 port map( A => RS2(0), B => RD_MEM(0), Z => n13);
   U13 : XNOR2_X1 port map( A => RD_MEM(3), B => RS2(3), ZN => n11);
   U14 : XNOR2_X1 port map( A => RD_MEM(4), B => RS2(4), ZN => n10);
   U15 : XNOR2_X1 port map( A => RD_MEM(2), B => RS2(2), ZN => n9);
   U16 : XNOR2_X1 port map( A => RD_WB(2), B => RS2(2), ZN => n8);
   U17 : XNOR2_X1 port map( A => RD_WB(0), B => RS2(0), ZN => n7);
   U18 : NOR4_X1 port map( A1 => n16, A2 => n17, A3 => n18, A4 => n19, ZN => 
                           FORWARD_A(1));
   U19 : XOR2_X1 port map( A => RS1(3), B => RD_WB(3), Z => n19);
   U20 : XOR2_X1 port map( A => RS1(1), B => RD_WB(1), Z => n18);
   U21 : XOR2_X1 port map( A => RS1(4), B => RD_WB(4), Z => n17);
   U22 : NAND4_X1 port map( A1 => n20, A2 => n21, A3 => RF_WE_WB, A4 => n1, ZN 
                           => n16);
   U23 : NAND4_X1 port map( A1 => n22, A2 => n23, A3 => n24, A4 => n25, ZN => 
                           n1);
   U24 : NOR3_X1 port map( A1 => n26, A2 => n14, A3 => n27, ZN => n25);
   U25 : XOR2_X1 port map( A => RS1(1), B => RD_MEM(1), Z => n27);
   U26 : INV_X1 port map( A => RF_WE_MEM, ZN => n14);
   U27 : XOR2_X1 port map( A => RS1(0), B => RD_MEM(0), Z => n26);
   U28 : XNOR2_X1 port map( A => RD_MEM(3), B => RS1(3), ZN => n24);
   U29 : XNOR2_X1 port map( A => RD_MEM(4), B => RS1(4), ZN => n23);
   U30 : XNOR2_X1 port map( A => RD_MEM(2), B => RS1(2), ZN => n22);
   U31 : XNOR2_X1 port map( A => RD_WB(2), B => RS1(2), ZN => n21);
   U32 : XNOR2_X1 port map( A => RD_WB(0), B => RS1(0), ZN => n20);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ZERO_DETECTOR_N32_1 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic);

end ZERO_DETECTOR_N32_1;

architecture SYN_STRUCTURAL of ZERO_DETECTOR_N32_1 is

   component AND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, M_4_1_port, M_4_0_port, M_3_3_port, M_3_2_port, 
      M_3_1_port, M_3_0_port, M_2_7_port, M_2_6_port, M_2_5_port, M_2_4_port, 
      M_2_3_port, M_2_2_port, M_2_1_port, M_2_0_port, M_1_15_port, M_1_14_port,
      M_1_13_port, M_1_12_port, M_1_11_port, M_1_10_port, M_1_9_port, 
      M_1_8_port, M_1_7_port, M_1_6_port, M_1_5_port, M_1_4_port, M_1_3_port, 
      M_1_2_port, M_1_1_port, M_1_0_port, M_0_31_port, M_0_30_port, M_0_29_port
      , M_0_28_port, M_0_27_port, M_0_26_port, M_0_25_port, M_0_24_port, 
      M_0_23_port, M_0_22_port, M_0_21_port, M_0_20_port, M_0_19_port, 
      M_0_18_port, M_0_17_port, M_0_16_port, M_0_15_port, M_0_14_port, 
      M_0_13_port, M_0_12_port, M_0_11_port, M_0_10_port, M_0_9_port, 
      M_0_8_port, M_0_7_port, M_0_6_port, M_0_5_port, M_0_4_port, M_0_3_port, 
      M_0_2_port, M_0_1_port, M_0_0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   XOR0_i_0_0 : XNOR2_63 port map( A => A(0), B => X_Logic0_port, Y => 
                           M_0_0_port);
   XOR0_i_0_1 : XNOR2_62 port map( A => A(1), B => X_Logic0_port, Y => 
                           M_0_1_port);
   XOR0_i_0_2 : XNOR2_61 port map( A => A(2), B => X_Logic0_port, Y => 
                           M_0_2_port);
   XOR0_i_0_3 : XNOR2_60 port map( A => A(3), B => X_Logic0_port, Y => 
                           M_0_3_port);
   XOR0_i_0_4 : XNOR2_59 port map( A => A(4), B => X_Logic0_port, Y => 
                           M_0_4_port);
   XOR0_i_0_5 : XNOR2_58 port map( A => A(5), B => X_Logic0_port, Y => 
                           M_0_5_port);
   XOR0_i_0_6 : XNOR2_57 port map( A => A(6), B => X_Logic0_port, Y => 
                           M_0_6_port);
   XOR0_i_0_7 : XNOR2_56 port map( A => A(7), B => X_Logic0_port, Y => 
                           M_0_7_port);
   XOR0_i_0_8 : XNOR2_55 port map( A => A(8), B => X_Logic0_port, Y => 
                           M_0_8_port);
   XOR0_i_0_9 : XNOR2_54 port map( A => A(9), B => X_Logic0_port, Y => 
                           M_0_9_port);
   XOR0_i_0_10 : XNOR2_53 port map( A => A(10), B => X_Logic0_port, Y => 
                           M_0_10_port);
   XOR0_i_0_11 : XNOR2_52 port map( A => A(11), B => X_Logic0_port, Y => 
                           M_0_11_port);
   XOR0_i_0_12 : XNOR2_51 port map( A => A(12), B => X_Logic0_port, Y => 
                           M_0_12_port);
   XOR0_i_0_13 : XNOR2_50 port map( A => A(13), B => X_Logic0_port, Y => 
                           M_0_13_port);
   XOR0_i_0_14 : XNOR2_49 port map( A => A(14), B => X_Logic0_port, Y => 
                           M_0_14_port);
   XOR0_i_0_15 : XNOR2_48 port map( A => A(15), B => X_Logic0_port, Y => 
                           M_0_15_port);
   XOR0_i_0_16 : XNOR2_47 port map( A => A(16), B => X_Logic0_port, Y => 
                           M_0_16_port);
   XOR0_i_0_17 : XNOR2_46 port map( A => A(17), B => X_Logic0_port, Y => 
                           M_0_17_port);
   XOR0_i_0_18 : XNOR2_45 port map( A => A(18), B => X_Logic0_port, Y => 
                           M_0_18_port);
   XOR0_i_0_19 : XNOR2_44 port map( A => A(19), B => X_Logic0_port, Y => 
                           M_0_19_port);
   XOR0_i_0_20 : XNOR2_43 port map( A => A(20), B => X_Logic0_port, Y => 
                           M_0_20_port);
   XOR0_i_0_21 : XNOR2_42 port map( A => A(21), B => X_Logic0_port, Y => 
                           M_0_21_port);
   XOR0_i_0_22 : XNOR2_41 port map( A => A(22), B => X_Logic0_port, Y => 
                           M_0_22_port);
   XOR0_i_0_23 : XNOR2_40 port map( A => A(23), B => X_Logic0_port, Y => 
                           M_0_23_port);
   XOR0_i_0_24 : XNOR2_39 port map( A => A(24), B => X_Logic0_port, Y => 
                           M_0_24_port);
   XOR0_i_0_25 : XNOR2_38 port map( A => A(25), B => X_Logic0_port, Y => 
                           M_0_25_port);
   XOR0_i_0_26 : XNOR2_37 port map( A => A(26), B => X_Logic0_port, Y => 
                           M_0_26_port);
   XOR0_i_0_27 : XNOR2_36 port map( A => A(27), B => X_Logic0_port, Y => 
                           M_0_27_port);
   XOR0_i_0_28 : XNOR2_35 port map( A => A(28), B => X_Logic0_port, Y => 
                           M_0_28_port);
   XOR0_i_0_29 : XNOR2_34 port map( A => A(29), B => X_Logic0_port, Y => 
                           M_0_29_port);
   XOR0_i_0_30 : XNOR2_33 port map( A => A(30), B => X_Logic0_port, Y => 
                           M_0_30_port);
   XOR0_i_0_31 : XNOR2_32 port map( A => A(31), B => X_Logic0_port, Y => 
                           M_0_31_port);
   AND_i_1_0 : AND2_61 port map( A => M_0_0_port, B => M_0_1_port, Y => 
                           M_1_0_port);
   AND_i_1_1 : AND2_60 port map( A => M_0_2_port, B => M_0_3_port, Y => 
                           M_1_1_port);
   AND_i_1_2 : AND2_59 port map( A => M_0_4_port, B => M_0_5_port, Y => 
                           M_1_2_port);
   AND_i_1_3 : AND2_58 port map( A => M_0_6_port, B => M_0_7_port, Y => 
                           M_1_3_port);
   AND_i_1_4 : AND2_57 port map( A => M_0_8_port, B => M_0_9_port, Y => 
                           M_1_4_port);
   AND_i_1_5 : AND2_56 port map( A => M_0_10_port, B => M_0_11_port, Y => 
                           M_1_5_port);
   AND_i_1_6 : AND2_55 port map( A => M_0_12_port, B => M_0_13_port, Y => 
                           M_1_6_port);
   AND_i_1_7 : AND2_54 port map( A => M_0_14_port, B => M_0_15_port, Y => 
                           M_1_7_port);
   AND_i_1_8 : AND2_53 port map( A => M_0_16_port, B => M_0_17_port, Y => 
                           M_1_8_port);
   AND_i_1_9 : AND2_52 port map( A => M_0_18_port, B => M_0_19_port, Y => 
                           M_1_9_port);
   AND_i_1_10 : AND2_51 port map( A => M_0_20_port, B => M_0_21_port, Y => 
                           M_1_10_port);
   AND_i_1_11 : AND2_50 port map( A => M_0_22_port, B => M_0_23_port, Y => 
                           M_1_11_port);
   AND_i_1_12 : AND2_49 port map( A => M_0_24_port, B => M_0_25_port, Y => 
                           M_1_12_port);
   AND_i_1_13 : AND2_48 port map( A => M_0_26_port, B => M_0_27_port, Y => 
                           M_1_13_port);
   AND_i_1_14 : AND2_47 port map( A => M_0_28_port, B => M_0_29_port, Y => 
                           M_1_14_port);
   AND_i_1_15 : AND2_46 port map( A => M_0_30_port, B => M_0_31_port, Y => 
                           M_1_15_port);
   AND_i_2_0 : AND2_45 port map( A => M_1_0_port, B => M_1_1_port, Y => 
                           M_2_0_port);
   AND_i_2_1 : AND2_44 port map( A => M_1_2_port, B => M_1_3_port, Y => 
                           M_2_1_port);
   AND_i_2_2 : AND2_43 port map( A => M_1_4_port, B => M_1_5_port, Y => 
                           M_2_2_port);
   AND_i_2_3 : AND2_42 port map( A => M_1_6_port, B => M_1_7_port, Y => 
                           M_2_3_port);
   AND_i_2_4 : AND2_41 port map( A => M_1_8_port, B => M_1_9_port, Y => 
                           M_2_4_port);
   AND_i_2_5 : AND2_40 port map( A => M_1_10_port, B => M_1_11_port, Y => 
                           M_2_5_port);
   AND_i_2_6 : AND2_39 port map( A => M_1_12_port, B => M_1_13_port, Y => 
                           M_2_6_port);
   AND_i_2_7 : AND2_38 port map( A => M_1_14_port, B => M_1_15_port, Y => 
                           M_2_7_port);
   AND_i_3_0 : AND2_37 port map( A => M_2_0_port, B => M_2_1_port, Y => 
                           M_3_0_port);
   AND_i_3_1 : AND2_36 port map( A => M_2_2_port, B => M_2_3_port, Y => 
                           M_3_1_port);
   AND_i_3_2 : AND2_35 port map( A => M_2_4_port, B => M_2_5_port, Y => 
                           M_3_2_port);
   AND_i_3_3 : AND2_34 port map( A => M_2_6_port, B => M_2_7_port, Y => 
                           M_3_3_port);
   AND_i_4_0 : AND2_33 port map( A => M_3_0_port, B => M_3_1_port, Y => 
                           M_4_0_port);
   AND_i_4_1 : AND2_32 port map( A => M_3_2_port, B => M_3_3_port, Y => 
                           M_4_1_port);
   AND_i_5_0 : AND2_31 port map( A => M_4_0_port, B => M_4_1_port, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_L_320 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_L_320;

architecture SYN_BEHAVIORAL of MUX21_L_320 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A, B => B, S => S, Z => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_NB8 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
         std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);  Z
         : out std_logic);

end ALU_N32_NB8;

architecture SYN_BEHAVIORAL of ALU_N32_NB8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X2
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component ZERO_DETECTOR_N32_0
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic);
   end component;
   
   component COMPARATOR_N32
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic_vector 
            (3 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component LOGIC_N32
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic_vector 
            (1 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component BARREL_SHIFTER_RIGHT_N32
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component BARREL_SHIFTER_LEFT_N32
      port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector
            (31 downto 0));
   end component;
   
   component BOOTH_MULTIPLIER_N32
      port( A, B : in std_logic_vector (15 downto 0);  P : out std_logic_vector
            (31 downto 0));
   end component;
   
   component P4_ADDER_N32_NB8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal Y_31_port, Y_30_port, Y_29_port, Y_28_port, Y_27_port, Y_26_port, 
      Y_25_port, Y_24_port, Y_23_port, Y_22_port, Y_21_port, Y_20_port, 
      Y_19_port, Y_18_port, Y_17_port, Y_16_port, Y_15_port, Y_14_port, 
      Y_13_port, Y_12_port, Y_11_port, Y_10_port, Y_9_port, Y_8_port, Y_7_port,
      Y_6_port, Y_5_port, Y_4_port, Y_3_port, Y_2_port, Y_1_port, Y_0_port, N96
      , OP_A_31_port, OP_A_30_port, OP_A_29_port, OP_A_28_port, OP_A_27_port, 
      OP_A_26_port, OP_A_25_port, OP_A_24_port, OP_A_23_port, OP_A_22_port, 
      OP_A_21_port, OP_A_20_port, OP_A_19_port, OP_A_18_port, OP_A_17_port, 
      OP_A_16_port, OP_A_15_port, OP_A_14_port, OP_A_13_port, OP_A_12_port, 
      OP_A_11_port, OP_A_10_port, OP_A_9_port, OP_A_8_port, OP_A_7_port, 
      OP_A_6_port, OP_A_5_port, OP_A_4_port, OP_A_3_port, OP_A_2_port, 
      OP_A_1_port, OP_A_0_port, OP_B_31_port, OP_B_30_port, OP_B_29_port, 
      OP_B_28_port, OP_B_27_port, OP_B_26_port, OP_B_25_port, OP_B_24_port, 
      OP_B_23_port, OP_B_22_port, OP_B_21_port, OP_B_20_port, OP_B_19_port, 
      OP_B_18_port, OP_B_17_port, OP_B_16_port, OP_B_15_port, OP_B_14_port, 
      OP_B_13_port, OP_B_12_port, OP_B_11_port, OP_B_10_port, OP_B_9_port, 
      OP_B_8_port, OP_B_7_port, OP_B_6_port, OP_B_5_port, OP_B_4_port, 
      OP_B_3_port, OP_B_2_port, OP_B_1_port, OP_B_0_port, Y_SHIFTL_31_port, 
      Y_SHIFTL_30_port, Y_SHIFTL_29_port, Y_SHIFTL_28_port, Y_SHIFTL_27_port, 
      Y_SHIFTL_26_port, Y_SHIFTL_25_port, Y_SHIFTL_24_port, Y_SHIFTL_23_port, 
      Y_SHIFTL_22_port, Y_SHIFTL_21_port, Y_SHIFTL_20_port, Y_SHIFTL_19_port, 
      Y_SHIFTL_18_port, Y_SHIFTL_17_port, Y_SHIFTL_16_port, Y_SHIFTL_15_port, 
      Y_SHIFTL_14_port, Y_SHIFTL_13_port, Y_SHIFTL_12_port, Y_SHIFTL_11_port, 
      Y_SHIFTL_10_port, Y_SHIFTL_9_port, Y_SHIFTL_8_port, Y_SHIFTL_7_port, 
      Y_SHIFTL_6_port, Y_SHIFTL_5_port, Y_SHIFTL_4_port, Y_SHIFTL_3_port, 
      Y_SHIFTL_2_port, Y_SHIFTL_1_port, Y_SHIFTL_0_port, Y_MUL_31_port, 
      Y_MUL_30_port, Y_MUL_29_port, Y_MUL_28_port, Y_MUL_27_port, Y_MUL_26_port
      , Y_MUL_25_port, Y_MUL_24_port, Y_MUL_23_port, Y_MUL_22_port, 
      Y_MUL_21_port, Y_MUL_20_port, Y_MUL_19_port, Y_MUL_18_port, Y_MUL_17_port
      , Y_MUL_16_port, Y_MUL_15_port, Y_MUL_14_port, Y_MUL_13_port, 
      Y_MUL_12_port, Y_MUL_11_port, Y_MUL_10_port, Y_MUL_9_port, Y_MUL_8_port, 
      Y_MUL_7_port, Y_MUL_6_port, Y_MUL_5_port, Y_MUL_4_port, Y_MUL_3_port, 
      Y_MUL_2_port, Y_MUL_1_port, Y_MUL_0_port, OP_Ci, Y_SUM_31_port, 
      Y_SUM_30_port, Y_SUM_29_port, Y_SUM_28_port, Y_SUM_27_port, Y_SUM_26_port
      , Y_SUM_25_port, Y_SUM_24_port, Y_SUM_23_port, Y_SUM_22_port, 
      Y_SUM_21_port, Y_SUM_20_port, Y_SUM_19_port, Y_SUM_18_port, Y_SUM_17_port
      , Y_SUM_16_port, Y_SUM_15_port, Y_SUM_14_port, Y_SUM_13_port, 
      Y_SUM_12_port, Y_SUM_11_port, Y_SUM_10_port, Y_SUM_9_port, Y_SUM_8_port, 
      Y_SUM_7_port, Y_SUM_6_port, Y_SUM_5_port, Y_SUM_4_port, Y_SUM_3_port, 
      Y_SUM_2_port, Y_SUM_1_port, Y_SUM_0_port, OP_LOGIC_1_port, 
      OP_LOGIC_0_port, Y_LOGIC_31_port, Y_LOGIC_30_port, Y_LOGIC_29_port, 
      Y_LOGIC_28_port, Y_LOGIC_27_port, Y_LOGIC_26_port, Y_LOGIC_25_port, 
      Y_LOGIC_24_port, Y_LOGIC_23_port, Y_LOGIC_22_port, Y_LOGIC_21_port, 
      Y_LOGIC_20_port, Y_LOGIC_19_port, Y_LOGIC_18_port, Y_LOGIC_17_port, 
      Y_LOGIC_16_port, Y_LOGIC_15_port, Y_LOGIC_14_port, Y_LOGIC_13_port, 
      Y_LOGIC_12_port, Y_LOGIC_11_port, Y_LOGIC_10_port, Y_LOGIC_9_port, 
      Y_LOGIC_8_port, Y_LOGIC_7_port, Y_LOGIC_6_port, Y_LOGIC_5_port, 
      Y_LOGIC_4_port, Y_LOGIC_3_port, Y_LOGIC_2_port, Y_LOGIC_1_port, 
      Y_LOGIC_0_port, OP_SHIFT, Y_SHIFTR_31_port, Y_SHIFTR_30_port, 
      Y_SHIFTR_29_port, Y_SHIFTR_28_port, Y_SHIFTR_27_port, Y_SHIFTR_26_port, 
      Y_SHIFTR_25_port, Y_SHIFTR_24_port, Y_SHIFTR_23_port, Y_SHIFTR_22_port, 
      Y_SHIFTR_21_port, Y_SHIFTR_20_port, Y_SHIFTR_19_port, Y_SHIFTR_18_port, 
      Y_SHIFTR_17_port, Y_SHIFTR_16_port, Y_SHIFTR_15_port, Y_SHIFTR_14_port, 
      Y_SHIFTR_13_port, Y_SHIFTR_12_port, Y_SHIFTR_11_port, Y_SHIFTR_10_port, 
      Y_SHIFTR_9_port, Y_SHIFTR_8_port, Y_SHIFTR_7_port, Y_SHIFTR_6_port, 
      Y_SHIFTR_5_port, Y_SHIFTR_4_port, Y_SHIFTR_3_port, Y_SHIFTR_2_port, 
      Y_SHIFTR_1_port, Y_SHIFTR_0_port, OP_COMPARE_3_port, OP_COMPARE_2_port, 
      OP_COMPARE_1_port, OP_COMPARE_0_port, Y_COMPARE_0_port, N246, N247, N248,
      N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, 
      N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, 
      N273, N274, N275, N276, N277, N278, N279, N280, N281, N285, N286, N287, 
      N288, N289, n225, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96_port, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, 
      n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, 
      n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, 
      n_1311, n_1312, n_1313, n_1314, n_1315 : std_logic;

begin
   Y <= ( Y_31_port, Y_30_port, Y_29_port, Y_28_port, Y_27_port, Y_26_port, 
      Y_25_port, Y_24_port, Y_23_port, Y_22_port, Y_21_port, Y_20_port, 
      Y_19_port, Y_18_port, Y_17_port, Y_16_port, Y_15_port, Y_14_port, 
      Y_13_port, Y_12_port, Y_11_port, Y_10_port, Y_9_port, Y_8_port, Y_7_port,
      Y_6_port, Y_5_port, Y_4_port, Y_3_port, Y_2_port, Y_1_port, Y_0_port );
   
   OP_COMPARE_reg_3_inst : DLH_X1 port map( G => N285, D => N289, Q => 
                           OP_COMPARE_3_port);
   OP_COMPARE_reg_2_inst : DLH_X1 port map( G => N285, D => N288, Q => 
                           OP_COMPARE_2_port);
   OP_COMPARE_reg_1_inst : DLH_X1 port map( G => N285, D => N287, Q => 
                           OP_COMPARE_1_port);
   OP_COMPARE_reg_0_inst : DLH_X1 port map( G => N285, D => N286, Q => 
                           OP_COMPARE_0_port);
   OP_A_reg_31_inst : DLH_X1 port map( G => N246, D => OP1(31), Q => 
                           OP_A_31_port);
   OP_A_reg_30_inst : DLH_X1 port map( G => N246, D => OP1(30), Q => 
                           OP_A_30_port);
   OP_A_reg_29_inst : DLH_X1 port map( G => N246, D => OP1(29), Q => 
                           OP_A_29_port);
   OP_A_reg_28_inst : DLH_X1 port map( G => N246, D => OP1(28), Q => 
                           OP_A_28_port);
   OP_A_reg_27_inst : DLH_X1 port map( G => N246, D => OP1(27), Q => 
                           OP_A_27_port);
   OP_A_reg_26_inst : DLH_X1 port map( G => N246, D => OP1(26), Q => 
                           OP_A_26_port);
   OP_A_reg_25_inst : DLH_X1 port map( G => N246, D => OP1(25), Q => 
                           OP_A_25_port);
   OP_A_reg_24_inst : DLH_X1 port map( G => N246, D => OP1(24), Q => 
                           OP_A_24_port);
   OP_A_reg_23_inst : DLH_X1 port map( G => N246, D => OP1(23), Q => 
                           OP_A_23_port);
   OP_A_reg_22_inst : DLH_X1 port map( G => N246, D => OP1(22), Q => 
                           OP_A_22_port);
   OP_A_reg_21_inst : DLH_X1 port map( G => N246, D => OP1(21), Q => 
                           OP_A_21_port);
   OP_A_reg_20_inst : DLH_X1 port map( G => N246, D => OP1(20), Q => 
                           OP_A_20_port);
   OP_A_reg_19_inst : DLH_X1 port map( G => N246, D => OP1(19), Q => 
                           OP_A_19_port);
   OP_A_reg_18_inst : DLH_X1 port map( G => N246, D => OP1(18), Q => 
                           OP_A_18_port);
   OP_A_reg_17_inst : DLH_X1 port map( G => N246, D => OP1(17), Q => 
                           OP_A_17_port);
   OP_A_reg_16_inst : DLH_X1 port map( G => N246, D => OP1(16), Q => 
                           OP_A_16_port);
   OP_A_reg_15_inst : DLH_X1 port map( G => N246, D => OP1(15), Q => 
                           OP_A_15_port);
   OP_A_reg_13_inst : DLH_X1 port map( G => N246, D => OP1(13), Q => 
                           OP_A_13_port);
   OP_A_reg_9_inst : DLH_X1 port map( G => N246, D => OP1(9), Q => OP_A_9_port)
                           ;
   OP_A_reg_5_inst : DLH_X1 port map( G => N246, D => OP1(5), Q => OP_A_5_port)
                           ;
   OP_B_reg_31_inst : DLH_X1 port map( G => N246, D => N278, Q => OP_B_31_port)
                           ;
   OP_B_reg_30_inst : DLH_X1 port map( G => N246, D => N277, Q => OP_B_30_port)
                           ;
   OP_B_reg_29_inst : DLH_X1 port map( G => N246, D => N276, Q => OP_B_29_port)
                           ;
   OP_B_reg_28_inst : DLH_X1 port map( G => N246, D => N275, Q => OP_B_28_port)
                           ;
   OP_B_reg_27_inst : DLH_X1 port map( G => N246, D => N274, Q => OP_B_27_port)
                           ;
   OP_B_reg_26_inst : DLH_X1 port map( G => N246, D => N273, Q => OP_B_26_port)
                           ;
   OP_B_reg_25_inst : DLH_X1 port map( G => N246, D => N272, Q => OP_B_25_port)
                           ;
   OP_B_reg_24_inst : DLH_X1 port map( G => N246, D => N271, Q => OP_B_24_port)
                           ;
   OP_B_reg_23_inst : DLH_X1 port map( G => N246, D => N270, Q => OP_B_23_port)
                           ;
   OP_B_reg_22_inst : DLH_X1 port map( G => N246, D => N269, Q => OP_B_22_port)
                           ;
   OP_B_reg_21_inst : DLH_X1 port map( G => N246, D => N268, Q => OP_B_21_port)
                           ;
   OP_B_reg_20_inst : DLH_X1 port map( G => N246, D => N267, Q => OP_B_20_port)
                           ;
   OP_B_reg_19_inst : DLH_X1 port map( G => N246, D => N266, Q => OP_B_19_port)
                           ;
   OP_B_reg_18_inst : DLH_X1 port map( G => N246, D => N265, Q => OP_B_18_port)
                           ;
   OP_B_reg_17_inst : DLH_X1 port map( G => N246, D => N264, Q => OP_B_17_port)
                           ;
   OP_B_reg_16_inst : DLH_X1 port map( G => N246, D => N263, Q => OP_B_16_port)
                           ;
   OP_B_reg_15_inst : DLH_X1 port map( G => N246, D => N262, Q => OP_B_15_port)
                           ;
   OP_B_reg_14_inst : DLH_X1 port map( G => N246, D => N261, Q => OP_B_14_port)
                           ;
   OP_B_reg_13_inst : DLH_X1 port map( G => N246, D => N260, Q => OP_B_13_port)
                           ;
   OP_B_reg_12_inst : DLH_X1 port map( G => N246, D => N259, Q => OP_B_12_port)
                           ;
   OP_B_reg_11_inst : DLH_X1 port map( G => N246, D => N258, Q => OP_B_11_port)
                           ;
   OP_B_reg_10_inst : DLH_X1 port map( G => N246, D => N257, Q => OP_B_10_port)
                           ;
   OP_B_reg_9_inst : DLH_X1 port map( G => N246, D => N256, Q => OP_B_9_port);
   OP_B_reg_8_inst : DLH_X1 port map( G => N246, D => N255, Q => OP_B_8_port);
   OP_B_reg_7_inst : DLH_X1 port map( G => N246, D => N254, Q => OP_B_7_port);
   OP_B_reg_6_inst : DLH_X1 port map( G => N246, D => N253, Q => OP_B_6_port);
   OP_B_reg_5_inst : DLH_X1 port map( G => N246, D => N252, Q => OP_B_5_port);
   OP_B_reg_4_inst : DLH_X1 port map( G => N246, D => N251, Q => OP_B_4_port);
   OP_B_reg_3_inst : DLH_X1 port map( G => N246, D => N250, Q => OP_B_3_port);
   OP_B_reg_2_inst : DLH_X1 port map( G => N246, D => N249, Q => OP_B_2_port);
   OP_B_reg_1_inst : DLH_X1 port map( G => N246, D => N248, Q => OP_B_1_port);
   OP_B_reg_0_inst : DLH_X1 port map( G => N246, D => N247, Q => OP_B_0_port);
   OP_Ci_reg : DLH_X1 port map( G => N279, D => N280, Q => OP_Ci);
   OP_LOGIC_reg_1_inst : DLH_X1 port map( G => N281, D => n182, Q => 
                           OP_LOGIC_1_port);
   OP_LOGIC_reg_0_inst : DLH_X1 port map( G => N281, D => n183, Q => 
                           OP_LOGIC_0_port);
   OP_SHIFT_reg : DLL_X1 port map( D => N96, GN => n225, Q => OP_SHIFT);
   SUM : P4_ADDER_N32_NB8 port map( A(31) => OP_A_31_port, A(30) => 
                           OP_A_30_port, A(29) => OP_A_29_port, A(28) => 
                           OP_A_28_port, A(27) => OP_A_27_port, A(26) => 
                           OP_A_26_port, A(25) => OP_A_25_port, A(24) => 
                           OP_A_24_port, A(23) => OP_A_23_port, A(22) => 
                           OP_A_22_port, A(21) => OP_A_21_port, A(20) => 
                           OP_A_20_port, A(19) => OP_A_19_port, A(18) => 
                           OP_A_18_port, A(17) => OP_A_17_port, A(16) => 
                           OP_A_16_port, A(15) => n18, A(14) => OP_A_14_port, 
                           A(13) => OP_A_13_port, A(12) => OP_A_12_port, A(11) 
                           => OP_A_11_port, A(10) => OP_A_10_port, A(9) => 
                           OP_A_9_port, A(8) => OP_A_8_port, A(7) => 
                           OP_A_7_port, A(6) => OP_A_6_port, A(5) => 
                           OP_A_5_port, A(4) => OP_A_4_port, A(3) => 
                           OP_A_3_port, A(2) => OP_A_2_port, A(1) => 
                           OP_A_1_port, A(0) => OP_A_0_port, B(31) => 
                           OP_B_31_port, B(30) => OP_B_30_port, B(29) => 
                           OP_B_29_port, B(28) => OP_B_28_port, B(27) => 
                           OP_B_27_port, B(26) => OP_B_26_port, B(25) => 
                           OP_B_25_port, B(24) => OP_B_24_port, B(23) => 
                           OP_B_23_port, B(22) => OP_B_22_port, B(21) => 
                           OP_B_21_port, B(20) => OP_B_20_port, B(19) => 
                           OP_B_19_port, B(18) => OP_B_18_port, B(17) => 
                           OP_B_17_port, B(16) => OP_B_16_port, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n12, B(3) => n14, B(2) => n8, 
                           B(1) => n16, B(0) => n10, Ci => OP_Ci, S(31) => 
                           Y_SUM_31_port, S(30) => Y_SUM_30_port, S(29) => 
                           Y_SUM_29_port, S(28) => Y_SUM_28_port, S(27) => 
                           Y_SUM_27_port, S(26) => Y_SUM_26_port, S(25) => 
                           Y_SUM_25_port, S(24) => Y_SUM_24_port, S(23) => 
                           Y_SUM_23_port, S(22) => Y_SUM_22_port, S(21) => 
                           Y_SUM_21_port, S(20) => Y_SUM_20_port, S(19) => 
                           Y_SUM_19_port, S(18) => Y_SUM_18_port, S(17) => 
                           Y_SUM_17_port, S(16) => Y_SUM_16_port, S(15) => 
                           Y_SUM_15_port, S(14) => Y_SUM_14_port, S(13) => 
                           Y_SUM_13_port, S(12) => Y_SUM_12_port, S(11) => 
                           Y_SUM_11_port, S(10) => Y_SUM_10_port, S(9) => 
                           Y_SUM_9_port, S(8) => Y_SUM_8_port, S(7) => 
                           Y_SUM_7_port, S(6) => Y_SUM_6_port, S(5) => 
                           Y_SUM_5_port, S(4) => Y_SUM_4_port, S(3) => 
                           Y_SUM_3_port, S(2) => Y_SUM_2_port, S(1) => 
                           Y_SUM_1_port, S(0) => Y_SUM_0_port, Co => n_1284);
   MUL : BOOTH_MULTIPLIER_N32 port map( A(15) => n18, A(14) => OP_A_14_port, 
                           A(13) => OP_A_13_port, A(12) => OP_A_12_port, A(11) 
                           => OP_A_11_port, A(10) => OP_A_10_port, A(9) => 
                           OP_A_9_port, A(8) => OP_A_8_port, A(7) => 
                           OP_A_7_port, A(6) => OP_A_6_port, A(5) => 
                           OP_A_5_port, A(4) => OP_A_4_port, A(3) => 
                           OP_A_3_port, A(2) => OP_A_2_port, A(1) => 
                           OP_A_1_port, A(0) => OP_A_0_port, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n12, B(3) => n14, B(2) => n8, 
                           B(1) => n16, B(0) => n10, P(31) => Y_MUL_31_port, 
                           P(30) => Y_MUL_30_port, P(29) => Y_MUL_29_port, 
                           P(28) => Y_MUL_28_port, P(27) => Y_MUL_27_port, 
                           P(26) => Y_MUL_26_port, P(25) => Y_MUL_25_port, 
                           P(24) => Y_MUL_24_port, P(23) => Y_MUL_23_port, 
                           P(22) => Y_MUL_22_port, P(21) => Y_MUL_21_port, 
                           P(20) => Y_MUL_20_port, P(19) => Y_MUL_19_port, 
                           P(18) => Y_MUL_18_port, P(17) => Y_MUL_17_port, 
                           P(16) => Y_MUL_16_port, P(15) => Y_MUL_15_port, 
                           P(14) => Y_MUL_14_port, P(13) => Y_MUL_13_port, 
                           P(12) => Y_MUL_12_port, P(11) => Y_MUL_11_port, 
                           P(10) => Y_MUL_10_port, P(9) => Y_MUL_9_port, P(8) 
                           => Y_MUL_8_port, P(7) => Y_MUL_7_port, P(6) => 
                           Y_MUL_6_port, P(5) => Y_MUL_5_port, P(4) => 
                           Y_MUL_4_port, P(3) => Y_MUL_3_port, P(2) => 
                           Y_MUL_2_port, P(1) => Y_MUL_1_port, P(0) => 
                           Y_MUL_0_port);
   BSL : BARREL_SHIFTER_LEFT_N32 port map( A(31) => OP_A_31_port, A(30) => 
                           OP_A_30_port, A(29) => OP_A_29_port, A(28) => 
                           OP_A_28_port, A(27) => OP_A_27_port, A(26) => 
                           OP_A_26_port, A(25) => OP_A_25_port, A(24) => 
                           OP_A_24_port, A(23) => OP_A_23_port, A(22) => 
                           OP_A_22_port, A(21) => OP_A_21_port, A(20) => 
                           OP_A_20_port, A(19) => OP_A_19_port, A(18) => 
                           OP_A_18_port, A(17) => OP_A_17_port, A(16) => 
                           OP_A_16_port, A(15) => n18, A(14) => OP_A_14_port, 
                           A(13) => OP_A_13_port, A(12) => OP_A_12_port, A(11) 
                           => OP_A_11_port, A(10) => OP_A_10_port, A(9) => 
                           OP_A_9_port, A(8) => OP_A_8_port, A(7) => 
                           OP_A_7_port, A(6) => OP_A_6_port, A(5) => 
                           OP_A_5_port, A(4) => OP_A_4_port, A(3) => 
                           OP_A_3_port, A(2) => OP_A_2_port, A(1) => 
                           OP_A_1_port, A(0) => OP_A_0_port, B(31) => 
                           OP_B_31_port, B(30) => OP_B_30_port, B(29) => 
                           OP_B_29_port, B(28) => OP_B_28_port, B(27) => 
                           OP_B_27_port, B(26) => OP_B_26_port, B(25) => 
                           OP_B_25_port, B(24) => OP_B_24_port, B(23) => 
                           OP_B_23_port, B(22) => OP_B_22_port, B(21) => 
                           OP_B_21_port, B(20) => OP_B_20_port, B(19) => 
                           OP_B_19_port, B(18) => OP_B_18_port, B(17) => 
                           OP_B_17_port, B(16) => OP_B_16_port, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n12, B(3) => n14, B(2) => n8, 
                           B(1) => n16, B(0) => n10, Y(31) => Y_SHIFTL_31_port,
                           Y(30) => Y_SHIFTL_30_port, Y(29) => Y_SHIFTL_29_port
                           , Y(28) => Y_SHIFTL_28_port, Y(27) => 
                           Y_SHIFTL_27_port, Y(26) => Y_SHIFTL_26_port, Y(25) 
                           => Y_SHIFTL_25_port, Y(24) => Y_SHIFTL_24_port, 
                           Y(23) => Y_SHIFTL_23_port, Y(22) => Y_SHIFTL_22_port
                           , Y(21) => Y_SHIFTL_21_port, Y(20) => 
                           Y_SHIFTL_20_port, Y(19) => Y_SHIFTL_19_port, Y(18) 
                           => Y_SHIFTL_18_port, Y(17) => Y_SHIFTL_17_port, 
                           Y(16) => Y_SHIFTL_16_port, Y(15) => Y_SHIFTL_15_port
                           , Y(14) => Y_SHIFTL_14_port, Y(13) => 
                           Y_SHIFTL_13_port, Y(12) => Y_SHIFTL_12_port, Y(11) 
                           => Y_SHIFTL_11_port, Y(10) => Y_SHIFTL_10_port, Y(9)
                           => Y_SHIFTL_9_port, Y(8) => Y_SHIFTL_8_port, Y(7) =>
                           Y_SHIFTL_7_port, Y(6) => Y_SHIFTL_6_port, Y(5) => 
                           Y_SHIFTL_5_port, Y(4) => Y_SHIFTL_4_port, Y(3) => 
                           Y_SHIFTL_3_port, Y(2) => Y_SHIFTL_2_port, Y(1) => 
                           Y_SHIFTL_1_port, Y(0) => Y_SHIFTL_0_port);
   BSR : BARREL_SHIFTER_RIGHT_N32 port map( A(31) => OP_A_31_port, A(30) => 
                           OP_A_30_port, A(29) => OP_A_29_port, A(28) => 
                           OP_A_28_port, A(27) => OP_A_27_port, A(26) => 
                           OP_A_26_port, A(25) => OP_A_25_port, A(24) => 
                           OP_A_24_port, A(23) => OP_A_23_port, A(22) => 
                           OP_A_22_port, A(21) => OP_A_21_port, A(20) => 
                           OP_A_20_port, A(19) => OP_A_19_port, A(18) => 
                           OP_A_18_port, A(17) => OP_A_17_port, A(16) => 
                           OP_A_16_port, A(15) => n18, A(14) => OP_A_14_port, 
                           A(13) => OP_A_13_port, A(12) => OP_A_12_port, A(11) 
                           => OP_A_11_port, A(10) => OP_A_10_port, A(9) => 
                           OP_A_9_port, A(8) => OP_A_8_port, A(7) => 
                           OP_A_7_port, A(6) => OP_A_6_port, A(5) => 
                           OP_A_5_port, A(4) => OP_A_4_port, A(3) => 
                           OP_A_3_port, A(2) => OP_A_2_port, A(1) => 
                           OP_A_1_port, A(0) => OP_A_0_port, B(31) => 
                           OP_B_31_port, B(30) => OP_B_30_port, B(29) => 
                           OP_B_29_port, B(28) => OP_B_28_port, B(27) => 
                           OP_B_27_port, B(26) => OP_B_26_port, B(25) => 
                           OP_B_25_port, B(24) => OP_B_24_port, B(23) => 
                           OP_B_23_port, B(22) => OP_B_22_port, B(21) => 
                           OP_B_21_port, B(20) => OP_B_20_port, B(19) => 
                           OP_B_19_port, B(18) => OP_B_18_port, B(17) => 
                           OP_B_17_port, B(16) => OP_B_16_port, B(15) => 
                           OP_B_15_port, B(14) => OP_B_14_port, B(13) => 
                           OP_B_13_port, B(12) => OP_B_12_port, B(11) => 
                           OP_B_11_port, B(10) => OP_B_10_port, B(9) => 
                           OP_B_9_port, B(8) => OP_B_8_port, B(7) => 
                           OP_B_7_port, B(6) => OP_B_6_port, B(5) => 
                           OP_B_5_port, B(4) => n12, B(3) => n14, B(2) => n8, 
                           B(1) => n16, B(0) => n10, S => OP_SHIFT, Y(31) => 
                           Y_SHIFTR_31_port, Y(30) => Y_SHIFTR_30_port, Y(29) 
                           => Y_SHIFTR_29_port, Y(28) => Y_SHIFTR_28_port, 
                           Y(27) => Y_SHIFTR_27_port, Y(26) => Y_SHIFTR_26_port
                           , Y(25) => Y_SHIFTR_25_port, Y(24) => 
                           Y_SHIFTR_24_port, Y(23) => Y_SHIFTR_23_port, Y(22) 
                           => Y_SHIFTR_22_port, Y(21) => Y_SHIFTR_21_port, 
                           Y(20) => Y_SHIFTR_20_port, Y(19) => Y_SHIFTR_19_port
                           , Y(18) => Y_SHIFTR_18_port, Y(17) => 
                           Y_SHIFTR_17_port, Y(16) => Y_SHIFTR_16_port, Y(15) 
                           => Y_SHIFTR_15_port, Y(14) => Y_SHIFTR_14_port, 
                           Y(13) => Y_SHIFTR_13_port, Y(12) => Y_SHIFTR_12_port
                           , Y(11) => Y_SHIFTR_11_port, Y(10) => 
                           Y_SHIFTR_10_port, Y(9) => Y_SHIFTR_9_port, Y(8) => 
                           Y_SHIFTR_8_port, Y(7) => Y_SHIFTR_7_port, Y(6) => 
                           Y_SHIFTR_6_port, Y(5) => Y_SHIFTR_5_port, Y(4) => 
                           Y_SHIFTR_4_port, Y(3) => Y_SHIFTR_3_port, Y(2) => 
                           Y_SHIFTR_2_port, Y(1) => Y_SHIFTR_1_port, Y(0) => 
                           Y_SHIFTR_0_port);
   LOG : LOGIC_N32 port map( A(31) => OP_A_31_port, A(30) => OP_A_30_port, 
                           A(29) => OP_A_29_port, A(28) => OP_A_28_port, A(27) 
                           => OP_A_27_port, A(26) => OP_A_26_port, A(25) => 
                           OP_A_25_port, A(24) => OP_A_24_port, A(23) => 
                           OP_A_23_port, A(22) => OP_A_22_port, A(21) => 
                           OP_A_21_port, A(20) => OP_A_20_port, A(19) => 
                           OP_A_19_port, A(18) => OP_A_18_port, A(17) => 
                           OP_A_17_port, A(16) => OP_A_16_port, A(15) => n18, 
                           A(14) => OP_A_14_port, A(13) => OP_A_13_port, A(12) 
                           => OP_A_12_port, A(11) => OP_A_11_port, A(10) => 
                           OP_A_10_port, A(9) => OP_A_9_port, A(8) => 
                           OP_A_8_port, A(7) => OP_A_7_port, A(6) => 
                           OP_A_6_port, A(5) => OP_A_5_port, A(4) => 
                           OP_A_4_port, A(3) => OP_A_3_port, A(2) => 
                           OP_A_2_port, A(1) => OP_A_1_port, A(0) => 
                           OP_A_0_port, B(31) => OP_B_31_port, B(30) => 
                           OP_B_30_port, B(29) => OP_B_29_port, B(28) => 
                           OP_B_28_port, B(27) => OP_B_27_port, B(26) => 
                           OP_B_26_port, B(25) => OP_B_25_port, B(24) => 
                           OP_B_24_port, B(23) => OP_B_23_port, B(22) => 
                           OP_B_22_port, B(21) => OP_B_21_port, B(20) => 
                           OP_B_20_port, B(19) => OP_B_19_port, B(18) => 
                           OP_B_18_port, B(17) => OP_B_17_port, B(16) => 
                           OP_B_16_port, B(15) => OP_B_15_port, B(14) => 
                           OP_B_14_port, B(13) => OP_B_13_port, B(12) => 
                           OP_B_12_port, B(11) => OP_B_11_port, B(10) => 
                           OP_B_10_port, B(9) => OP_B_9_port, B(8) => 
                           OP_B_8_port, B(7) => OP_B_7_port, B(6) => 
                           OP_B_6_port, B(5) => OP_B_5_port, B(4) => n12, B(3) 
                           => n14, B(2) => n8, B(1) => n16, B(0) => n10, S(1) 
                           => OP_LOGIC_1_port, S(0) => OP_LOGIC_0_port, Y(31) 
                           => Y_LOGIC_31_port, Y(30) => Y_LOGIC_30_port, Y(29) 
                           => Y_LOGIC_29_port, Y(28) => Y_LOGIC_28_port, Y(27) 
                           => Y_LOGIC_27_port, Y(26) => Y_LOGIC_26_port, Y(25) 
                           => Y_LOGIC_25_port, Y(24) => Y_LOGIC_24_port, Y(23) 
                           => Y_LOGIC_23_port, Y(22) => Y_LOGIC_22_port, Y(21) 
                           => Y_LOGIC_21_port, Y(20) => Y_LOGIC_20_port, Y(19) 
                           => Y_LOGIC_19_port, Y(18) => Y_LOGIC_18_port, Y(17) 
                           => Y_LOGIC_17_port, Y(16) => Y_LOGIC_16_port, Y(15) 
                           => Y_LOGIC_15_port, Y(14) => Y_LOGIC_14_port, Y(13) 
                           => Y_LOGIC_13_port, Y(12) => Y_LOGIC_12_port, Y(11) 
                           => Y_LOGIC_11_port, Y(10) => Y_LOGIC_10_port, Y(9) 
                           => Y_LOGIC_9_port, Y(8) => Y_LOGIC_8_port, Y(7) => 
                           Y_LOGIC_7_port, Y(6) => Y_LOGIC_6_port, Y(5) => 
                           Y_LOGIC_5_port, Y(4) => Y_LOGIC_4_port, Y(3) => 
                           Y_LOGIC_3_port, Y(2) => Y_LOGIC_2_port, Y(1) => 
                           Y_LOGIC_1_port, Y(0) => Y_LOGIC_0_port);
   CMP : COMPARATOR_N32 port map( A(31) => OP_A_31_port, A(30) => OP_A_30_port,
                           A(29) => OP_A_29_port, A(28) => OP_A_28_port, A(27) 
                           => OP_A_27_port, A(26) => OP_A_26_port, A(25) => 
                           OP_A_25_port, A(24) => OP_A_24_port, A(23) => 
                           OP_A_23_port, A(22) => OP_A_22_port, A(21) => 
                           OP_A_21_port, A(20) => OP_A_20_port, A(19) => 
                           OP_A_19_port, A(18) => OP_A_18_port, A(17) => 
                           OP_A_17_port, A(16) => OP_A_16_port, A(15) => n18, 
                           A(14) => OP_A_14_port, A(13) => OP_A_13_port, A(12) 
                           => OP_A_12_port, A(11) => OP_A_11_port, A(10) => 
                           OP_A_10_port, A(9) => OP_A_9_port, A(8) => 
                           OP_A_8_port, A(7) => OP_A_7_port, A(6) => 
                           OP_A_6_port, A(5) => OP_A_5_port, A(4) => 
                           OP_A_4_port, A(3) => OP_A_3_port, A(2) => 
                           OP_A_2_port, A(1) => OP_A_1_port, A(0) => 
                           OP_A_0_port, B(31) => OP_B_31_port, B(30) => 
                           OP_B_30_port, B(29) => OP_B_29_port, B(28) => 
                           OP_B_28_port, B(27) => OP_B_27_port, B(26) => 
                           OP_B_26_port, B(25) => OP_B_25_port, B(24) => 
                           OP_B_24_port, B(23) => OP_B_23_port, B(22) => 
                           OP_B_22_port, B(21) => OP_B_21_port, B(20) => 
                           OP_B_20_port, B(19) => OP_B_19_port, B(18) => 
                           OP_B_18_port, B(17) => OP_B_17_port, B(16) => 
                           OP_B_16_port, B(15) => OP_B_15_port, B(14) => 
                           OP_B_14_port, B(13) => OP_B_13_port, B(12) => 
                           OP_B_12_port, B(11) => OP_B_11_port, B(10) => 
                           OP_B_10_port, B(9) => OP_B_9_port, B(8) => 
                           OP_B_8_port, B(7) => OP_B_7_port, B(6) => 
                           OP_B_6_port, B(5) => OP_B_5_port, B(4) => n12, B(3) 
                           => n14, B(2) => n8, B(1) => n16, B(0) => n10, S(3) 
                           => OP_COMPARE_3_port, S(2) => OP_COMPARE_2_port, 
                           S(1) => OP_COMPARE_1_port, S(0) => OP_COMPARE_0_port
                           , Y(31) => n_1285, Y(30) => n_1286, Y(29) => n_1287,
                           Y(28) => n_1288, Y(27) => n_1289, Y(26) => n_1290, 
                           Y(25) => n_1291, Y(24) => n_1292, Y(23) => n_1293, 
                           Y(22) => n_1294, Y(21) => n_1295, Y(20) => n_1296, 
                           Y(19) => n_1297, Y(18) => n_1298, Y(17) => n_1299, 
                           Y(16) => n_1300, Y(15) => n_1301, Y(14) => n_1302, 
                           Y(13) => n_1303, Y(12) => n_1304, Y(11) => n_1305, 
                           Y(10) => n_1306, Y(9) => n_1307, Y(8) => n_1308, 
                           Y(7) => n_1309, Y(6) => n_1310, Y(5) => n_1311, Y(4)
                           => n_1312, Y(3) => n_1313, Y(2) => n_1314, Y(1) => 
                           n_1315, Y(0) => Y_COMPARE_0_port);
   ZDET : ZERO_DETECTOR_N32_0 port map( A(31) => Y_31_port, A(30) => Y_30_port,
                           A(29) => Y_29_port, A(28) => Y_28_port, A(27) => 
                           Y_27_port, A(26) => Y_26_port, A(25) => Y_25_port, 
                           A(24) => Y_24_port, A(23) => Y_23_port, A(22) => 
                           Y_22_port, A(21) => Y_21_port, A(20) => Y_20_port, 
                           A(19) => Y_19_port, A(18) => Y_18_port, A(17) => 
                           Y_17_port, A(16) => Y_16_port, A(15) => Y_15_port, 
                           A(14) => Y_14_port, A(13) => Y_13_port, A(12) => 
                           Y_12_port, A(11) => Y_11_port, A(10) => Y_10_port, 
                           A(9) => Y_9_port, A(8) => Y_8_port, A(7) => Y_7_port
                           , A(6) => Y_6_port, A(5) => Y_5_port, A(4) => 
                           Y_4_port, A(3) => Y_3_port, A(2) => Y_2_port, A(1) 
                           => Y_1_port, A(0) => Y_0_port, Y => Z);
   OP_A_reg_0_inst : DLH_X2 port map( G => N246, D => OP1(0), Q => OP_A_0_port)
                           ;
   OP_A_reg_1_inst : DLH_X2 port map( G => N246, D => OP1(1), Q => OP_A_1_port)
                           ;
   OP_A_reg_7_inst : DLH_X2 port map( G => N246, D => OP1(7), Q => OP_A_7_port)
                           ;
   OP_A_reg_3_inst : DLH_X2 port map( G => N246, D => OP1(3), Q => OP_A_3_port)
                           ;
   OP_A_reg_11_inst : DLH_X2 port map( G => N246, D => OP1(11), Q => 
                           OP_A_11_port);
   OP_A_reg_14_inst : DLH_X2 port map( G => N246, D => OP1(14), Q => 
                           OP_A_14_port);
   OP_A_reg_10_inst : DLH_X2 port map( G => N246, D => OP1(10), Q => 
                           OP_A_10_port);
   OP_A_reg_6_inst : DLH_X2 port map( G => N246, D => OP1(6), Q => OP_A_6_port)
                           ;
   OP_A_reg_2_inst : DLH_X2 port map( G => N246, D => OP1(2), Q => OP_A_2_port)
                           ;
   OP_A_reg_8_inst : DLH_X2 port map( G => N246, D => OP1(8), Q => OP_A_8_port)
                           ;
   OP_A_reg_12_inst : DLH_X2 port map( G => N246, D => OP1(12), Q => 
                           OP_A_12_port);
   OP_A_reg_4_inst : DLH_X2 port map( G => N246, D => OP1(4), Q => OP_A_4_port)
                           ;
   U3 : OR2_X1 port map( A1 => n121, A2 => n122, ZN => n1);
   U4 : OR2_X1 port map( A1 => n119, A2 => n120, ZN => n2);
   U5 : INV_X2 port map( A => n2, ZN => n3);
   U6 : INV_X2 port map( A => n1, ZN => n4);
   U7 : INV_X1 port map( A => n24, ZN => n5);
   U8 : INV_X2 port map( A => n5, ZN => n6);
   U9 : NAND2_X2 port map( A1 => n139, A2 => n144, ZN => N246);
   U10 : INV_X1 port map( A => OP_B_2_port, ZN => n7);
   U11 : INV_X4 port map( A => n7, ZN => n8);
   U12 : INV_X1 port map( A => OP_B_0_port, ZN => n9);
   U13 : INV_X4 port map( A => n9, ZN => n10);
   U14 : INV_X1 port map( A => OP_B_4_port, ZN => n11);
   U15 : INV_X4 port map( A => n11, ZN => n12);
   U16 : INV_X1 port map( A => OP_B_3_port, ZN => n13);
   U17 : INV_X4 port map( A => n13, ZN => n14);
   U18 : INV_X1 port map( A => OP_B_1_port, ZN => n15);
   U19 : INV_X4 port map( A => n15, ZN => n16);
   U20 : INV_X1 port map( A => OP_A_15_port, ZN => n17);
   U21 : INV_X8 port map( A => n17, ZN => n18);
   U22 : NAND4_X2 port map( A1 => n139, A2 => n140, A3 => n141, A4 => n142, ZN 
                           => n138);
   U23 : INV_X2 port map( A => n225, ZN => n22);
   U24 : AND4_X2 port map( A1 => OPC(1), A2 => n167, A3 => n168, A4 => n150, ZN
                           => n23);
   U25 : OR3_X2 port map( A1 => n183, A2 => n182, A3 => n181, ZN => N281);
   U26 : NAND4_X2 port map( A1 => n140, A2 => n141, A3 => n142, A4 => n143, ZN 
                           => N279);
   U27 : NAND3_X1 port map( A1 => n19, A2 => n20, A3 => n21, ZN => Y_9_port);
   U28 : AOI222_X1 port map( A1 => Y_SHIFTR_9_port, A2 => n22, B1 => 
                           Y_SUM_9_port, B2 => N279, C1 => Y_LOGIC_9_port, C2 
                           => N281, ZN => n21);
   U29 : AOI22_X1 port map( A1 => OP2(9), A2 => n4, B1 => OP1(9), B2 => n3, ZN 
                           => n20);
   U30 : AOI22_X1 port map( A1 => Y_MUL_9_port, A2 => n23, B1 => 
                           Y_SHIFTL_9_port, B2 => n6, ZN => n19);
   U31 : NAND3_X1 port map( A1 => n25, A2 => n26, A3 => n27, ZN => Y_8_port);
   U32 : AOI222_X1 port map( A1 => Y_SHIFTR_8_port, A2 => n22, B1 => 
                           Y_SUM_8_port, B2 => N279, C1 => Y_LOGIC_8_port, C2 
                           => N281, ZN => n27);
   U33 : AOI22_X1 port map( A1 => OP2(8), A2 => n4, B1 => OP1(8), B2 => n3, ZN 
                           => n26);
   U34 : AOI22_X1 port map( A1 => Y_MUL_8_port, A2 => n23, B1 => 
                           Y_SHIFTL_8_port, B2 => n6, ZN => n25);
   U35 : NAND3_X1 port map( A1 => n28, A2 => n29, A3 => n30, ZN => Y_7_port);
   U36 : AOI222_X1 port map( A1 => Y_SHIFTR_7_port, A2 => n22, B1 => 
                           Y_SUM_7_port, B2 => N279, C1 => Y_LOGIC_7_port, C2 
                           => N281, ZN => n30);
   U37 : AOI22_X1 port map( A1 => OP2(7), A2 => n4, B1 => OP1(7), B2 => n3, ZN 
                           => n29);
   U38 : AOI22_X1 port map( A1 => Y_MUL_7_port, A2 => n23, B1 => 
                           Y_SHIFTL_7_port, B2 => n6, ZN => n28);
   U39 : NAND3_X1 port map( A1 => n31, A2 => n32, A3 => n33, ZN => Y_6_port);
   U40 : AOI222_X1 port map( A1 => Y_SHIFTR_6_port, A2 => n22, B1 => 
                           Y_SUM_6_port, B2 => N279, C1 => Y_LOGIC_6_port, C2 
                           => N281, ZN => n33);
   U41 : AOI22_X1 port map( A1 => OP2(6), A2 => n4, B1 => OP1(6), B2 => n3, ZN 
                           => n32);
   U42 : AOI22_X1 port map( A1 => Y_MUL_6_port, A2 => n23, B1 => 
                           Y_SHIFTL_6_port, B2 => n6, ZN => n31);
   U43 : NAND3_X1 port map( A1 => n34, A2 => n35, A3 => n36, ZN => Y_5_port);
   U44 : AOI222_X1 port map( A1 => Y_SHIFTR_5_port, A2 => n22, B1 => 
                           Y_SUM_5_port, B2 => N279, C1 => Y_LOGIC_5_port, C2 
                           => N281, ZN => n36);
   U45 : AOI22_X1 port map( A1 => OP2(5), A2 => n4, B1 => OP1(5), B2 => n3, ZN 
                           => n35);
   U46 : AOI22_X1 port map( A1 => Y_MUL_5_port, A2 => n23, B1 => 
                           Y_SHIFTL_5_port, B2 => n6, ZN => n34);
   U47 : NAND3_X1 port map( A1 => n37, A2 => n38, A3 => n39, ZN => Y_4_port);
   U48 : AOI222_X1 port map( A1 => Y_SHIFTR_4_port, A2 => n22, B1 => 
                           Y_SUM_4_port, B2 => N279, C1 => Y_LOGIC_4_port, C2 
                           => N281, ZN => n39);
   U49 : AOI22_X1 port map( A1 => OP2(4), A2 => n4, B1 => OP1(4), B2 => n3, ZN 
                           => n38);
   U50 : AOI22_X1 port map( A1 => Y_MUL_4_port, A2 => n23, B1 => 
                           Y_SHIFTL_4_port, B2 => n6, ZN => n37);
   U51 : NAND3_X1 port map( A1 => n40, A2 => n41, A3 => n42, ZN => Y_3_port);
   U52 : AOI222_X1 port map( A1 => Y_SHIFTR_3_port, A2 => n22, B1 => 
                           Y_SUM_3_port, B2 => N279, C1 => Y_LOGIC_3_port, C2 
                           => N281, ZN => n42);
   U53 : AOI22_X1 port map( A1 => OP2(3), A2 => n4, B1 => OP1(3), B2 => n3, ZN 
                           => n41);
   U54 : AOI22_X1 port map( A1 => Y_MUL_3_port, A2 => n23, B1 => 
                           Y_SHIFTL_3_port, B2 => n6, ZN => n40);
   U55 : NAND3_X1 port map( A1 => n43, A2 => n44, A3 => n45, ZN => Y_31_port);
   U56 : AOI222_X1 port map( A1 => Y_SHIFTR_31_port, A2 => n22, B1 => 
                           Y_SUM_31_port, B2 => N279, C1 => Y_LOGIC_31_port, C2
                           => N281, ZN => n45);
   U57 : AOI22_X1 port map( A1 => OP2(31), A2 => n4, B1 => OP1(31), B2 => n3, 
                           ZN => n44);
   U58 : AOI22_X1 port map( A1 => Y_MUL_31_port, A2 => n23, B1 => 
                           Y_SHIFTL_31_port, B2 => n6, ZN => n43);
   U59 : NAND3_X1 port map( A1 => n46, A2 => n47, A3 => n48, ZN => Y_30_port);
   U60 : AOI222_X1 port map( A1 => Y_SHIFTR_30_port, A2 => n22, B1 => 
                           Y_SUM_30_port, B2 => N279, C1 => Y_LOGIC_30_port, C2
                           => N281, ZN => n48);
   U61 : AOI22_X1 port map( A1 => OP2(30), A2 => n4, B1 => OP1(30), B2 => n3, 
                           ZN => n47);
   U62 : AOI22_X1 port map( A1 => Y_MUL_30_port, A2 => n23, B1 => 
                           Y_SHIFTL_30_port, B2 => n6, ZN => n46);
   U63 : NAND3_X1 port map( A1 => n49, A2 => n50, A3 => n51, ZN => Y_2_port);
   U64 : AOI222_X1 port map( A1 => Y_SHIFTR_2_port, A2 => n22, B1 => 
                           Y_SUM_2_port, B2 => N279, C1 => Y_LOGIC_2_port, C2 
                           => N281, ZN => n51);
   U65 : AOI22_X1 port map( A1 => OP2(2), A2 => n4, B1 => OP1(2), B2 => n3, ZN 
                           => n50);
   U66 : AOI22_X1 port map( A1 => Y_MUL_2_port, A2 => n23, B1 => 
                           Y_SHIFTL_2_port, B2 => n6, ZN => n49);
   U67 : NAND3_X1 port map( A1 => n52, A2 => n53, A3 => n54, ZN => Y_29_port);
   U68 : AOI222_X1 port map( A1 => Y_SHIFTR_29_port, A2 => n22, B1 => 
                           Y_SUM_29_port, B2 => N279, C1 => Y_LOGIC_29_port, C2
                           => N281, ZN => n54);
   U69 : AOI22_X1 port map( A1 => OP2(29), A2 => n4, B1 => OP1(29), B2 => n3, 
                           ZN => n53);
   U70 : AOI22_X1 port map( A1 => Y_MUL_29_port, A2 => n23, B1 => 
                           Y_SHIFTL_29_port, B2 => n6, ZN => n52);
   U71 : NAND3_X1 port map( A1 => n55, A2 => n56, A3 => n57, ZN => Y_28_port);
   U72 : AOI222_X1 port map( A1 => Y_SHIFTR_28_port, A2 => n22, B1 => 
                           Y_SUM_28_port, B2 => N279, C1 => Y_LOGIC_28_port, C2
                           => N281, ZN => n57);
   U73 : AOI22_X1 port map( A1 => OP2(28), A2 => n4, B1 => OP1(28), B2 => n3, 
                           ZN => n56);
   U74 : AOI22_X1 port map( A1 => Y_MUL_28_port, A2 => n23, B1 => 
                           Y_SHIFTL_28_port, B2 => n6, ZN => n55);
   U75 : NAND3_X1 port map( A1 => n58, A2 => n59, A3 => n60, ZN => Y_27_port);
   U76 : AOI222_X1 port map( A1 => Y_SHIFTR_27_port, A2 => n22, B1 => 
                           Y_SUM_27_port, B2 => N279, C1 => Y_LOGIC_27_port, C2
                           => N281, ZN => n60);
   U77 : AOI22_X1 port map( A1 => OP2(27), A2 => n4, B1 => OP1(27), B2 => n3, 
                           ZN => n59);
   U78 : AOI22_X1 port map( A1 => Y_MUL_27_port, A2 => n23, B1 => 
                           Y_SHIFTL_27_port, B2 => n6, ZN => n58);
   U79 : NAND3_X1 port map( A1 => n61, A2 => n62, A3 => n63, ZN => Y_26_port);
   U80 : AOI222_X1 port map( A1 => Y_SHIFTR_26_port, A2 => n22, B1 => 
                           Y_SUM_26_port, B2 => N279, C1 => Y_LOGIC_26_port, C2
                           => N281, ZN => n63);
   U81 : AOI22_X1 port map( A1 => OP2(26), A2 => n4, B1 => OP1(26), B2 => n3, 
                           ZN => n62);
   U82 : AOI22_X1 port map( A1 => Y_MUL_26_port, A2 => n23, B1 => 
                           Y_SHIFTL_26_port, B2 => n6, ZN => n61);
   U83 : NAND3_X1 port map( A1 => n64, A2 => n65, A3 => n66, ZN => Y_25_port);
   U84 : AOI222_X1 port map( A1 => Y_SHIFTR_25_port, A2 => n22, B1 => 
                           Y_SUM_25_port, B2 => N279, C1 => Y_LOGIC_25_port, C2
                           => N281, ZN => n66);
   U85 : AOI22_X1 port map( A1 => OP2(25), A2 => n4, B1 => OP1(25), B2 => n3, 
                           ZN => n65);
   U86 : AOI22_X1 port map( A1 => Y_MUL_25_port, A2 => n23, B1 => 
                           Y_SHIFTL_25_port, B2 => n6, ZN => n64);
   U87 : NAND3_X1 port map( A1 => n67, A2 => n68, A3 => n69, ZN => Y_24_port);
   U88 : AOI222_X1 port map( A1 => Y_SHIFTR_24_port, A2 => n22, B1 => 
                           Y_SUM_24_port, B2 => N279, C1 => Y_LOGIC_24_port, C2
                           => N281, ZN => n69);
   U89 : AOI22_X1 port map( A1 => OP2(24), A2 => n4, B1 => OP1(24), B2 => n3, 
                           ZN => n68);
   U90 : AOI22_X1 port map( A1 => Y_MUL_24_port, A2 => n23, B1 => 
                           Y_SHIFTL_24_port, B2 => n6, ZN => n67);
   U91 : NAND3_X1 port map( A1 => n70, A2 => n71, A3 => n72, ZN => Y_23_port);
   U92 : AOI222_X1 port map( A1 => Y_SHIFTR_23_port, A2 => n22, B1 => 
                           Y_SUM_23_port, B2 => N279, C1 => Y_LOGIC_23_port, C2
                           => N281, ZN => n72);
   U93 : AOI22_X1 port map( A1 => OP2(23), A2 => n4, B1 => OP1(23), B2 => n3, 
                           ZN => n71);
   U94 : AOI22_X1 port map( A1 => Y_MUL_23_port, A2 => n23, B1 => 
                           Y_SHIFTL_23_port, B2 => n6, ZN => n70);
   U95 : NAND3_X1 port map( A1 => n73, A2 => n74, A3 => n75, ZN => Y_22_port);
   U96 : AOI222_X1 port map( A1 => Y_SHIFTR_22_port, A2 => n22, B1 => 
                           Y_SUM_22_port, B2 => N279, C1 => Y_LOGIC_22_port, C2
                           => N281, ZN => n75);
   U97 : AOI22_X1 port map( A1 => OP2(22), A2 => n4, B1 => OP1(22), B2 => n3, 
                           ZN => n74);
   U98 : AOI22_X1 port map( A1 => Y_MUL_22_port, A2 => n23, B1 => 
                           Y_SHIFTL_22_port, B2 => n6, ZN => n73);
   U99 : NAND3_X1 port map( A1 => n76, A2 => n77, A3 => n78, ZN => Y_21_port);
   U100 : AOI222_X1 port map( A1 => Y_SHIFTR_21_port, A2 => n22, B1 => 
                           Y_SUM_21_port, B2 => N279, C1 => Y_LOGIC_21_port, C2
                           => N281, ZN => n78);
   U101 : AOI22_X1 port map( A1 => OP2(21), A2 => n4, B1 => OP1(21), B2 => n3, 
                           ZN => n77);
   U102 : AOI22_X1 port map( A1 => Y_MUL_21_port, A2 => n23, B1 => 
                           Y_SHIFTL_21_port, B2 => n6, ZN => n76);
   U103 : NAND3_X1 port map( A1 => n79, A2 => n80, A3 => n81, ZN => Y_20_port);
   U104 : AOI222_X1 port map( A1 => Y_SHIFTR_20_port, A2 => n22, B1 => 
                           Y_SUM_20_port, B2 => N279, C1 => Y_LOGIC_20_port, C2
                           => N281, ZN => n81);
   U105 : AOI22_X1 port map( A1 => OP2(20), A2 => n4, B1 => OP1(20), B2 => n3, 
                           ZN => n80);
   U106 : AOI22_X1 port map( A1 => Y_MUL_20_port, A2 => n23, B1 => 
                           Y_SHIFTL_20_port, B2 => n6, ZN => n79);
   U107 : NAND3_X1 port map( A1 => n82, A2 => n83, A3 => n84, ZN => Y_1_port);
   U108 : AOI222_X1 port map( A1 => Y_SHIFTR_1_port, A2 => n22, B1 => 
                           Y_SUM_1_port, B2 => N279, C1 => Y_LOGIC_1_port, C2 
                           => N281, ZN => n84);
   U109 : AOI22_X1 port map( A1 => OP2(1), A2 => n4, B1 => OP1(1), B2 => n3, ZN
                           => n83);
   U110 : AOI22_X1 port map( A1 => Y_MUL_1_port, A2 => n23, B1 => 
                           Y_SHIFTL_1_port, B2 => n6, ZN => n82);
   U111 : NAND3_X1 port map( A1 => n85, A2 => n86, A3 => n87, ZN => Y_19_port);
   U112 : AOI222_X1 port map( A1 => Y_SHIFTR_19_port, A2 => n22, B1 => 
                           Y_SUM_19_port, B2 => N279, C1 => Y_LOGIC_19_port, C2
                           => N281, ZN => n87);
   U113 : AOI22_X1 port map( A1 => OP2(19), A2 => n4, B1 => OP1(19), B2 => n3, 
                           ZN => n86);
   U114 : AOI22_X1 port map( A1 => Y_MUL_19_port, A2 => n23, B1 => 
                           Y_SHIFTL_19_port, B2 => n6, ZN => n85);
   U115 : NAND3_X1 port map( A1 => n88, A2 => n89, A3 => n90, ZN => Y_18_port);
   U116 : AOI222_X1 port map( A1 => Y_SHIFTR_18_port, A2 => n22, B1 => 
                           Y_SUM_18_port, B2 => N279, C1 => Y_LOGIC_18_port, C2
                           => N281, ZN => n90);
   U117 : AOI22_X1 port map( A1 => OP2(18), A2 => n4, B1 => OP1(18), B2 => n3, 
                           ZN => n89);
   U118 : AOI22_X1 port map( A1 => Y_MUL_18_port, A2 => n23, B1 => 
                           Y_SHIFTL_18_port, B2 => n6, ZN => n88);
   U119 : NAND3_X1 port map( A1 => n91, A2 => n92, A3 => n93, ZN => Y_17_port);
   U120 : AOI222_X1 port map( A1 => Y_SHIFTR_17_port, A2 => n22, B1 => 
                           Y_SUM_17_port, B2 => N279, C1 => Y_LOGIC_17_port, C2
                           => N281, ZN => n93);
   U121 : AOI22_X1 port map( A1 => OP2(17), A2 => n4, B1 => OP1(17), B2 => n3, 
                           ZN => n92);
   U122 : AOI22_X1 port map( A1 => Y_MUL_17_port, A2 => n23, B1 => 
                           Y_SHIFTL_17_port, B2 => n6, ZN => n91);
   U123 : NAND3_X1 port map( A1 => n94, A2 => n95, A3 => n96_port, ZN => 
                           Y_16_port);
   U124 : AOI222_X1 port map( A1 => Y_SHIFTR_16_port, A2 => n22, B1 => 
                           Y_SUM_16_port, B2 => N279, C1 => Y_LOGIC_16_port, C2
                           => N281, ZN => n96_port);
   U125 : AOI22_X1 port map( A1 => OP2(16), A2 => n4, B1 => OP1(16), B2 => n3, 
                           ZN => n95);
   U126 : AOI22_X1 port map( A1 => Y_MUL_16_port, A2 => n23, B1 => 
                           Y_SHIFTL_16_port, B2 => n6, ZN => n94);
   U127 : NAND3_X1 port map( A1 => n97, A2 => n98, A3 => n99, ZN => Y_15_port);
   U128 : AOI222_X1 port map( A1 => Y_SHIFTR_15_port, A2 => n22, B1 => 
                           Y_SUM_15_port, B2 => N279, C1 => Y_LOGIC_15_port, C2
                           => N281, ZN => n99);
   U129 : AOI22_X1 port map( A1 => OP2(15), A2 => n4, B1 => OP1(15), B2 => n3, 
                           ZN => n98);
   U130 : AOI22_X1 port map( A1 => Y_MUL_15_port, A2 => n23, B1 => 
                           Y_SHIFTL_15_port, B2 => n6, ZN => n97);
   U131 : NAND3_X1 port map( A1 => n100, A2 => n101, A3 => n102, ZN => 
                           Y_14_port);
   U132 : AOI222_X1 port map( A1 => Y_SHIFTR_14_port, A2 => n22, B1 => 
                           Y_SUM_14_port, B2 => N279, C1 => Y_LOGIC_14_port, C2
                           => N281, ZN => n102);
   U133 : AOI22_X1 port map( A1 => OP2(14), A2 => n4, B1 => OP1(14), B2 => n3, 
                           ZN => n101);
   U134 : AOI22_X1 port map( A1 => Y_MUL_14_port, A2 => n23, B1 => 
                           Y_SHIFTL_14_port, B2 => n6, ZN => n100);
   U135 : NAND3_X1 port map( A1 => n103, A2 => n104, A3 => n105, ZN => 
                           Y_13_port);
   U136 : AOI222_X1 port map( A1 => Y_SHIFTR_13_port, A2 => n22, B1 => 
                           Y_SUM_13_port, B2 => N279, C1 => Y_LOGIC_13_port, C2
                           => N281, ZN => n105);
   U137 : AOI22_X1 port map( A1 => OP2(13), A2 => n4, B1 => OP1(13), B2 => n3, 
                           ZN => n104);
   U138 : AOI22_X1 port map( A1 => Y_MUL_13_port, A2 => n23, B1 => 
                           Y_SHIFTL_13_port, B2 => n6, ZN => n103);
   U139 : NAND3_X1 port map( A1 => n106, A2 => n107, A3 => n108, ZN => 
                           Y_12_port);
   U140 : AOI222_X1 port map( A1 => Y_SHIFTR_12_port, A2 => n22, B1 => 
                           Y_SUM_12_port, B2 => N279, C1 => Y_LOGIC_12_port, C2
                           => N281, ZN => n108);
   U141 : AOI22_X1 port map( A1 => OP2(12), A2 => n4, B1 => OP1(12), B2 => n3, 
                           ZN => n107);
   U142 : AOI22_X1 port map( A1 => Y_MUL_12_port, A2 => n23, B1 => 
                           Y_SHIFTL_12_port, B2 => n6, ZN => n106);
   U143 : NAND3_X1 port map( A1 => n109, A2 => n110, A3 => n111, ZN => 
                           Y_11_port);
   U144 : AOI222_X1 port map( A1 => Y_SHIFTR_11_port, A2 => n22, B1 => 
                           Y_SUM_11_port, B2 => N279, C1 => Y_LOGIC_11_port, C2
                           => N281, ZN => n111);
   U145 : AOI22_X1 port map( A1 => OP2(11), A2 => n4, B1 => OP1(11), B2 => n3, 
                           ZN => n110);
   U146 : AOI22_X1 port map( A1 => Y_MUL_11_port, A2 => n23, B1 => 
                           Y_SHIFTL_11_port, B2 => n6, ZN => n109);
   U147 : NAND3_X1 port map( A1 => n112, A2 => n113, A3 => n114, ZN => 
                           Y_10_port);
   U148 : AOI222_X1 port map( A1 => Y_SHIFTR_10_port, A2 => n22, B1 => 
                           Y_SUM_10_port, B2 => N279, C1 => Y_LOGIC_10_port, C2
                           => N281, ZN => n114);
   U149 : AOI22_X1 port map( A1 => OP2(10), A2 => n4, B1 => OP1(10), B2 => n3, 
                           ZN => n113);
   U150 : AOI22_X1 port map( A1 => Y_MUL_10_port, A2 => n23, B1 => 
                           Y_SHIFTL_10_port, B2 => n6, ZN => n112);
   U151 : NAND4_X1 port map( A1 => n115, A2 => n116, A3 => n117, A4 => n118, ZN
                           => Y_0_port);
   U152 : AOI22_X1 port map( A1 => OP2(0), A2 => n4, B1 => OP1(0), B2 => n3, ZN
                           => n118);
   U153 : AOI22_X1 port map( A1 => Y_MUL_0_port, A2 => n23, B1 => 
                           Y_SHIFTL_0_port, B2 => n6, ZN => n117);
   U154 : AOI22_X1 port map( A1 => Y_SUM_0_port, A2 => N279, B1 => 
                           Y_LOGIC_0_port, B2 => N281, ZN => n116);
   U155 : AOI22_X1 port map( A1 => Y_COMPARE_0_port, A2 => N285, B1 => 
                           Y_SHIFTR_0_port, B2 => n22, ZN => n115);
   U156 : OAI21_X1 port map( B1 => n123, B2 => n124, A => n125, ZN => N289);
   U157 : OAI211_X1 port map( C1 => n123, C2 => n126, A => n127, B => n128, ZN 
                           => N288);
   U158 : OAI211_X1 port map( C1 => n129, C2 => n130, A => n131, B => n132, ZN 
                           => N287);
   U159 : AOI221_X1 port map( B1 => n133, B2 => n134, C1 => n135, C2 => n136, A
                           => n137, ZN => n132);
   U160 : MUX2_X1 port map( A => N280, B => n138, S => OP2(31), Z => N278);
   U161 : MUX2_X1 port map( A => N280, B => n138, S => OP2(30), Z => N277);
   U162 : MUX2_X1 port map( A => N280, B => n138, S => OP2(29), Z => N276);
   U163 : MUX2_X1 port map( A => N280, B => n138, S => OP2(28), Z => N275);
   U164 : MUX2_X1 port map( A => N280, B => n138, S => OP2(27), Z => N274);
   U165 : MUX2_X1 port map( A => N280, B => n138, S => OP2(26), Z => N273);
   U166 : MUX2_X1 port map( A => N280, B => n138, S => OP2(25), Z => N272);
   U167 : MUX2_X1 port map( A => N280, B => n138, S => OP2(24), Z => N271);
   U168 : MUX2_X1 port map( A => N280, B => n138, S => OP2(23), Z => N270);
   U169 : MUX2_X1 port map( A => N280, B => n138, S => OP2(22), Z => N269);
   U170 : MUX2_X1 port map( A => N280, B => n138, S => OP2(21), Z => N268);
   U171 : MUX2_X1 port map( A => N280, B => n138, S => OP2(20), Z => N267);
   U172 : MUX2_X1 port map( A => N280, B => n138, S => OP2(19), Z => N266);
   U173 : MUX2_X1 port map( A => N280, B => n138, S => OP2(18), Z => N265);
   U174 : MUX2_X1 port map( A => N280, B => n138, S => OP2(17), Z => N264);
   U175 : MUX2_X1 port map( A => N280, B => n138, S => OP2(16), Z => N263);
   U176 : MUX2_X1 port map( A => N280, B => n138, S => OP2(15), Z => N262);
   U177 : MUX2_X1 port map( A => N280, B => n138, S => OP2(14), Z => N261);
   U178 : MUX2_X1 port map( A => N280, B => n138, S => OP2(13), Z => N260);
   U179 : MUX2_X1 port map( A => N280, B => n138, S => OP2(12), Z => N259);
   U180 : MUX2_X1 port map( A => N280, B => n138, S => OP2(11), Z => N258);
   U181 : MUX2_X1 port map( A => N280, B => n138, S => OP2(10), Z => N257);
   U182 : MUX2_X1 port map( A => N280, B => n138, S => OP2(9), Z => N256);
   U183 : MUX2_X1 port map( A => N280, B => n138, S => OP2(8), Z => N255);
   U184 : MUX2_X1 port map( A => N280, B => n138, S => OP2(7), Z => N254);
   U185 : MUX2_X1 port map( A => N280, B => n138, S => OP2(6), Z => N253);
   U186 : MUX2_X1 port map( A => N280, B => n138, S => OP2(5), Z => N252);
   U187 : MUX2_X1 port map( A => N280, B => n138, S => OP2(4), Z => N251);
   U188 : MUX2_X1 port map( A => N280, B => n138, S => OP2(3), Z => N250);
   U189 : MUX2_X1 port map( A => N280, B => n138, S => OP2(2), Z => N249);
   U190 : MUX2_X1 port map( A => N280, B => n138, S => OP2(1), Z => N248);
   U191 : MUX2_X1 port map( A => N280, B => n138, S => OP2(0), Z => N247);
   U192 : INV_X1 port map( A => n143, ZN => N280);
   U193 : INV_X1 port map( A => N279, ZN => n144);
   U194 : AOI22_X1 port map( A1 => n145, A2 => n146, B1 => n147, B2 => n148, ZN
                           => n143);
   U195 : INV_X1 port map( A => n122, ZN => n146);
   U196 : NAND4_X1 port map( A1 => n149, A2 => n150, A3 => OPC(3), A4 => n151, 
                           ZN => n142);
   U197 : NOR2_X1 port map( A1 => n152, A2 => n153, ZN => n151);
   U198 : NAND4_X1 port map( A1 => n154, A2 => n124, A3 => n155, A4 => n130, ZN
                           => n149);
   U199 : OAI21_X1 port map( B1 => n133, B2 => n156, A => n157, ZN => n141);
   U200 : INV_X1 port map( A => n158, ZN => n140);
   U201 : OAI22_X1 port map( A1 => n124, A2 => n159, B1 => n160, B2 => n161, ZN
                           => n158);
   U202 : AOI211_X1 port map( C1 => n162, C2 => OPC(3), A => n156, B => n148, 
                           ZN => n160);
   U203 : NOR4_X1 port map( A1 => N281, A2 => N285, A3 => n23, A4 => n163, ZN 
                           => n139);
   U204 : OR2_X1 port map( A1 => n6, A2 => n22, ZN => n163);
   U205 : AOI221_X1 port map( B1 => n164, B2 => n165, C1 => n134, C2 => n148, A
                           => N96, ZN => n225);
   U206 : OAI22_X1 port map( A1 => n159, A2 => n154, B1 => n161, B2 => n119, ZN
                           => N96);
   U207 : OAI22_X1 port map( A1 => n119, A2 => n154, B1 => n166, B2 => n159, ZN
                           => n24);
   U208 : XNOR2_X1 port map( A => n152, B => OPC(3), ZN => n168);
   U209 : NAND4_X1 port map( A1 => n131, A2 => n128, A3 => n125, A4 => n169, ZN
                           => N285);
   U210 : AOI221_X1 port map( B1 => n157, B2 => n165, C1 => n167, C2 => n170, A
                           => N286, ZN => n169);
   U211 : NAND3_X1 port map( A1 => n171, A2 => n127, A3 => n172, ZN => N286);
   U212 : INV_X1 port map( A => n173, ZN => n172);
   U213 : OAI22_X1 port map( A1 => n124, A2 => n129, B1 => n130, B2 => n119, ZN
                           => n173);
   U214 : INV_X1 port map( A => n137, ZN => n127);
   U215 : NOR2_X1 port map( A1 => n154, A2 => n123, ZN => n137);
   U216 : OAI21_X1 port map( B1 => n164, B2 => n145, A => n136, ZN => n171);
   U217 : INV_X1 port map( A => n123, ZN => n136);
   U218 : AOI21_X1 port map( B1 => n174, B2 => OPC(2), A => n156, ZN => n123);
   U219 : NOR4_X1 port map( A1 => n153, A2 => n150, A3 => OPC(3), A4 => OPC(2),
                           ZN => n156);
   U220 : INV_X1 port map( A => OPC(1), ZN => n153);
   U221 : INV_X1 port map( A => n121, ZN => n157);
   U222 : AOI22_X1 port map( A1 => n167, A2 => n133, B1 => n170, B2 => n175, ZN
                           => n125);
   U223 : AOI22_X1 port map( A1 => n145, A2 => n133, B1 => n147, B2 => n170, ZN
                           => n128);
   U224 : NAND2_X1 port map( A1 => n121, A2 => n130, ZN => n147);
   U225 : NAND3_X1 port map( A1 => OPC(4), A2 => n176, A3 => OPC(5), ZN => n130
                           );
   U226 : NAND3_X1 port map( A1 => OPC(4), A2 => n177, A3 => OPC(6), ZN => n121
                           );
   U227 : AND2_X1 port map( A1 => n162, A2 => n178, ZN => n133);
   U228 : NOR3_X1 port map( A1 => n150, A2 => OPC(1), A3 => n152, ZN => n162);
   U229 : INV_X1 port map( A => n120, ZN => n145);
   U230 : NOR2_X1 port map( A1 => n135, A2 => n134, ZN => n120);
   U231 : AOI22_X1 port map( A1 => n165, A2 => n175, B1 => n179, B2 => n170, ZN
                           => n131);
   U232 : INV_X1 port map( A => n129, ZN => n170);
   U233 : INV_X1 port map( A => n161, ZN => n179);
   U234 : INV_X1 port map( A => n155, ZN => n175);
   U235 : INV_X1 port map( A => n119, ZN => n165);
   U236 : NAND2_X1 port map( A1 => OPC(3), A2 => n180, ZN => n119);
   U237 : OAI22_X1 port map( A1 => n154, A2 => n122, B1 => n155, B2 => n159, ZN
                           => n181);
   U238 : INV_X1 port map( A => n148, ZN => n159);
   U239 : NOR4_X1 port map( A1 => OPC(3), A2 => OPC(2), A3 => OPC(1), A4 => 
                           OPC(0), ZN => n148);
   U240 : NAND3_X1 port map( A1 => OPC(6), A2 => OPC(4), A3 => OPC(5), ZN => 
                           n155);
   U241 : INV_X1 port map( A => n167, ZN => n154);
   U242 : NOR3_X1 port map( A1 => OPC(6), A2 => OPC(4), A3 => n177, ZN => n167)
                           ;
   U243 : OAI22_X1 port map( A1 => n126, A2 => n129, B1 => n122, B2 => n161, ZN
                           => n182);
   U244 : NAND3_X1 port map( A1 => n176, A2 => n177, A3 => OPC(4), ZN => n161);
   U245 : INV_X1 port map( A => n134, ZN => n126);
   U246 : NOR3_X1 port map( A1 => OPC(5), A2 => OPC(4), A3 => n176, ZN => n134)
                           ;
   U247 : OAI22_X1 port map( A1 => n129, A2 => n166, B1 => n122, B2 => n124, ZN
                           => n183);
   U248 : INV_X1 port map( A => n164, ZN => n124);
   U249 : NOR3_X1 port map( A1 => n176, A2 => OPC(4), A3 => n177, ZN => n164);
   U250 : INV_X1 port map( A => OPC(5), ZN => n177);
   U251 : INV_X1 port map( A => OPC(6), ZN => n176);
   U252 : NAND2_X1 port map( A1 => n180, A2 => n178, ZN => n122);
   U253 : NOR3_X1 port map( A1 => OPC(2), A2 => OPC(1), A3 => n150, ZN => n180)
                           ;
   U254 : INV_X1 port map( A => OPC(0), ZN => n150);
   U255 : INV_X1 port map( A => n135, ZN => n166);
   U256 : NOR3_X1 port map( A1 => OPC(5), A2 => OPC(4), A3 => OPC(6), ZN => 
                           n135);
   U257 : NAND2_X1 port map( A1 => n174, A2 => n152, ZN => n129);
   U258 : INV_X1 port map( A => OPC(2), ZN => n152);
   U259 : NOR3_X1 port map( A1 => OPC(1), A2 => OPC(0), A3 => n178, ZN => n174)
                           ;
   U260 : INV_X1 port map( A => OPC(3), ZN => n178);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX41_N32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX41_N32_1;

architecture SYN_BEHAVIORAL of MUX41_N32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n1);
   U2 : OR2_X1 port map( A1 => n71, A2 => S(1), ZN => n2);
   U3 : INV_X2 port map( A => n2, ZN => n3);
   U4 : INV_X2 port map( A => n1, ZN => n4);
   U5 : AND2_X2 port map( A1 => S(0), A2 => S(1), ZN => n8);
   U6 : AND2_X2 port map( A1 => S(1), A2 => n71, ZN => n7);
   U7 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Y(9));
   U8 : AOI22_X1 port map( A1 => C(9), A2 => n7, B1 => D(9), B2 => n8, ZN => n6
                           );
   U9 : AOI22_X1 port map( A1 => A(9), A2 => n4, B1 => B(9), B2 => n3, ZN => n5
                           );
   U10 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => Y(8));
   U11 : AOI22_X1 port map( A1 => C(8), A2 => n7, B1 => D(8), B2 => n8, ZN => 
                           n10);
   U12 : AOI22_X1 port map( A1 => A(8), A2 => n4, B1 => B(8), B2 => n3, ZN => 
                           n9);
   U13 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => Y(7));
   U14 : AOI22_X1 port map( A1 => C(7), A2 => n7, B1 => D(7), B2 => n8, ZN => 
                           n12);
   U15 : AOI22_X1 port map( A1 => A(7), A2 => n4, B1 => B(7), B2 => n3, ZN => 
                           n11);
   U16 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => Y(6));
   U17 : AOI22_X1 port map( A1 => C(6), A2 => n7, B1 => D(6), B2 => n8, ZN => 
                           n14);
   U18 : AOI22_X1 port map( A1 => A(6), A2 => n4, B1 => B(6), B2 => n3, ZN => 
                           n13);
   U19 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => Y(5));
   U20 : AOI22_X1 port map( A1 => C(5), A2 => n7, B1 => D(5), B2 => n8, ZN => 
                           n16);
   U21 : AOI22_X1 port map( A1 => A(5), A2 => n4, B1 => B(5), B2 => n3, ZN => 
                           n15);
   U22 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => Y(4));
   U23 : AOI22_X1 port map( A1 => C(4), A2 => n7, B1 => D(4), B2 => n8, ZN => 
                           n18);
   U24 : AOI22_X1 port map( A1 => A(4), A2 => n4, B1 => B(4), B2 => n3, ZN => 
                           n17);
   U25 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => Y(3));
   U26 : AOI22_X1 port map( A1 => C(3), A2 => n7, B1 => D(3), B2 => n8, ZN => 
                           n20);
   U27 : AOI22_X1 port map( A1 => A(3), A2 => n4, B1 => B(3), B2 => n3, ZN => 
                           n19);
   U28 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => Y(31));
   U29 : AOI22_X1 port map( A1 => C(31), A2 => n7, B1 => D(31), B2 => n8, ZN =>
                           n22);
   U30 : AOI22_X1 port map( A1 => A(31), A2 => n4, B1 => B(31), B2 => n3, ZN =>
                           n21);
   U31 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => Y(30));
   U32 : AOI22_X1 port map( A1 => C(30), A2 => n7, B1 => D(30), B2 => n8, ZN =>
                           n24);
   U33 : AOI22_X1 port map( A1 => A(30), A2 => n4, B1 => B(30), B2 => n3, ZN =>
                           n23);
   U34 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => Y(2));
   U35 : AOI22_X1 port map( A1 => C(2), A2 => n7, B1 => D(2), B2 => n8, ZN => 
                           n26);
   U36 : AOI22_X1 port map( A1 => A(2), A2 => n4, B1 => B(2), B2 => n3, ZN => 
                           n25);
   U37 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => Y(29));
   U38 : AOI22_X1 port map( A1 => C(29), A2 => n7, B1 => D(29), B2 => n8, ZN =>
                           n28);
   U39 : AOI22_X1 port map( A1 => A(29), A2 => n4, B1 => B(29), B2 => n3, ZN =>
                           n27);
   U40 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => Y(28));
   U41 : AOI22_X1 port map( A1 => C(28), A2 => n7, B1 => D(28), B2 => n8, ZN =>
                           n30);
   U42 : AOI22_X1 port map( A1 => A(28), A2 => n4, B1 => B(28), B2 => n3, ZN =>
                           n29);
   U43 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => Y(27));
   U44 : AOI22_X1 port map( A1 => C(27), A2 => n7, B1 => D(27), B2 => n8, ZN =>
                           n32);
   U45 : AOI22_X1 port map( A1 => A(27), A2 => n4, B1 => B(27), B2 => n3, ZN =>
                           n31);
   U46 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => Y(26));
   U47 : AOI22_X1 port map( A1 => C(26), A2 => n7, B1 => D(26), B2 => n8, ZN =>
                           n34);
   U48 : AOI22_X1 port map( A1 => A(26), A2 => n4, B1 => B(26), B2 => n3, ZN =>
                           n33);
   U49 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => Y(25));
   U50 : AOI22_X1 port map( A1 => C(25), A2 => n7, B1 => D(25), B2 => n8, ZN =>
                           n36);
   U51 : AOI22_X1 port map( A1 => A(25), A2 => n4, B1 => B(25), B2 => n3, ZN =>
                           n35);
   U52 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => Y(24));
   U53 : AOI22_X1 port map( A1 => C(24), A2 => n7, B1 => D(24), B2 => n8, ZN =>
                           n38);
   U54 : AOI22_X1 port map( A1 => A(24), A2 => n4, B1 => B(24), B2 => n3, ZN =>
                           n37);
   U55 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => Y(23));
   U56 : AOI22_X1 port map( A1 => C(23), A2 => n7, B1 => D(23), B2 => n8, ZN =>
                           n40);
   U57 : AOI22_X1 port map( A1 => A(23), A2 => n4, B1 => B(23), B2 => n3, ZN =>
                           n39);
   U58 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => Y(22));
   U59 : AOI22_X1 port map( A1 => C(22), A2 => n7, B1 => D(22), B2 => n8, ZN =>
                           n42);
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n4, B1 => B(22), B2 => n3, ZN =>
                           n41);
   U61 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => Y(21));
   U62 : AOI22_X1 port map( A1 => C(21), A2 => n7, B1 => D(21), B2 => n8, ZN =>
                           n44);
   U63 : AOI22_X1 port map( A1 => A(21), A2 => n4, B1 => B(21), B2 => n3, ZN =>
                           n43);
   U64 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => Y(20));
   U65 : AOI22_X1 port map( A1 => C(20), A2 => n7, B1 => D(20), B2 => n8, ZN =>
                           n46);
   U66 : AOI22_X1 port map( A1 => A(20), A2 => n4, B1 => B(20), B2 => n3, ZN =>
                           n45);
   U67 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => Y(1));
   U68 : AOI22_X1 port map( A1 => C(1), A2 => n7, B1 => D(1), B2 => n8, ZN => 
                           n48);
   U69 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n3, ZN => 
                           n47);
   U70 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => Y(19));
   U71 : AOI22_X1 port map( A1 => C(19), A2 => n7, B1 => D(19), B2 => n8, ZN =>
                           n50);
   U72 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n3, ZN =>
                           n49);
   U73 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => Y(18));
   U74 : AOI22_X1 port map( A1 => C(18), A2 => n7, B1 => D(18), B2 => n8, ZN =>
                           n52);
   U75 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n3, ZN =>
                           n51);
   U76 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => Y(17));
   U77 : AOI22_X1 port map( A1 => C(17), A2 => n7, B1 => D(17), B2 => n8, ZN =>
                           n54);
   U78 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n3, ZN =>
                           n53);
   U79 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => Y(16));
   U80 : AOI22_X1 port map( A1 => C(16), A2 => n7, B1 => D(16), B2 => n8, ZN =>
                           n56);
   U81 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n3, ZN =>
                           n55);
   U82 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => Y(15));
   U83 : AOI22_X1 port map( A1 => C(15), A2 => n7, B1 => D(15), B2 => n8, ZN =>
                           n58);
   U84 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n3, ZN =>
                           n57);
   U85 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => Y(14));
   U86 : AOI22_X1 port map( A1 => C(14), A2 => n7, B1 => D(14), B2 => n8, ZN =>
                           n60);
   U87 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n3, ZN =>
                           n59);
   U88 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => Y(13));
   U89 : AOI22_X1 port map( A1 => C(13), A2 => n7, B1 => D(13), B2 => n8, ZN =>
                           n62);
   U90 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n3, ZN =>
                           n61);
   U91 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => Y(12));
   U92 : AOI22_X1 port map( A1 => C(12), A2 => n7, B1 => D(12), B2 => n8, ZN =>
                           n64);
   U93 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n3, ZN =>
                           n63);
   U94 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => Y(11));
   U95 : AOI22_X1 port map( A1 => C(11), A2 => n7, B1 => D(11), B2 => n8, ZN =>
                           n66);
   U96 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n3, ZN =>
                           n65);
   U97 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => Y(10));
   U98 : AOI22_X1 port map( A1 => C(10), A2 => n7, B1 => D(10), B2 => n8, ZN =>
                           n68);
   U99 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n3, ZN =>
                           n67);
   U100 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => Y(0));
   U101 : AOI22_X1 port map( A1 => C(0), A2 => n7, B1 => D(0), B2 => n8, ZN => 
                           n70);
   U102 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n3, ZN => 
                           n69);
   U103 : INV_X1 port map( A => S(0), ZN => n71);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity REGADDR_N32_OPC6_REG5 is

   port( INSTR : in std_logic_vector (31 downto 0);  RS1, RS2, RD : out 
         std_logic_vector (4 downto 0));

end REGADDR_N32_OPC6_REG5;

architecture SYN_BEHAVIORAL of REGADDR_N32_OPC6_REG5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32 : std_logic;

begin
   
   U3 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => RS2(4));
   U4 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => RS2(3));
   U5 : NOR2_X1 port map( A1 => n1, A2 => n4, ZN => RS2(2));
   U6 : NOR2_X1 port map( A1 => n1, A2 => n5, ZN => RS2(1));
   U7 : NOR2_X1 port map( A1 => n1, A2 => n6, ZN => RS2(0));
   U8 : OAI211_X1 port map( C1 => n7, C2 => n8, A => n9, B => n10, ZN => n1);
   U9 : NOR2_X1 port map( A1 => INSTR(30), A2 => INSTR(28), ZN => n10);
   U10 : MUX2_X1 port map( A => n11, B => INSTR(31), S => n12, Z => n9);
   U11 : XNOR2_X1 port map( A => n13, B => n14, ZN => n12);
   U12 : INV_X1 port map( A => INSTR(31), ZN => n8);
   U13 : INV_X1 port map( A => n11, ZN => n7);
   U14 : AOI21_X1 port map( B1 => n14, B2 => INSTR(29), A => n15, ZN => n11);
   U15 : XNOR2_X1 port map( A => INSTR(26), B => n16, ZN => n14);
   U16 : AND2_X1 port map( A1 => INSTR(25), A2 => n17, ZN => RS1(4));
   U17 : AND2_X1 port map( A1 => INSTR(24), A2 => n17, ZN => RS1(3));
   U18 : AND2_X1 port map( A1 => INSTR(23), A2 => n17, ZN => RS1(2));
   U19 : AND2_X1 port map( A1 => INSTR(22), A2 => n17, ZN => RS1(1));
   U20 : AND2_X1 port map( A1 => INSTR(21), A2 => n17, ZN => RS1(0));
   U21 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n17);
   U22 : OAI221_X1 port map( B1 => n2, B2 => n20, C1 => n21, C2 => n22, A => 
                           n23, ZN => RD(4));
   U23 : INV_X1 port map( A => INSTR(15), ZN => n22);
   U24 : INV_X1 port map( A => INSTR(20), ZN => n2);
   U25 : OAI221_X1 port map( B1 => n3, B2 => n20, C1 => n21, C2 => n24, A => 
                           n23, ZN => RD(3));
   U26 : INV_X1 port map( A => INSTR(14), ZN => n24);
   U27 : INV_X1 port map( A => INSTR(19), ZN => n3);
   U28 : OAI221_X1 port map( B1 => n4, B2 => n20, C1 => n21, C2 => n25, A => 
                           n23, ZN => RD(2));
   U29 : INV_X1 port map( A => INSTR(13), ZN => n25);
   U30 : INV_X1 port map( A => INSTR(18), ZN => n4);
   U31 : OAI221_X1 port map( B1 => n5, B2 => n20, C1 => n21, C2 => n26, A => 
                           n23, ZN => RD(1));
   U32 : INV_X1 port map( A => INSTR(12), ZN => n26);
   U33 : INV_X1 port map( A => INSTR(17), ZN => n5);
   U34 : OAI221_X1 port map( B1 => n6, B2 => n20, C1 => n21, C2 => n27, A => 
                           n23, ZN => RD(0));
   U35 : NAND2_X1 port map( A1 => n18, A2 => INSTR(26), ZN => n23);
   U36 : INV_X1 port map( A => n28, ZN => n18);
   U37 : INV_X1 port map( A => INSTR(11), ZN => n27);
   U38 : NAND3_X1 port map( A1 => n21, A2 => n28, A3 => n29, ZN => n20);
   U39 : NAND3_X1 port map( A1 => n15, A2 => INSTR(31), A3 => n30, ZN => n29);
   U40 : NOR3_X1 port map( A1 => n13, A2 => INSTR(30), A3 => INSTR(28), ZN => 
                           n30);
   U41 : INV_X1 port map( A => INSTR(29), ZN => n13);
   U42 : NOR2_X1 port map( A1 => n31, A2 => n16, ZN => n15);
   U43 : NAND2_X1 port map( A1 => n32, A2 => INSTR(27), ZN => n28);
   U44 : NAND4_X1 port map( A1 => n32, A2 => n31, A3 => n16, A4 => n19, ZN => 
                           n21);
   U45 : INV_X1 port map( A => INSTR(30), ZN => n19);
   U46 : INV_X1 port map( A => INSTR(27), ZN => n16);
   U47 : INV_X1 port map( A => INSTR(26), ZN => n31);
   U48 : NOR3_X1 port map( A1 => INSTR(29), A2 => INSTR(31), A3 => INSTR(28), 
                           ZN => n32);
   U49 : INV_X1 port map( A => INSTR(16), ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SIGNEX_N32_OPC6_REG5 is

   port( INSTR : in std_logic_vector (31 downto 0);  IMM : out std_logic_vector
         (31 downto 0));

end SIGNEX_N32_OPC6_REG5;

architecture SYN_BEHAVIORAL of SIGNEX_N32_OPC6_REG5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50 : std_logic;

begin
   
   U2 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           IMM(31));
   U3 : NOR2_X1 port map( A1 => n5, A2 => n6, ZN => IMM(9));
   U4 : NOR2_X1 port map( A1 => n5, A2 => n7, ZN => IMM(8));
   U5 : NOR2_X1 port map( A1 => n5, A2 => n8, ZN => IMM(7));
   U6 : NOR2_X1 port map( A1 => n5, A2 => n9, ZN => IMM(6));
   U7 : NOR2_X1 port map( A1 => n5, A2 => n10, ZN => IMM(5));
   U8 : NOR2_X1 port map( A1 => n5, A2 => n11, ZN => IMM(4));
   U9 : NOR2_X1 port map( A1 => n5, A2 => n12, ZN => IMM(3));
   U10 : OAI21_X1 port map( B1 => n13, B2 => n14, A => n15, ZN => IMM(30));
   U11 : NOR2_X1 port map( A1 => n5, A2 => n16, ZN => IMM(2));
   U12 : OAI21_X1 port map( B1 => n13, B2 => n17, A => n15, ZN => IMM(29));
   U13 : OAI21_X1 port map( B1 => n13, B2 => n18, A => n15, ZN => IMM(28));
   U14 : OAI21_X1 port map( B1 => n13, B2 => n19, A => n15, ZN => IMM(27));
   U15 : OAI21_X1 port map( B1 => n13, B2 => n20, A => n15, ZN => IMM(26));
   U16 : OAI21_X1 port map( B1 => n6, B2 => n13, A => n15, ZN => IMM(25));
   U17 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => n15);
   U18 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n23, B2 => n4, ZN => n22)
                           ;
   U19 : INV_X1 port map( A => n13, ZN => n23);
   U20 : INV_X1 port map( A => INSTR(25), ZN => n2);
   U21 : INV_X1 port map( A => INSTR(9), ZN => n6);
   U22 : OAI21_X1 port map( B1 => n7, B2 => n13, A => n24, ZN => IMM(24));
   U23 : AOI21_X1 port map( B1 => INSTR(24), B2 => n25, A => n26, ZN => n24);
   U24 : INV_X1 port map( A => INSTR(8), ZN => n7);
   U25 : OAI21_X1 port map( B1 => n8, B2 => n13, A => n27, ZN => IMM(23));
   U26 : AOI21_X1 port map( B1 => INSTR(23), B2 => n25, A => n26, ZN => n27);
   U27 : INV_X1 port map( A => INSTR(7), ZN => n8);
   U28 : OAI21_X1 port map( B1 => n9, B2 => n13, A => n28, ZN => IMM(22));
   U29 : AOI21_X1 port map( B1 => INSTR(22), B2 => n25, A => n26, ZN => n28);
   U30 : INV_X1 port map( A => INSTR(6), ZN => n9);
   U31 : OAI21_X1 port map( B1 => n10, B2 => n13, A => n29, ZN => IMM(21));
   U32 : AOI21_X1 port map( B1 => INSTR(21), B2 => n25, A => n26, ZN => n29);
   U33 : INV_X1 port map( A => INSTR(5), ZN => n10);
   U34 : OAI21_X1 port map( B1 => n11, B2 => n13, A => n30, ZN => IMM(20));
   U35 : AOI21_X1 port map( B1 => INSTR(20), B2 => n25, A => n26, ZN => n30);
   U36 : INV_X1 port map( A => INSTR(4), ZN => n11);
   U37 : NOR2_X1 port map( A1 => n5, A2 => n31, ZN => IMM(1));
   U38 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n32, ZN => IMM(19));
   U39 : AOI21_X1 port map( B1 => INSTR(19), B2 => n25, A => n26, ZN => n32);
   U40 : INV_X1 port map( A => INSTR(3), ZN => n12);
   U41 : OAI21_X1 port map( B1 => n13, B2 => n16, A => n33, ZN => IMM(18));
   U42 : AOI21_X1 port map( B1 => INSTR(18), B2 => n25, A => n26, ZN => n33);
   U43 : INV_X1 port map( A => INSTR(2), ZN => n16);
   U44 : OAI21_X1 port map( B1 => n13, B2 => n31, A => n34, ZN => IMM(17));
   U45 : AOI21_X1 port map( B1 => INSTR(17), B2 => n25, A => n26, ZN => n34);
   U46 : INV_X1 port map( A => INSTR(1), ZN => n31);
   U47 : OAI21_X1 port map( B1 => n13, B2 => n35, A => n36, ZN => IMM(16));
   U48 : AOI21_X1 port map( B1 => INSTR(16), B2 => n25, A => n26, ZN => n36);
   U49 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => n26);
   U50 : NAND3_X1 port map( A1 => INSTR(15), A2 => n1, A3 => n37, ZN => n4);
   U51 : MUX2_X1 port map( A => n38, B => n39, S => INSTR(31), Z => n37);
   U52 : NAND4_X1 port map( A1 => INSTR(30), A2 => INSTR(29), A3 => n40, A4 => 
                           n41, ZN => n39);
   U53 : INV_X1 port map( A => n42, ZN => n41);
   U54 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => n40);
   U55 : OAI211_X1 port map( C1 => n42, C2 => n45, A => n46, B => INSTR(26), ZN
                           => n38);
   U56 : MUX2_X1 port map( A => n44, B => INSTR(30), S => n47, Z => n46);
   U57 : INV_X1 port map( A => INSTR(30), ZN => n45);
   U58 : INV_X1 port map( A => n25, ZN => n1);
   U59 : NOR2_X1 port map( A1 => n43, A2 => n48, ZN => n25);
   U60 : NOR2_X1 port map( A1 => n49, A2 => n5, ZN => IMM(15));
   U61 : INV_X1 port map( A => INSTR(15), ZN => n49);
   U62 : NOR2_X1 port map( A1 => n5, A2 => n14, ZN => IMM(14));
   U63 : INV_X1 port map( A => INSTR(14), ZN => n14);
   U64 : NOR2_X1 port map( A1 => n5, A2 => n17, ZN => IMM(13));
   U65 : INV_X1 port map( A => INSTR(13), ZN => n17);
   U66 : NOR2_X1 port map( A1 => n5, A2 => n18, ZN => IMM(12));
   U67 : INV_X1 port map( A => INSTR(12), ZN => n18);
   U68 : NOR2_X1 port map( A1 => n5, A2 => n19, ZN => IMM(11));
   U69 : INV_X1 port map( A => INSTR(11), ZN => n19);
   U70 : NOR2_X1 port map( A1 => n5, A2 => n20, ZN => IMM(10));
   U71 : INV_X1 port map( A => INSTR(10), ZN => n20);
   U72 : NOR2_X1 port map( A1 => n5, A2 => n35, ZN => IMM(0));
   U73 : INV_X1 port map( A => INSTR(0), ZN => n35);
   U74 : NAND2_X1 port map( A1 => n13, A2 => n21, ZN => n5);
   U75 : INV_X1 port map( A => n3, ZN => n21);
   U76 : NOR3_X1 port map( A1 => INSTR(26), A2 => INSTR(27), A3 => n48, ZN => 
                           n3);
   U77 : OR4_X1 port map( A1 => INSTR(28), A2 => INSTR(29), A3 => INSTR(30), A4
                           => INSTR(31), ZN => n48);
   U78 : NAND3_X1 port map( A1 => n42, A2 => INSTR(26), A3 => n50, ZN => n13);
   U79 : NOR3_X1 port map( A1 => n47, A2 => INSTR(31), A3 => INSTR(30), ZN => 
                           n50);
   U80 : INV_X1 port map( A => INSTR(29), ZN => n47);
   U81 : NOR2_X1 port map( A1 => n44, A2 => n43, ZN => n42);
   U82 : INV_X1 port map( A => INSTR(27), ZN => n43);
   U83 : INV_X1 port map( A => INSTR(28), ZN => n44);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RF_N32_NA5 is

   port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
         ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_N32_NA5;

architecture SYN_BEHAVIORAL of RF_N32_NA5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REG_0_31_port, REG_0_30_port, REG_0_29_port, REG_0_28_port, 
      REG_0_27_port, REG_0_26_port, REG_0_25_port, REG_0_24_port, REG_0_23_port
      , REG_0_22_port, REG_0_21_port, REG_0_20_port, REG_0_19_port, 
      REG_0_18_port, REG_0_17_port, REG_0_16_port, REG_0_15_port, REG_0_14_port
      , REG_0_13_port, REG_0_12_port, REG_0_11_port, REG_0_10_port, 
      REG_0_9_port, REG_0_8_port, REG_0_7_port, REG_0_6_port, REG_0_5_port, 
      REG_0_4_port, REG_0_3_port, REG_0_2_port, REG_0_1_port, REG_0_0_port, 
      REG_1_31_port, REG_1_30_port, REG_1_29_port, REG_1_28_port, REG_1_27_port
      , REG_1_26_port, REG_1_25_port, REG_1_24_port, REG_1_23_port, 
      REG_1_22_port, REG_1_21_port, REG_1_20_port, REG_1_19_port, REG_1_18_port
      , REG_1_17_port, REG_1_16_port, REG_1_15_port, REG_1_14_port, 
      REG_1_13_port, REG_1_12_port, REG_1_11_port, REG_1_10_port, REG_1_9_port,
      REG_1_8_port, REG_1_7_port, REG_1_6_port, REG_1_5_port, REG_1_4_port, 
      REG_1_3_port, REG_1_2_port, REG_1_1_port, REG_1_0_port, REG_2_31_port, 
      REG_2_30_port, REG_2_29_port, REG_2_28_port, REG_2_27_port, REG_2_26_port
      , REG_2_25_port, REG_2_24_port, REG_2_23_port, REG_2_22_port, 
      REG_2_21_port, REG_2_20_port, REG_2_19_port, REG_2_18_port, REG_2_17_port
      , REG_2_16_port, REG_2_15_port, REG_2_14_port, REG_2_13_port, 
      REG_2_12_port, REG_2_11_port, REG_2_10_port, REG_2_9_port, REG_2_8_port, 
      REG_2_7_port, REG_2_6_port, REG_2_5_port, REG_2_4_port, REG_2_3_port, 
      REG_2_2_port, REG_2_1_port, REG_2_0_port, REG_3_31_port, REG_3_30_port, 
      REG_3_29_port, REG_3_28_port, REG_3_27_port, REG_3_26_port, REG_3_25_port
      , REG_3_24_port, REG_3_23_port, REG_3_22_port, REG_3_21_port, 
      REG_3_20_port, REG_3_19_port, REG_3_18_port, REG_3_17_port, REG_3_16_port
      , REG_3_15_port, REG_3_14_port, REG_3_13_port, REG_3_12_port, 
      REG_3_11_port, REG_3_10_port, REG_3_9_port, REG_3_8_port, REG_3_7_port, 
      REG_3_6_port, REG_3_5_port, REG_3_4_port, REG_3_3_port, REG_3_2_port, 
      REG_3_1_port, REG_3_0_port, REG_4_31_port, REG_4_30_port, REG_4_29_port, 
      REG_4_28_port, REG_4_27_port, REG_4_26_port, REG_4_25_port, REG_4_24_port
      , REG_4_23_port, REG_4_22_port, REG_4_21_port, REG_4_20_port, 
      REG_4_19_port, REG_4_18_port, REG_4_17_port, REG_4_16_port, REG_4_15_port
      , REG_4_14_port, REG_4_13_port, REG_4_12_port, REG_4_11_port, 
      REG_4_10_port, REG_4_9_port, REG_4_8_port, REG_4_7_port, REG_4_6_port, 
      REG_4_5_port, REG_4_4_port, REG_4_3_port, REG_4_2_port, REG_4_1_port, 
      REG_4_0_port, REG_5_31_port, REG_5_30_port, REG_5_29_port, REG_5_28_port,
      REG_5_27_port, REG_5_26_port, REG_5_25_port, REG_5_24_port, REG_5_23_port
      , REG_5_22_port, REG_5_21_port, REG_5_20_port, REG_5_19_port, 
      REG_5_18_port, REG_5_17_port, REG_5_16_port, REG_5_15_port, REG_5_14_port
      , REG_5_13_port, REG_5_12_port, REG_5_11_port, REG_5_10_port, 
      REG_5_9_port, REG_5_8_port, REG_5_7_port, REG_5_6_port, REG_5_5_port, 
      REG_5_4_port, REG_5_3_port, REG_5_2_port, REG_5_1_port, REG_5_0_port, 
      REG_6_31_port, REG_6_30_port, REG_6_29_port, REG_6_28_port, REG_6_27_port
      , REG_6_26_port, REG_6_25_port, REG_6_24_port, REG_6_23_port, 
      REG_6_22_port, REG_6_21_port, REG_6_20_port, REG_6_19_port, REG_6_18_port
      , REG_6_17_port, REG_6_16_port, REG_6_15_port, REG_6_14_port, 
      REG_6_13_port, REG_6_12_port, REG_6_11_port, REG_6_10_port, REG_6_9_port,
      REG_6_8_port, REG_6_7_port, REG_6_6_port, REG_6_5_port, REG_6_4_port, 
      REG_6_3_port, REG_6_2_port, REG_6_1_port, REG_6_0_port, REG_7_31_port, 
      REG_7_30_port, REG_7_29_port, REG_7_28_port, REG_7_27_port, REG_7_26_port
      , REG_7_25_port, REG_7_24_port, REG_7_23_port, REG_7_22_port, 
      REG_7_21_port, REG_7_20_port, REG_7_19_port, REG_7_18_port, REG_7_17_port
      , REG_7_16_port, REG_7_15_port, REG_7_14_port, REG_7_13_port, 
      REG_7_12_port, REG_7_11_port, REG_7_10_port, REG_7_9_port, REG_7_8_port, 
      REG_7_7_port, REG_7_6_port, REG_7_5_port, REG_7_4_port, REG_7_3_port, 
      REG_7_2_port, REG_7_1_port, REG_7_0_port, REG_8_31_port, REG_8_30_port, 
      REG_8_29_port, REG_8_28_port, REG_8_27_port, REG_8_26_port, REG_8_25_port
      , REG_8_24_port, REG_8_23_port, REG_8_22_port, REG_8_21_port, 
      REG_8_20_port, REG_8_19_port, REG_8_18_port, REG_8_17_port, REG_8_16_port
      , REG_8_15_port, REG_8_14_port, REG_8_13_port, REG_8_12_port, 
      REG_8_11_port, REG_8_10_port, REG_8_9_port, REG_8_8_port, REG_8_7_port, 
      REG_8_6_port, REG_8_5_port, REG_8_4_port, REG_8_3_port, REG_8_2_port, 
      REG_8_1_port, REG_8_0_port, REG_9_31_port, REG_9_30_port, REG_9_29_port, 
      REG_9_28_port, REG_9_27_port, REG_9_26_port, REG_9_25_port, REG_9_24_port
      , REG_9_23_port, REG_9_22_port, REG_9_21_port, REG_9_20_port, 
      REG_9_19_port, REG_9_18_port, REG_9_17_port, REG_9_16_port, REG_9_15_port
      , REG_9_14_port, REG_9_13_port, REG_9_12_port, REG_9_11_port, 
      REG_9_10_port, REG_9_9_port, REG_9_8_port, REG_9_7_port, REG_9_6_port, 
      REG_9_5_port, REG_9_4_port, REG_9_3_port, REG_9_2_port, REG_9_1_port, 
      REG_9_0_port, REG_10_31_port, REG_10_30_port, REG_10_29_port, 
      REG_10_28_port, REG_10_27_port, REG_10_26_port, REG_10_25_port, 
      REG_10_24_port, REG_10_23_port, REG_10_22_port, REG_10_21_port, 
      REG_10_20_port, REG_10_19_port, REG_10_18_port, REG_10_17_port, 
      REG_10_16_port, REG_10_15_port, REG_10_14_port, REG_10_13_port, 
      REG_10_12_port, REG_10_11_port, REG_10_10_port, REG_10_9_port, 
      REG_10_8_port, REG_10_7_port, REG_10_6_port, REG_10_5_port, REG_10_4_port
      , REG_10_3_port, REG_10_2_port, REG_10_1_port, REG_10_0_port, 
      REG_11_31_port, REG_11_30_port, REG_11_29_port, REG_11_28_port, 
      REG_11_27_port, REG_11_26_port, REG_11_25_port, REG_11_24_port, 
      REG_11_23_port, REG_11_22_port, REG_11_21_port, REG_11_20_port, 
      REG_11_19_port, REG_11_18_port, REG_11_17_port, REG_11_16_port, 
      REG_11_15_port, REG_11_14_port, REG_11_13_port, REG_11_12_port, 
      REG_11_11_port, REG_11_10_port, REG_11_9_port, REG_11_8_port, 
      REG_11_7_port, REG_11_6_port, REG_11_5_port, REG_11_4_port, REG_11_3_port
      , REG_11_2_port, REG_11_1_port, REG_11_0_port, REG_12_31_port, 
      REG_12_30_port, REG_12_29_port, REG_12_28_port, REG_12_27_port, 
      REG_12_26_port, REG_12_25_port, REG_12_24_port, REG_12_23_port, 
      REG_12_22_port, REG_12_21_port, REG_12_20_port, REG_12_19_port, 
      REG_12_18_port, REG_12_17_port, REG_12_16_port, REG_12_15_port, 
      REG_12_14_port, REG_12_13_port, REG_12_12_port, REG_12_11_port, 
      REG_12_10_port, REG_12_9_port, REG_12_8_port, REG_12_7_port, 
      REG_12_6_port, REG_12_5_port, REG_12_4_port, REG_12_3_port, REG_12_2_port
      , REG_12_1_port, REG_12_0_port, REG_13_31_port, REG_13_30_port, 
      REG_13_29_port, REG_13_28_port, REG_13_27_port, REG_13_26_port, 
      REG_13_25_port, REG_13_24_port, REG_13_23_port, REG_13_22_port, 
      REG_13_21_port, REG_13_20_port, REG_13_19_port, REG_13_18_port, 
      REG_13_17_port, REG_13_16_port, REG_13_15_port, REG_13_14_port, 
      REG_13_13_port, REG_13_12_port, REG_13_11_port, REG_13_10_port, 
      REG_13_9_port, REG_13_8_port, REG_13_7_port, REG_13_6_port, REG_13_5_port
      , REG_13_4_port, REG_13_3_port, REG_13_2_port, REG_13_1_port, 
      REG_13_0_port, REG_14_31_port, REG_14_30_port, REG_14_29_port, 
      REG_14_28_port, REG_14_27_port, REG_14_26_port, REG_14_25_port, 
      REG_14_24_port, REG_14_23_port, REG_14_22_port, REG_14_21_port, 
      REG_14_20_port, REG_14_19_port, REG_14_18_port, REG_14_17_port, 
      REG_14_16_port, REG_14_15_port, REG_14_14_port, REG_14_13_port, 
      REG_14_12_port, REG_14_11_port, REG_14_10_port, REG_14_9_port, 
      REG_14_8_port, REG_14_7_port, REG_14_6_port, REG_14_5_port, REG_14_4_port
      , REG_14_3_port, REG_14_2_port, REG_14_1_port, REG_14_0_port, 
      REG_15_31_port, REG_15_30_port, REG_15_29_port, REG_15_28_port, 
      REG_15_27_port, REG_15_26_port, REG_15_25_port, REG_15_24_port, 
      REG_15_23_port, REG_15_22_port, REG_15_21_port, REG_15_20_port, 
      REG_15_19_port, REG_15_18_port, REG_15_17_port, REG_15_16_port, 
      REG_15_15_port, REG_15_14_port, REG_15_13_port, REG_15_12_port, 
      REG_15_11_port, REG_15_10_port, REG_15_9_port, REG_15_8_port, 
      REG_15_7_port, REG_15_6_port, REG_15_5_port, REG_15_4_port, REG_15_3_port
      , REG_15_2_port, REG_15_1_port, REG_15_0_port, REG_16_31_port, 
      REG_16_30_port, REG_16_29_port, REG_16_28_port, REG_16_27_port, 
      REG_16_26_port, REG_16_25_port, REG_16_24_port, REG_16_23_port, 
      REG_16_22_port, REG_16_21_port, REG_16_20_port, REG_16_19_port, 
      REG_16_18_port, REG_16_17_port, REG_16_16_port, REG_16_15_port, 
      REG_16_14_port, REG_16_13_port, REG_16_12_port, REG_16_11_port, 
      REG_16_10_port, REG_16_9_port, REG_16_8_port, REG_16_7_port, 
      REG_16_6_port, REG_16_5_port, REG_16_4_port, REG_16_3_port, REG_16_2_port
      , REG_16_1_port, REG_16_0_port, REG_17_31_port, REG_17_30_port, 
      REG_17_29_port, REG_17_28_port, REG_17_27_port, REG_17_26_port, 
      REG_17_25_port, REG_17_24_port, REG_17_23_port, REG_17_22_port, 
      REG_17_21_port, REG_17_20_port, REG_17_19_port, REG_17_18_port, 
      REG_17_17_port, REG_17_16_port, REG_17_15_port, REG_17_14_port, 
      REG_17_13_port, REG_17_12_port, REG_17_11_port, REG_17_10_port, 
      REG_17_9_port, REG_17_8_port, REG_17_7_port, REG_17_6_port, REG_17_5_port
      , REG_17_4_port, REG_17_3_port, REG_17_2_port, REG_17_1_port, 
      REG_17_0_port, REG_18_31_port, REG_18_30_port, REG_18_29_port, 
      REG_18_28_port, REG_18_27_port, REG_18_26_port, REG_18_25_port, 
      REG_18_24_port, REG_18_23_port, REG_18_22_port, REG_18_21_port, 
      REG_18_20_port, REG_18_19_port, REG_18_18_port, REG_18_17_port, 
      REG_18_16_port, REG_18_15_port, REG_18_14_port, REG_18_13_port, 
      REG_18_12_port, REG_18_11_port, REG_18_10_port, REG_18_9_port, 
      REG_18_8_port, REG_18_7_port, REG_18_6_port, REG_18_5_port, REG_18_4_port
      , REG_18_3_port, REG_18_2_port, REG_18_1_port, REG_18_0_port, 
      REG_19_31_port, REG_19_30_port, REG_19_29_port, REG_19_28_port, 
      REG_19_27_port, REG_19_26_port, REG_19_25_port, REG_19_24_port, 
      REG_19_23_port, REG_19_22_port, REG_19_21_port, REG_19_20_port, 
      REG_19_19_port, REG_19_18_port, REG_19_17_port, REG_19_16_port, 
      REG_19_15_port, REG_19_14_port, REG_19_13_port, REG_19_12_port, 
      REG_19_11_port, REG_19_10_port, REG_19_9_port, REG_19_8_port, 
      REG_19_7_port, REG_19_6_port, REG_19_5_port, REG_19_4_port, REG_19_3_port
      , REG_19_2_port, REG_19_1_port, REG_19_0_port, REG_20_31_port, 
      REG_20_30_port, REG_20_29_port, REG_20_28_port, REG_20_27_port, 
      REG_20_26_port, REG_20_25_port, REG_20_24_port, REG_20_23_port, 
      REG_20_22_port, REG_20_21_port, REG_20_20_port, REG_20_19_port, 
      REG_20_18_port, REG_20_17_port, REG_20_16_port, REG_20_15_port, 
      REG_20_14_port, REG_20_13_port, REG_20_12_port, REG_20_11_port, 
      REG_20_10_port, REG_20_9_port, REG_20_8_port, REG_20_7_port, 
      REG_20_6_port, REG_20_5_port, REG_20_4_port, REG_20_3_port, REG_20_2_port
      , REG_20_1_port, REG_20_0_port, REG_21_31_port, REG_21_30_port, 
      REG_21_29_port, REG_21_28_port, REG_21_27_port, REG_21_26_port, 
      REG_21_25_port, REG_21_24_port, REG_21_23_port, REG_21_22_port, 
      REG_21_21_port, REG_21_20_port, REG_21_19_port, REG_21_18_port, 
      REG_21_17_port, REG_21_16_port, REG_21_15_port, REG_21_14_port, 
      REG_21_13_port, REG_21_12_port, REG_21_11_port, REG_21_10_port, 
      REG_21_9_port, REG_21_8_port, REG_21_7_port, REG_21_6_port, REG_21_5_port
      , REG_21_4_port, REG_21_3_port, REG_21_2_port, REG_21_1_port, 
      REG_21_0_port, REG_22_31_port, REG_22_30_port, REG_22_29_port, 
      REG_22_28_port, REG_22_27_port, REG_22_26_port, REG_22_25_port, 
      REG_22_24_port, REG_22_23_port, REG_22_22_port, REG_22_21_port, 
      REG_22_20_port, REG_22_19_port, REG_22_18_port, REG_22_17_port, 
      REG_22_16_port, REG_22_15_port, REG_22_14_port, REG_22_13_port, 
      REG_22_12_port, REG_22_11_port, REG_22_10_port, REG_22_9_port, 
      REG_22_8_port, REG_22_7_port, REG_22_6_port, REG_22_5_port, REG_22_4_port
      , REG_22_3_port, REG_22_2_port, REG_22_1_port, REG_22_0_port, 
      REG_23_31_port, REG_23_30_port, REG_23_29_port, REG_23_28_port, 
      REG_23_27_port, REG_23_26_port, REG_23_25_port, REG_23_24_port, 
      REG_23_23_port, REG_23_22_port, REG_23_21_port, REG_23_20_port, 
      REG_23_19_port, REG_23_18_port, REG_23_17_port, REG_23_16_port, 
      REG_23_15_port, REG_23_14_port, REG_23_13_port, REG_23_12_port, 
      REG_23_11_port, REG_23_10_port, REG_23_9_port, REG_23_8_port, 
      REG_23_7_port, REG_23_6_port, REG_23_5_port, REG_23_4_port, REG_23_3_port
      , REG_23_2_port, REG_23_1_port, REG_23_0_port, REG_24_31_port, 
      REG_24_30_port, REG_24_29_port, REG_24_28_port, REG_24_27_port, 
      REG_24_26_port, REG_24_25_port, REG_24_24_port, REG_24_23_port, 
      REG_24_22_port, REG_24_21_port, REG_24_20_port, REG_24_19_port, 
      REG_24_18_port, REG_24_17_port, REG_24_16_port, REG_24_15_port, 
      REG_24_14_port, REG_24_13_port, REG_24_12_port, REG_24_11_port, 
      REG_24_10_port, REG_24_9_port, REG_24_8_port, REG_24_7_port, 
      REG_24_6_port, REG_24_5_port, REG_24_4_port, REG_24_3_port, REG_24_2_port
      , REG_24_1_port, REG_24_0_port, REG_25_31_port, REG_25_30_port, 
      REG_25_29_port, REG_25_28_port, REG_25_27_port, REG_25_26_port, 
      REG_25_25_port, REG_25_24_port, REG_25_23_port, REG_25_22_port, 
      REG_25_21_port, REG_25_20_port, REG_25_19_port, REG_25_18_port, 
      REG_25_17_port, REG_25_16_port, REG_25_15_port, REG_25_14_port, 
      REG_25_13_port, REG_25_12_port, REG_25_11_port, REG_25_10_port, 
      REG_25_9_port, REG_25_8_port, REG_25_7_port, REG_25_6_port, REG_25_5_port
      , REG_25_4_port, REG_25_3_port, REG_25_2_port, REG_25_1_port, 
      REG_25_0_port, REG_26_31_port, REG_26_30_port, REG_26_29_port, 
      REG_26_28_port, REG_26_27_port, REG_26_26_port, REG_26_25_port, 
      REG_26_24_port, REG_26_23_port, REG_26_22_port, REG_26_21_port, 
      REG_26_20_port, REG_26_19_port, REG_26_18_port, REG_26_17_port, 
      REG_26_16_port, REG_26_15_port, REG_26_14_port, REG_26_13_port, 
      REG_26_12_port, REG_26_11_port, REG_26_10_port, REG_26_9_port, 
      REG_26_8_port, REG_26_7_port, REG_26_6_port, REG_26_5_port, REG_26_4_port
      , REG_26_3_port, REG_26_2_port, REG_26_1_port, REG_26_0_port, 
      REG_27_31_port, REG_27_30_port, REG_27_29_port, REG_27_28_port, 
      REG_27_27_port, REG_27_26_port, REG_27_25_port, REG_27_24_port, 
      REG_27_23_port, REG_27_22_port, REG_27_21_port, REG_27_20_port, 
      REG_27_19_port, REG_27_18_port, REG_27_17_port, REG_27_16_port, 
      REG_27_15_port, REG_27_14_port, REG_27_13_port, REG_27_12_port, 
      REG_27_11_port, REG_27_10_port, REG_27_9_port, REG_27_8_port, 
      REG_27_7_port, REG_27_6_port, REG_27_5_port, REG_27_4_port, REG_27_3_port
      , REG_27_2_port, REG_27_1_port, REG_27_0_port, REG_28_31_port, 
      REG_28_30_port, REG_28_29_port, REG_28_28_port, REG_28_27_port, 
      REG_28_26_port, REG_28_25_port, REG_28_24_port, REG_28_23_port, 
      REG_28_22_port, REG_28_21_port, REG_28_20_port, REG_28_19_port, 
      REG_28_18_port, REG_28_17_port, REG_28_16_port, REG_28_15_port, 
      REG_28_14_port, REG_28_13_port, REG_28_12_port, REG_28_11_port, 
      REG_28_10_port, REG_28_9_port, REG_28_8_port, REG_28_7_port, 
      REG_28_6_port, REG_28_5_port, REG_28_4_port, REG_28_3_port, REG_28_2_port
      , REG_28_1_port, REG_28_0_port, REG_29_31_port, REG_29_30_port, 
      REG_29_29_port, REG_29_28_port, REG_29_27_port, REG_29_26_port, 
      REG_29_25_port, REG_29_24_port, REG_29_23_port, REG_29_22_port, 
      REG_29_21_port, REG_29_20_port, REG_29_19_port, REG_29_18_port, 
      REG_29_17_port, REG_29_16_port, REG_29_15_port, REG_29_14_port, 
      REG_29_13_port, REG_29_12_port, REG_29_11_port, REG_29_10_port, 
      REG_29_9_port, REG_29_8_port, REG_29_7_port, REG_29_6_port, REG_29_5_port
      , REG_29_4_port, REG_29_3_port, REG_29_2_port, REG_29_1_port, 
      REG_29_0_port, REG_30_31_port, REG_30_30_port, REG_30_29_port, 
      REG_30_28_port, REG_30_27_port, REG_30_26_port, REG_30_25_port, 
      REG_30_24_port, REG_30_23_port, REG_30_22_port, REG_30_21_port, 
      REG_30_20_port, REG_30_19_port, REG_30_18_port, REG_30_17_port, 
      REG_30_16_port, REG_30_15_port, REG_30_14_port, REG_30_13_port, 
      REG_30_12_port, REG_30_11_port, REG_30_10_port, REG_30_9_port, 
      REG_30_8_port, REG_30_7_port, REG_30_6_port, REG_30_5_port, REG_30_4_port
      , REG_30_3_port, REG_30_2_port, REG_30_1_port, REG_30_0_port, 
      REG_31_31_port, REG_31_30_port, REG_31_29_port, REG_31_28_port, 
      REG_31_27_port, REG_31_26_port, REG_31_25_port, REG_31_24_port, 
      REG_31_23_port, REG_31_22_port, REG_31_21_port, REG_31_20_port, 
      REG_31_19_port, REG_31_18_port, REG_31_17_port, REG_31_16_port, 
      REG_31_15_port, REG_31_14_port, REG_31_13_port, REG_31_12_port, 
      REG_31_11_port, REG_31_10_port, REG_31_9_port, REG_31_8_port, 
      REG_31_7_port, REG_31_6_port, REG_31_5_port, REG_31_4_port, REG_31_3_port
      , REG_31_2_port, REG_31_1_port, REG_31_0_port, N155, N188, N189, N190, 
      N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, 
      N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, 
      N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, 
      N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, 
      N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, 
      N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, 
      N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, 
      N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, 
      N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, 
      N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, 
      N312, N313, N314, N315, N316, N317, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109
      , n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155_port, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188_port, n189_port, n190_port
      , n191_port, n192_port, n193_port, n194_port, n195_port, n196_port, 
      n197_port, n198_port, n199_port, n200_port, n201_port, n202_port, 
      n203_port, n204_port, n205_port, n206_port, n207_port, n208_port, 
      n209_port, n210_port, n211_port, n212_port, n213_port, n214_port, 
      n215_port, n216_port, n217_port, n218_port, n219_port, n220_port, 
      n221_port, n222_port, n223_port, n224_port, n225_port, n226_port, 
      n227_port, n228_port, n229_port, n230_port, n231_port, n232_port, 
      n233_port, n234_port, n235_port, n236_port, n237_port, n238_port, 
      n239_port, n240_port, n241_port, n242_port, n243_port, n244_port, 
      n245_port, n246_port, n247_port, n248_port, n249_port, n250_port, n251, 
      n252_port, n253_port, n254_port, n255_port, n256_port, n257_port, 
      n258_port, n259_port, n260_port, n261_port, n262_port, n263_port, 
      n264_port, n265_port, n266_port, n267_port, n268_port, n269_port, 
      n270_port, n271_port, n272_port, n273_port, n274_port, n275_port, 
      n276_port, n277_port, n278_port, n279_port, n280_port, n281_port, 
      n282_port, n283_port, n284_port, n285_port, n286_port, n287_port, 
      n288_port, n289_port, n290_port, n291_port, n292_port, n293_port, 
      n294_port, n295_port, n296_port, n297_port, n298_port, n299_port, 
      n300_port, n301_port, n302_port, n303_port, n304_port, n305_port, 
      n306_port, n307_port, n308_port, n309_port, n310_port, n311_port, 
      n312_port, n313_port, n314_port, n315_port, n316_port, n317_port, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832 : 
      std_logic;

begin
   
   REG_reg_0_31_inst : DLH_X1 port map( G => N218, D => N250, Q => 
                           REG_0_31_port);
   REG_reg_0_30_inst : DLH_X1 port map( G => N218, D => N249, Q => 
                           REG_0_30_port);
   REG_reg_0_29_inst : DLH_X1 port map( G => N218, D => N248, Q => 
                           REG_0_29_port);
   REG_reg_0_28_inst : DLH_X1 port map( G => N218, D => N247, Q => 
                           REG_0_28_port);
   REG_reg_0_27_inst : DLH_X1 port map( G => N218, D => N246, Q => 
                           REG_0_27_port);
   REG_reg_0_26_inst : DLH_X1 port map( G => N218, D => N245, Q => 
                           REG_0_26_port);
   REG_reg_0_25_inst : DLH_X1 port map( G => N218, D => N244, Q => 
                           REG_0_25_port);
   REG_reg_0_24_inst : DLH_X1 port map( G => N218, D => N243, Q => 
                           REG_0_24_port);
   REG_reg_0_23_inst : DLH_X1 port map( G => N218, D => N242, Q => 
                           REG_0_23_port);
   REG_reg_0_22_inst : DLH_X1 port map( G => N218, D => N241, Q => 
                           REG_0_22_port);
   REG_reg_0_21_inst : DLH_X1 port map( G => N218, D => N240, Q => 
                           REG_0_21_port);
   REG_reg_0_20_inst : DLH_X1 port map( G => N218, D => N239, Q => 
                           REG_0_20_port);
   REG_reg_0_19_inst : DLH_X1 port map( G => N218, D => N238, Q => 
                           REG_0_19_port);
   REG_reg_0_18_inst : DLH_X1 port map( G => N218, D => N237, Q => 
                           REG_0_18_port);
   REG_reg_0_17_inst : DLH_X1 port map( G => N218, D => N236, Q => 
                           REG_0_17_port);
   REG_reg_0_16_inst : DLH_X1 port map( G => N218, D => N235, Q => 
                           REG_0_16_port);
   REG_reg_0_15_inst : DLH_X1 port map( G => N218, D => N234, Q => 
                           REG_0_15_port);
   REG_reg_0_14_inst : DLH_X1 port map( G => N218, D => N233, Q => 
                           REG_0_14_port);
   REG_reg_0_13_inst : DLH_X1 port map( G => N218, D => N232, Q => 
                           REG_0_13_port);
   REG_reg_0_12_inst : DLH_X1 port map( G => N218, D => N231, Q => 
                           REG_0_12_port);
   REG_reg_0_11_inst : DLH_X1 port map( G => N218, D => N230, Q => 
                           REG_0_11_port);
   REG_reg_0_10_inst : DLH_X1 port map( G => N218, D => N229, Q => 
                           REG_0_10_port);
   REG_reg_0_9_inst : DLH_X1 port map( G => N218, D => N228, Q => REG_0_9_port)
                           ;
   REG_reg_0_8_inst : DLH_X1 port map( G => N218, D => N227, Q => REG_0_8_port)
                           ;
   REG_reg_0_7_inst : DLH_X1 port map( G => N218, D => N226, Q => REG_0_7_port)
                           ;
   REG_reg_0_6_inst : DLH_X1 port map( G => N218, D => N225, Q => REG_0_6_port)
                           ;
   REG_reg_0_5_inst : DLH_X1 port map( G => N218, D => N224, Q => REG_0_5_port)
                           ;
   REG_reg_0_4_inst : DLH_X1 port map( G => N218, D => N223, Q => REG_0_4_port)
                           ;
   REG_reg_0_3_inst : DLH_X1 port map( G => N218, D => N222, Q => REG_0_3_port)
                           ;
   REG_reg_0_2_inst : DLH_X1 port map( G => N218, D => N221, Q => REG_0_2_port)
                           ;
   REG_reg_0_1_inst : DLH_X1 port map( G => N218, D => N220, Q => REG_0_1_port)
                           ;
   REG_reg_0_0_inst : DLH_X1 port map( G => N218, D => N219, Q => REG_0_0_port)
                           ;
   REG_reg_1_31_inst : DLH_X1 port map( G => n74, D => n1801, Q => 
                           REG_1_31_port);
   REG_reg_1_30_inst : DLH_X1 port map( G => n74, D => n1802, Q => 
                           REG_1_30_port);
   REG_reg_1_29_inst : DLH_X1 port map( G => n74, D => n1803, Q => 
                           REG_1_29_port);
   REG_reg_1_28_inst : DLH_X1 port map( G => n74, D => n1804, Q => 
                           REG_1_28_port);
   REG_reg_1_27_inst : DLH_X1 port map( G => n74, D => n1805, Q => 
                           REG_1_27_port);
   REG_reg_1_26_inst : DLH_X1 port map( G => n74, D => n1806, Q => 
                           REG_1_26_port);
   REG_reg_1_25_inst : DLH_X1 port map( G => n74, D => n1807, Q => 
                           REG_1_25_port);
   REG_reg_1_24_inst : DLH_X1 port map( G => n74, D => n1808, Q => 
                           REG_1_24_port);
   REG_reg_1_23_inst : DLH_X1 port map( G => n74, D => n1809, Q => 
                           REG_1_23_port);
   REG_reg_1_22_inst : DLH_X1 port map( G => n74, D => n1810, Q => 
                           REG_1_22_port);
   REG_reg_1_21_inst : DLH_X1 port map( G => n74, D => n1811, Q => 
                           REG_1_21_port);
   REG_reg_1_20_inst : DLH_X1 port map( G => n74, D => n1812, Q => 
                           REG_1_20_port);
   REG_reg_1_19_inst : DLH_X1 port map( G => n74, D => n1813, Q => 
                           REG_1_19_port);
   REG_reg_1_18_inst : DLH_X1 port map( G => n74, D => n1814, Q => 
                           REG_1_18_port);
   REG_reg_1_17_inst : DLH_X1 port map( G => n74, D => n1815, Q => 
                           REG_1_17_port);
   REG_reg_1_16_inst : DLH_X1 port map( G => n74, D => n1816, Q => 
                           REG_1_16_port);
   REG_reg_1_15_inst : DLH_X1 port map( G => n74, D => n1817, Q => 
                           REG_1_15_port);
   REG_reg_1_14_inst : DLH_X1 port map( G => n74, D => n1818, Q => 
                           REG_1_14_port);
   REG_reg_1_13_inst : DLH_X1 port map( G => n74, D => n1819, Q => 
                           REG_1_13_port);
   REG_reg_1_12_inst : DLH_X1 port map( G => n74, D => n1820, Q => 
                           REG_1_12_port);
   REG_reg_1_11_inst : DLH_X1 port map( G => n74, D => n1821, Q => 
                           REG_1_11_port);
   REG_reg_1_10_inst : DLH_X1 port map( G => n74, D => n1822, Q => 
                           REG_1_10_port);
   REG_reg_1_9_inst : DLH_X1 port map( G => n74, D => n1823, Q => REG_1_9_port)
                           ;
   REG_reg_1_8_inst : DLH_X1 port map( G => n74, D => n1824, Q => REG_1_8_port)
                           ;
   REG_reg_1_7_inst : DLH_X1 port map( G => n74, D => n1825, Q => REG_1_7_port)
                           ;
   REG_reg_1_6_inst : DLH_X1 port map( G => n74, D => n1826, Q => REG_1_6_port)
                           ;
   REG_reg_1_5_inst : DLH_X1 port map( G => n74, D => n1827, Q => REG_1_5_port)
                           ;
   REG_reg_1_4_inst : DLH_X1 port map( G => n74, D => n1828, Q => REG_1_4_port)
                           ;
   REG_reg_1_3_inst : DLH_X1 port map( G => n74, D => n1829, Q => REG_1_3_port)
                           ;
   REG_reg_1_2_inst : DLH_X1 port map( G => n74, D => n1830, Q => REG_1_2_port)
                           ;
   REG_reg_1_1_inst : DLH_X1 port map( G => n74, D => n1831, Q => REG_1_1_port)
                           ;
   REG_reg_1_0_inst : DLH_X1 port map( G => n74, D => n1832, Q => REG_1_0_port)
                           ;
   REG_reg_2_31_inst : DLH_X1 port map( G => n76, D => n1801, Q => 
                           REG_2_31_port);
   REG_reg_2_30_inst : DLH_X1 port map( G => n76, D => n1802, Q => 
                           REG_2_30_port);
   REG_reg_2_29_inst : DLH_X1 port map( G => n76, D => n1803, Q => 
                           REG_2_29_port);
   REG_reg_2_28_inst : DLH_X1 port map( G => n76, D => n1804, Q => 
                           REG_2_28_port);
   REG_reg_2_27_inst : DLH_X1 port map( G => n76, D => n1805, Q => 
                           REG_2_27_port);
   REG_reg_2_26_inst : DLH_X1 port map( G => n76, D => n1806, Q => 
                           REG_2_26_port);
   REG_reg_2_25_inst : DLH_X1 port map( G => n76, D => n1807, Q => 
                           REG_2_25_port);
   REG_reg_2_24_inst : DLH_X1 port map( G => n76, D => n1808, Q => 
                           REG_2_24_port);
   REG_reg_2_23_inst : DLH_X1 port map( G => n76, D => n1809, Q => 
                           REG_2_23_port);
   REG_reg_2_22_inst : DLH_X1 port map( G => n76, D => n1810, Q => 
                           REG_2_22_port);
   REG_reg_2_21_inst : DLH_X1 port map( G => n76, D => n1811, Q => 
                           REG_2_21_port);
   REG_reg_2_20_inst : DLH_X1 port map( G => n76, D => n1812, Q => 
                           REG_2_20_port);
   REG_reg_2_19_inst : DLH_X1 port map( G => n76, D => n1813, Q => 
                           REG_2_19_port);
   REG_reg_2_18_inst : DLH_X1 port map( G => n76, D => n1814, Q => 
                           REG_2_18_port);
   REG_reg_2_17_inst : DLH_X1 port map( G => n76, D => n1815, Q => 
                           REG_2_17_port);
   REG_reg_2_16_inst : DLH_X1 port map( G => n76, D => n1816, Q => 
                           REG_2_16_port);
   REG_reg_2_15_inst : DLH_X1 port map( G => n76, D => n1817, Q => 
                           REG_2_15_port);
   REG_reg_2_14_inst : DLH_X1 port map( G => n76, D => n1818, Q => 
                           REG_2_14_port);
   REG_reg_2_13_inst : DLH_X1 port map( G => n76, D => n1819, Q => 
                           REG_2_13_port);
   REG_reg_2_12_inst : DLH_X1 port map( G => n76, D => n1820, Q => 
                           REG_2_12_port);
   REG_reg_2_11_inst : DLH_X1 port map( G => n76, D => n1821, Q => 
                           REG_2_11_port);
   REG_reg_2_10_inst : DLH_X1 port map( G => n76, D => n1822, Q => 
                           REG_2_10_port);
   REG_reg_2_9_inst : DLH_X1 port map( G => n76, D => n1823, Q => REG_2_9_port)
                           ;
   REG_reg_2_8_inst : DLH_X1 port map( G => n76, D => n1824, Q => REG_2_8_port)
                           ;
   REG_reg_2_7_inst : DLH_X1 port map( G => n76, D => n1825, Q => REG_2_7_port)
                           ;
   REG_reg_2_6_inst : DLH_X1 port map( G => n76, D => n1826, Q => REG_2_6_port)
                           ;
   REG_reg_2_5_inst : DLH_X1 port map( G => n76, D => n1827, Q => REG_2_5_port)
                           ;
   REG_reg_2_4_inst : DLH_X1 port map( G => n76, D => n1828, Q => REG_2_4_port)
                           ;
   REG_reg_2_3_inst : DLH_X1 port map( G => n76, D => n1829, Q => REG_2_3_port)
                           ;
   REG_reg_2_2_inst : DLH_X1 port map( G => n76, D => n1830, Q => REG_2_2_port)
                           ;
   REG_reg_2_1_inst : DLH_X1 port map( G => n76, D => n1831, Q => REG_2_1_port)
                           ;
   REG_reg_2_0_inst : DLH_X1 port map( G => n76, D => n1832, Q => REG_2_0_port)
                           ;
   REG_reg_3_31_inst : DLH_X1 port map( G => n34, D => n1801, Q => 
                           REG_3_31_port);
   REG_reg_3_30_inst : DLH_X1 port map( G => n34, D => n1802, Q => 
                           REG_3_30_port);
   REG_reg_3_29_inst : DLH_X1 port map( G => n34, D => n1803, Q => 
                           REG_3_29_port);
   REG_reg_3_28_inst : DLH_X1 port map( G => n34, D => n1804, Q => 
                           REG_3_28_port);
   REG_reg_3_27_inst : DLH_X1 port map( G => n34, D => n1805, Q => 
                           REG_3_27_port);
   REG_reg_3_26_inst : DLH_X1 port map( G => n34, D => n1806, Q => 
                           REG_3_26_port);
   REG_reg_3_25_inst : DLH_X1 port map( G => n34, D => n1807, Q => 
                           REG_3_25_port);
   REG_reg_3_24_inst : DLH_X1 port map( G => n34, D => n1808, Q => 
                           REG_3_24_port);
   REG_reg_3_23_inst : DLH_X1 port map( G => n34, D => n1809, Q => 
                           REG_3_23_port);
   REG_reg_3_22_inst : DLH_X1 port map( G => n34, D => n1810, Q => 
                           REG_3_22_port);
   REG_reg_3_21_inst : DLH_X1 port map( G => n34, D => n1811, Q => 
                           REG_3_21_port);
   REG_reg_3_20_inst : DLH_X1 port map( G => n34, D => n1812, Q => 
                           REG_3_20_port);
   REG_reg_3_19_inst : DLH_X1 port map( G => n34, D => n1813, Q => 
                           REG_3_19_port);
   REG_reg_3_18_inst : DLH_X1 port map( G => n34, D => n1814, Q => 
                           REG_3_18_port);
   REG_reg_3_17_inst : DLH_X1 port map( G => n34, D => n1815, Q => 
                           REG_3_17_port);
   REG_reg_3_16_inst : DLH_X1 port map( G => n34, D => n1816, Q => 
                           REG_3_16_port);
   REG_reg_3_15_inst : DLH_X1 port map( G => n34, D => n1817, Q => 
                           REG_3_15_port);
   REG_reg_3_14_inst : DLH_X1 port map( G => n34, D => n1818, Q => 
                           REG_3_14_port);
   REG_reg_3_13_inst : DLH_X1 port map( G => n34, D => n1819, Q => 
                           REG_3_13_port);
   REG_reg_3_12_inst : DLH_X1 port map( G => n34, D => n1820, Q => 
                           REG_3_12_port);
   REG_reg_3_11_inst : DLH_X1 port map( G => n34, D => n1821, Q => 
                           REG_3_11_port);
   REG_reg_3_10_inst : DLH_X1 port map( G => n34, D => n1822, Q => 
                           REG_3_10_port);
   REG_reg_3_9_inst : DLH_X1 port map( G => n34, D => n1823, Q => REG_3_9_port)
                           ;
   REG_reg_3_8_inst : DLH_X1 port map( G => n34, D => n1824, Q => REG_3_8_port)
                           ;
   REG_reg_3_7_inst : DLH_X1 port map( G => n34, D => n1825, Q => REG_3_7_port)
                           ;
   REG_reg_3_6_inst : DLH_X1 port map( G => n34, D => n1826, Q => REG_3_6_port)
                           ;
   REG_reg_3_5_inst : DLH_X1 port map( G => n34, D => n1827, Q => REG_3_5_port)
                           ;
   REG_reg_3_4_inst : DLH_X1 port map( G => n34, D => n1828, Q => REG_3_4_port)
                           ;
   REG_reg_3_3_inst : DLH_X1 port map( G => n34, D => n1829, Q => REG_3_3_port)
                           ;
   REG_reg_3_2_inst : DLH_X1 port map( G => n34, D => n1830, Q => REG_3_2_port)
                           ;
   REG_reg_3_1_inst : DLH_X1 port map( G => n34, D => n1831, Q => REG_3_1_port)
                           ;
   REG_reg_3_0_inst : DLH_X1 port map( G => n34, D => n1832, Q => REG_3_0_port)
                           ;
   REG_reg_4_31_inst : DLH_X1 port map( G => n22, D => n1801, Q => 
                           REG_4_31_port);
   REG_reg_4_30_inst : DLH_X1 port map( G => n22, D => n1802, Q => 
                           REG_4_30_port);
   REG_reg_4_29_inst : DLH_X1 port map( G => n22, D => n1803, Q => 
                           REG_4_29_port);
   REG_reg_4_28_inst : DLH_X1 port map( G => n22, D => n1804, Q => 
                           REG_4_28_port);
   REG_reg_4_27_inst : DLH_X1 port map( G => n22, D => n1805, Q => 
                           REG_4_27_port);
   REG_reg_4_26_inst : DLH_X1 port map( G => n22, D => n1806, Q => 
                           REG_4_26_port);
   REG_reg_4_25_inst : DLH_X1 port map( G => n22, D => n1807, Q => 
                           REG_4_25_port);
   REG_reg_4_24_inst : DLH_X1 port map( G => n22, D => n1808, Q => 
                           REG_4_24_port);
   REG_reg_4_23_inst : DLH_X1 port map( G => n22, D => n1809, Q => 
                           REG_4_23_port);
   REG_reg_4_22_inst : DLH_X1 port map( G => n22, D => n1810, Q => 
                           REG_4_22_port);
   REG_reg_4_21_inst : DLH_X1 port map( G => n22, D => n1811, Q => 
                           REG_4_21_port);
   REG_reg_4_20_inst : DLH_X1 port map( G => n22, D => n1812, Q => 
                           REG_4_20_port);
   REG_reg_4_19_inst : DLH_X1 port map( G => n22, D => n1813, Q => 
                           REG_4_19_port);
   REG_reg_4_18_inst : DLH_X1 port map( G => n22, D => n1814, Q => 
                           REG_4_18_port);
   REG_reg_4_17_inst : DLH_X1 port map( G => n22, D => n1815, Q => 
                           REG_4_17_port);
   REG_reg_4_16_inst : DLH_X1 port map( G => n22, D => n1816, Q => 
                           REG_4_16_port);
   REG_reg_4_15_inst : DLH_X1 port map( G => n22, D => n1817, Q => 
                           REG_4_15_port);
   REG_reg_4_14_inst : DLH_X1 port map( G => n22, D => n1818, Q => 
                           REG_4_14_port);
   REG_reg_4_13_inst : DLH_X1 port map( G => n22, D => n1819, Q => 
                           REG_4_13_port);
   REG_reg_4_12_inst : DLH_X1 port map( G => n22, D => n1820, Q => 
                           REG_4_12_port);
   REG_reg_4_11_inst : DLH_X1 port map( G => n22, D => n1821, Q => 
                           REG_4_11_port);
   REG_reg_4_10_inst : DLH_X1 port map( G => n22, D => n1822, Q => 
                           REG_4_10_port);
   REG_reg_4_9_inst : DLH_X1 port map( G => n22, D => n1823, Q => REG_4_9_port)
                           ;
   REG_reg_4_8_inst : DLH_X1 port map( G => n22, D => n1824, Q => REG_4_8_port)
                           ;
   REG_reg_4_7_inst : DLH_X1 port map( G => n22, D => n1825, Q => REG_4_7_port)
                           ;
   REG_reg_4_6_inst : DLH_X1 port map( G => n22, D => n1826, Q => REG_4_6_port)
                           ;
   REG_reg_4_5_inst : DLH_X1 port map( G => n22, D => n1827, Q => REG_4_5_port)
                           ;
   REG_reg_4_4_inst : DLH_X1 port map( G => n22, D => n1828, Q => REG_4_4_port)
                           ;
   REG_reg_4_3_inst : DLH_X1 port map( G => n22, D => n1829, Q => REG_4_3_port)
                           ;
   REG_reg_4_2_inst : DLH_X1 port map( G => n22, D => n1830, Q => REG_4_2_port)
                           ;
   REG_reg_4_1_inst : DLH_X1 port map( G => n22, D => n1831, Q => REG_4_1_port)
                           ;
   REG_reg_4_0_inst : DLH_X1 port map( G => n22, D => n1832, Q => REG_4_0_port)
                           ;
   REG_reg_5_31_inst : DLH_X1 port map( G => n24, D => n1801, Q => 
                           REG_5_31_port);
   REG_reg_5_30_inst : DLH_X1 port map( G => n24, D => n1802, Q => 
                           REG_5_30_port);
   REG_reg_5_29_inst : DLH_X1 port map( G => n24, D => n1803, Q => 
                           REG_5_29_port);
   REG_reg_5_28_inst : DLH_X1 port map( G => n24, D => n1804, Q => 
                           REG_5_28_port);
   REG_reg_5_27_inst : DLH_X1 port map( G => n24, D => n1805, Q => 
                           REG_5_27_port);
   REG_reg_5_26_inst : DLH_X1 port map( G => n24, D => n1806, Q => 
                           REG_5_26_port);
   REG_reg_5_25_inst : DLH_X1 port map( G => n24, D => n1807, Q => 
                           REG_5_25_port);
   REG_reg_5_24_inst : DLH_X1 port map( G => n24, D => n1808, Q => 
                           REG_5_24_port);
   REG_reg_5_23_inst : DLH_X1 port map( G => n24, D => n1809, Q => 
                           REG_5_23_port);
   REG_reg_5_22_inst : DLH_X1 port map( G => n24, D => n1810, Q => 
                           REG_5_22_port);
   REG_reg_5_21_inst : DLH_X1 port map( G => n24, D => n1811, Q => 
                           REG_5_21_port);
   REG_reg_5_20_inst : DLH_X1 port map( G => n24, D => n1812, Q => 
                           REG_5_20_port);
   REG_reg_5_19_inst : DLH_X1 port map( G => n24, D => n1813, Q => 
                           REG_5_19_port);
   REG_reg_5_18_inst : DLH_X1 port map( G => n24, D => n1814, Q => 
                           REG_5_18_port);
   REG_reg_5_17_inst : DLH_X1 port map( G => n24, D => n1815, Q => 
                           REG_5_17_port);
   REG_reg_5_16_inst : DLH_X1 port map( G => n24, D => n1816, Q => 
                           REG_5_16_port);
   REG_reg_5_15_inst : DLH_X1 port map( G => n24, D => n1817, Q => 
                           REG_5_15_port);
   REG_reg_5_14_inst : DLH_X1 port map( G => n24, D => n1818, Q => 
                           REG_5_14_port);
   REG_reg_5_13_inst : DLH_X1 port map( G => n24, D => n1819, Q => 
                           REG_5_13_port);
   REG_reg_5_12_inst : DLH_X1 port map( G => n24, D => n1820, Q => 
                           REG_5_12_port);
   REG_reg_5_11_inst : DLH_X1 port map( G => n24, D => n1821, Q => 
                           REG_5_11_port);
   REG_reg_5_10_inst : DLH_X1 port map( G => n24, D => n1822, Q => 
                           REG_5_10_port);
   REG_reg_5_9_inst : DLH_X1 port map( G => n24, D => n1823, Q => REG_5_9_port)
                           ;
   REG_reg_5_8_inst : DLH_X1 port map( G => n24, D => n1824, Q => REG_5_8_port)
                           ;
   REG_reg_5_7_inst : DLH_X1 port map( G => n24, D => n1825, Q => REG_5_7_port)
                           ;
   REG_reg_5_6_inst : DLH_X1 port map( G => n24, D => n1826, Q => REG_5_6_port)
                           ;
   REG_reg_5_5_inst : DLH_X1 port map( G => n24, D => n1827, Q => REG_5_5_port)
                           ;
   REG_reg_5_4_inst : DLH_X1 port map( G => n24, D => n1828, Q => REG_5_4_port)
                           ;
   REG_reg_5_3_inst : DLH_X1 port map( G => n24, D => n1829, Q => REG_5_3_port)
                           ;
   REG_reg_5_2_inst : DLH_X1 port map( G => n24, D => n1830, Q => REG_5_2_port)
                           ;
   REG_reg_5_1_inst : DLH_X1 port map( G => n24, D => n1831, Q => REG_5_1_port)
                           ;
   REG_reg_5_0_inst : DLH_X1 port map( G => n24, D => n1832, Q => REG_5_0_port)
                           ;
   REG_reg_6_31_inst : DLH_X1 port map( G => n26, D => n1801, Q => 
                           REG_6_31_port);
   REG_reg_6_30_inst : DLH_X1 port map( G => n26, D => n1802, Q => 
                           REG_6_30_port);
   REG_reg_6_29_inst : DLH_X1 port map( G => n26, D => n1803, Q => 
                           REG_6_29_port);
   REG_reg_6_28_inst : DLH_X1 port map( G => n26, D => n1804, Q => 
                           REG_6_28_port);
   REG_reg_6_27_inst : DLH_X1 port map( G => n26, D => n1805, Q => 
                           REG_6_27_port);
   REG_reg_6_26_inst : DLH_X1 port map( G => n26, D => n1806, Q => 
                           REG_6_26_port);
   REG_reg_6_25_inst : DLH_X1 port map( G => n26, D => n1807, Q => 
                           REG_6_25_port);
   REG_reg_6_24_inst : DLH_X1 port map( G => n26, D => n1808, Q => 
                           REG_6_24_port);
   REG_reg_6_23_inst : DLH_X1 port map( G => n26, D => n1809, Q => 
                           REG_6_23_port);
   REG_reg_6_22_inst : DLH_X1 port map( G => n26, D => n1810, Q => 
                           REG_6_22_port);
   REG_reg_6_21_inst : DLH_X1 port map( G => n26, D => n1811, Q => 
                           REG_6_21_port);
   REG_reg_6_20_inst : DLH_X1 port map( G => n26, D => n1812, Q => 
                           REG_6_20_port);
   REG_reg_6_19_inst : DLH_X1 port map( G => n26, D => n1813, Q => 
                           REG_6_19_port);
   REG_reg_6_18_inst : DLH_X1 port map( G => n26, D => n1814, Q => 
                           REG_6_18_port);
   REG_reg_6_17_inst : DLH_X1 port map( G => n26, D => n1815, Q => 
                           REG_6_17_port);
   REG_reg_6_16_inst : DLH_X1 port map( G => n26, D => n1816, Q => 
                           REG_6_16_port);
   REG_reg_6_15_inst : DLH_X1 port map( G => n26, D => n1817, Q => 
                           REG_6_15_port);
   REG_reg_6_14_inst : DLH_X1 port map( G => n26, D => n1818, Q => 
                           REG_6_14_port);
   REG_reg_6_13_inst : DLH_X1 port map( G => n26, D => n1819, Q => 
                           REG_6_13_port);
   REG_reg_6_12_inst : DLH_X1 port map( G => n26, D => n1820, Q => 
                           REG_6_12_port);
   REG_reg_6_11_inst : DLH_X1 port map( G => n26, D => n1821, Q => 
                           REG_6_11_port);
   REG_reg_6_10_inst : DLH_X1 port map( G => n26, D => n1822, Q => 
                           REG_6_10_port);
   REG_reg_6_9_inst : DLH_X1 port map( G => n26, D => n1823, Q => REG_6_9_port)
                           ;
   REG_reg_6_8_inst : DLH_X1 port map( G => n26, D => n1824, Q => REG_6_8_port)
                           ;
   REG_reg_6_7_inst : DLH_X1 port map( G => n26, D => n1825, Q => REG_6_7_port)
                           ;
   REG_reg_6_6_inst : DLH_X1 port map( G => n26, D => n1826, Q => REG_6_6_port)
                           ;
   REG_reg_6_5_inst : DLH_X1 port map( G => n26, D => n1827, Q => REG_6_5_port)
                           ;
   REG_reg_6_4_inst : DLH_X1 port map( G => n26, D => n1828, Q => REG_6_4_port)
                           ;
   REG_reg_6_3_inst : DLH_X1 port map( G => n26, D => n1829, Q => REG_6_3_port)
                           ;
   REG_reg_6_2_inst : DLH_X1 port map( G => n26, D => n1830, Q => REG_6_2_port)
                           ;
   REG_reg_6_1_inst : DLH_X1 port map( G => n26, D => n1831, Q => REG_6_1_port)
                           ;
   REG_reg_6_0_inst : DLH_X1 port map( G => n26, D => n1832, Q => REG_6_0_port)
                           ;
   REG_reg_7_31_inst : DLH_X1 port map( G => n28, D => n1801, Q => 
                           REG_7_31_port);
   REG_reg_7_30_inst : DLH_X1 port map( G => n28, D => n1802, Q => 
                           REG_7_30_port);
   REG_reg_7_29_inst : DLH_X1 port map( G => n28, D => n1803, Q => 
                           REG_7_29_port);
   REG_reg_7_28_inst : DLH_X1 port map( G => n28, D => n1804, Q => 
                           REG_7_28_port);
   REG_reg_7_27_inst : DLH_X1 port map( G => n28, D => n1805, Q => 
                           REG_7_27_port);
   REG_reg_7_26_inst : DLH_X1 port map( G => n28, D => n1806, Q => 
                           REG_7_26_port);
   REG_reg_7_25_inst : DLH_X1 port map( G => n28, D => n1807, Q => 
                           REG_7_25_port);
   REG_reg_7_24_inst : DLH_X1 port map( G => n28, D => n1808, Q => 
                           REG_7_24_port);
   REG_reg_7_23_inst : DLH_X1 port map( G => n28, D => n1809, Q => 
                           REG_7_23_port);
   REG_reg_7_22_inst : DLH_X1 port map( G => n28, D => n1810, Q => 
                           REG_7_22_port);
   REG_reg_7_21_inst : DLH_X1 port map( G => n28, D => n1811, Q => 
                           REG_7_21_port);
   REG_reg_7_20_inst : DLH_X1 port map( G => n28, D => n1812, Q => 
                           REG_7_20_port);
   REG_reg_7_19_inst : DLH_X1 port map( G => n28, D => n1813, Q => 
                           REG_7_19_port);
   REG_reg_7_18_inst : DLH_X1 port map( G => n28, D => n1814, Q => 
                           REG_7_18_port);
   REG_reg_7_17_inst : DLH_X1 port map( G => n28, D => n1815, Q => 
                           REG_7_17_port);
   REG_reg_7_16_inst : DLH_X1 port map( G => n28, D => n1816, Q => 
                           REG_7_16_port);
   REG_reg_7_15_inst : DLH_X1 port map( G => n28, D => n1817, Q => 
                           REG_7_15_port);
   REG_reg_7_14_inst : DLH_X1 port map( G => n28, D => n1818, Q => 
                           REG_7_14_port);
   REG_reg_7_13_inst : DLH_X1 port map( G => n28, D => n1819, Q => 
                           REG_7_13_port);
   REG_reg_7_12_inst : DLH_X1 port map( G => n28, D => n1820, Q => 
                           REG_7_12_port);
   REG_reg_7_11_inst : DLH_X1 port map( G => n28, D => n1821, Q => 
                           REG_7_11_port);
   REG_reg_7_10_inst : DLH_X1 port map( G => n28, D => n1822, Q => 
                           REG_7_10_port);
   REG_reg_7_9_inst : DLH_X1 port map( G => n28, D => n1823, Q => REG_7_9_port)
                           ;
   REG_reg_7_8_inst : DLH_X1 port map( G => n28, D => n1824, Q => REG_7_8_port)
                           ;
   REG_reg_7_7_inst : DLH_X1 port map( G => n28, D => n1825, Q => REG_7_7_port)
                           ;
   REG_reg_7_6_inst : DLH_X1 port map( G => n28, D => n1826, Q => REG_7_6_port)
                           ;
   REG_reg_7_5_inst : DLH_X1 port map( G => n28, D => n1827, Q => REG_7_5_port)
                           ;
   REG_reg_7_4_inst : DLH_X1 port map( G => n28, D => n1828, Q => REG_7_4_port)
                           ;
   REG_reg_7_3_inst : DLH_X1 port map( G => n28, D => n1829, Q => REG_7_3_port)
                           ;
   REG_reg_7_2_inst : DLH_X1 port map( G => n28, D => n1830, Q => REG_7_2_port)
                           ;
   REG_reg_7_1_inst : DLH_X1 port map( G => n28, D => n1831, Q => REG_7_1_port)
                           ;
   REG_reg_7_0_inst : DLH_X1 port map( G => n28, D => n1832, Q => REG_7_0_port)
                           ;
   REG_reg_8_31_inst : DLH_X1 port map( G => n30, D => n1801, Q => 
                           REG_8_31_port);
   REG_reg_8_30_inst : DLH_X1 port map( G => n30, D => n1802, Q => 
                           REG_8_30_port);
   REG_reg_8_29_inst : DLH_X1 port map( G => n30, D => n1803, Q => 
                           REG_8_29_port);
   REG_reg_8_28_inst : DLH_X1 port map( G => n30, D => n1804, Q => 
                           REG_8_28_port);
   REG_reg_8_27_inst : DLH_X1 port map( G => n30, D => n1805, Q => 
                           REG_8_27_port);
   REG_reg_8_26_inst : DLH_X1 port map( G => n30, D => n1806, Q => 
                           REG_8_26_port);
   REG_reg_8_25_inst : DLH_X1 port map( G => n30, D => n1807, Q => 
                           REG_8_25_port);
   REG_reg_8_24_inst : DLH_X1 port map( G => n30, D => n1808, Q => 
                           REG_8_24_port);
   REG_reg_8_23_inst : DLH_X1 port map( G => n30, D => n1809, Q => 
                           REG_8_23_port);
   REG_reg_8_22_inst : DLH_X1 port map( G => n30, D => n1810, Q => 
                           REG_8_22_port);
   REG_reg_8_21_inst : DLH_X1 port map( G => n30, D => n1811, Q => 
                           REG_8_21_port);
   REG_reg_8_20_inst : DLH_X1 port map( G => n30, D => n1812, Q => 
                           REG_8_20_port);
   REG_reg_8_19_inst : DLH_X1 port map( G => n30, D => n1813, Q => 
                           REG_8_19_port);
   REG_reg_8_18_inst : DLH_X1 port map( G => n30, D => n1814, Q => 
                           REG_8_18_port);
   REG_reg_8_17_inst : DLH_X1 port map( G => n30, D => n1815, Q => 
                           REG_8_17_port);
   REG_reg_8_16_inst : DLH_X1 port map( G => n30, D => n1816, Q => 
                           REG_8_16_port);
   REG_reg_8_15_inst : DLH_X1 port map( G => n30, D => n1817, Q => 
                           REG_8_15_port);
   REG_reg_8_14_inst : DLH_X1 port map( G => n30, D => n1818, Q => 
                           REG_8_14_port);
   REG_reg_8_13_inst : DLH_X1 port map( G => n30, D => n1819, Q => 
                           REG_8_13_port);
   REG_reg_8_12_inst : DLH_X1 port map( G => n30, D => n1820, Q => 
                           REG_8_12_port);
   REG_reg_8_11_inst : DLH_X1 port map( G => n30, D => n1821, Q => 
                           REG_8_11_port);
   REG_reg_8_10_inst : DLH_X1 port map( G => n30, D => n1822, Q => 
                           REG_8_10_port);
   REG_reg_8_9_inst : DLH_X1 port map( G => n30, D => n1823, Q => REG_8_9_port)
                           ;
   REG_reg_8_8_inst : DLH_X1 port map( G => n30, D => n1824, Q => REG_8_8_port)
                           ;
   REG_reg_8_7_inst : DLH_X1 port map( G => n30, D => n1825, Q => REG_8_7_port)
                           ;
   REG_reg_8_6_inst : DLH_X1 port map( G => n30, D => n1826, Q => REG_8_6_port)
                           ;
   REG_reg_8_5_inst : DLH_X1 port map( G => n30, D => n1827, Q => REG_8_5_port)
                           ;
   REG_reg_8_4_inst : DLH_X1 port map( G => n30, D => n1828, Q => REG_8_4_port)
                           ;
   REG_reg_8_3_inst : DLH_X1 port map( G => n30, D => n1829, Q => REG_8_3_port)
                           ;
   REG_reg_8_2_inst : DLH_X1 port map( G => n30, D => n1830, Q => REG_8_2_port)
                           ;
   REG_reg_8_1_inst : DLH_X1 port map( G => n30, D => n1831, Q => REG_8_1_port)
                           ;
   REG_reg_8_0_inst : DLH_X1 port map( G => n30, D => n1832, Q => REG_8_0_port)
                           ;
   REG_reg_9_31_inst : DLH_X1 port map( G => n32, D => n1801, Q => 
                           REG_9_31_port);
   REG_reg_9_30_inst : DLH_X1 port map( G => n32, D => n1802, Q => 
                           REG_9_30_port);
   REG_reg_9_29_inst : DLH_X1 port map( G => n32, D => n1803, Q => 
                           REG_9_29_port);
   REG_reg_9_28_inst : DLH_X1 port map( G => n32, D => n1804, Q => 
                           REG_9_28_port);
   REG_reg_9_27_inst : DLH_X1 port map( G => n32, D => n1805, Q => 
                           REG_9_27_port);
   REG_reg_9_26_inst : DLH_X1 port map( G => n32, D => n1806, Q => 
                           REG_9_26_port);
   REG_reg_9_25_inst : DLH_X1 port map( G => n32, D => n1807, Q => 
                           REG_9_25_port);
   REG_reg_9_24_inst : DLH_X1 port map( G => n32, D => n1808, Q => 
                           REG_9_24_port);
   REG_reg_9_23_inst : DLH_X1 port map( G => n32, D => n1809, Q => 
                           REG_9_23_port);
   REG_reg_9_22_inst : DLH_X1 port map( G => n32, D => n1810, Q => 
                           REG_9_22_port);
   REG_reg_9_21_inst : DLH_X1 port map( G => n32, D => n1811, Q => 
                           REG_9_21_port);
   REG_reg_9_20_inst : DLH_X1 port map( G => n32, D => n1812, Q => 
                           REG_9_20_port);
   REG_reg_9_19_inst : DLH_X1 port map( G => n32, D => n1813, Q => 
                           REG_9_19_port);
   REG_reg_9_18_inst : DLH_X1 port map( G => n32, D => n1814, Q => 
                           REG_9_18_port);
   REG_reg_9_17_inst : DLH_X1 port map( G => n32, D => n1815, Q => 
                           REG_9_17_port);
   REG_reg_9_16_inst : DLH_X1 port map( G => n32, D => n1816, Q => 
                           REG_9_16_port);
   REG_reg_9_15_inst : DLH_X1 port map( G => n32, D => n1817, Q => 
                           REG_9_15_port);
   REG_reg_9_14_inst : DLH_X1 port map( G => n32, D => n1818, Q => 
                           REG_9_14_port);
   REG_reg_9_13_inst : DLH_X1 port map( G => n32, D => n1819, Q => 
                           REG_9_13_port);
   REG_reg_9_12_inst : DLH_X1 port map( G => n32, D => n1820, Q => 
                           REG_9_12_port);
   REG_reg_9_11_inst : DLH_X1 port map( G => n32, D => n1821, Q => 
                           REG_9_11_port);
   REG_reg_9_10_inst : DLH_X1 port map( G => n32, D => n1822, Q => 
                           REG_9_10_port);
   REG_reg_9_9_inst : DLH_X1 port map( G => n32, D => n1823, Q => REG_9_9_port)
                           ;
   REG_reg_9_8_inst : DLH_X1 port map( G => n32, D => n1824, Q => REG_9_8_port)
                           ;
   REG_reg_9_7_inst : DLH_X1 port map( G => n32, D => n1825, Q => REG_9_7_port)
                           ;
   REG_reg_9_6_inst : DLH_X1 port map( G => n32, D => n1826, Q => REG_9_6_port)
                           ;
   REG_reg_9_5_inst : DLH_X1 port map( G => n32, D => n1827, Q => REG_9_5_port)
                           ;
   REG_reg_9_4_inst : DLH_X1 port map( G => n32, D => n1828, Q => REG_9_4_port)
                           ;
   REG_reg_9_3_inst : DLH_X1 port map( G => n32, D => n1829, Q => REG_9_3_port)
                           ;
   REG_reg_9_2_inst : DLH_X1 port map( G => n32, D => n1830, Q => REG_9_2_port)
                           ;
   REG_reg_9_1_inst : DLH_X1 port map( G => n32, D => n1831, Q => REG_9_1_port)
                           ;
   REG_reg_9_0_inst : DLH_X1 port map( G => n32, D => n1832, Q => REG_9_0_port)
                           ;
   REG_reg_10_31_inst : DLH_X1 port map( G => n36, D => n1801, Q => 
                           REG_10_31_port);
   REG_reg_10_30_inst : DLH_X1 port map( G => n36, D => n1802, Q => 
                           REG_10_30_port);
   REG_reg_10_29_inst : DLH_X1 port map( G => n36, D => n1803, Q => 
                           REG_10_29_port);
   REG_reg_10_28_inst : DLH_X1 port map( G => n36, D => n1804, Q => 
                           REG_10_28_port);
   REG_reg_10_27_inst : DLH_X1 port map( G => n36, D => n1805, Q => 
                           REG_10_27_port);
   REG_reg_10_26_inst : DLH_X1 port map( G => n36, D => n1806, Q => 
                           REG_10_26_port);
   REG_reg_10_25_inst : DLH_X1 port map( G => n36, D => n1807, Q => 
                           REG_10_25_port);
   REG_reg_10_24_inst : DLH_X1 port map( G => n36, D => n1808, Q => 
                           REG_10_24_port);
   REG_reg_10_23_inst : DLH_X1 port map( G => n36, D => n1809, Q => 
                           REG_10_23_port);
   REG_reg_10_22_inst : DLH_X1 port map( G => n36, D => n1810, Q => 
                           REG_10_22_port);
   REG_reg_10_21_inst : DLH_X1 port map( G => n36, D => n1811, Q => 
                           REG_10_21_port);
   REG_reg_10_20_inst : DLH_X1 port map( G => n36, D => n1812, Q => 
                           REG_10_20_port);
   REG_reg_10_19_inst : DLH_X1 port map( G => n36, D => n1813, Q => 
                           REG_10_19_port);
   REG_reg_10_18_inst : DLH_X1 port map( G => n36, D => n1814, Q => 
                           REG_10_18_port);
   REG_reg_10_17_inst : DLH_X1 port map( G => n36, D => n1815, Q => 
                           REG_10_17_port);
   REG_reg_10_16_inst : DLH_X1 port map( G => n36, D => n1816, Q => 
                           REG_10_16_port);
   REG_reg_10_15_inst : DLH_X1 port map( G => n36, D => n1817, Q => 
                           REG_10_15_port);
   REG_reg_10_14_inst : DLH_X1 port map( G => n36, D => n1818, Q => 
                           REG_10_14_port);
   REG_reg_10_13_inst : DLH_X1 port map( G => n36, D => n1819, Q => 
                           REG_10_13_port);
   REG_reg_10_12_inst : DLH_X1 port map( G => n36, D => n1820, Q => 
                           REG_10_12_port);
   REG_reg_10_11_inst : DLH_X1 port map( G => n36, D => n1821, Q => 
                           REG_10_11_port);
   REG_reg_10_10_inst : DLH_X1 port map( G => n36, D => n1822, Q => 
                           REG_10_10_port);
   REG_reg_10_9_inst : DLH_X1 port map( G => n36, D => n1823, Q => 
                           REG_10_9_port);
   REG_reg_10_8_inst : DLH_X1 port map( G => n36, D => n1824, Q => 
                           REG_10_8_port);
   REG_reg_10_7_inst : DLH_X1 port map( G => n36, D => n1825, Q => 
                           REG_10_7_port);
   REG_reg_10_6_inst : DLH_X1 port map( G => n36, D => n1826, Q => 
                           REG_10_6_port);
   REG_reg_10_5_inst : DLH_X1 port map( G => n36, D => n1827, Q => 
                           REG_10_5_port);
   REG_reg_10_4_inst : DLH_X1 port map( G => n36, D => n1828, Q => 
                           REG_10_4_port);
   REG_reg_10_3_inst : DLH_X1 port map( G => n36, D => n1829, Q => 
                           REG_10_3_port);
   REG_reg_10_2_inst : DLH_X1 port map( G => n36, D => n1830, Q => 
                           REG_10_2_port);
   REG_reg_10_1_inst : DLH_X1 port map( G => n36, D => n1831, Q => 
                           REG_10_1_port);
   REG_reg_10_0_inst : DLH_X1 port map( G => n36, D => n1832, Q => 
                           REG_10_0_port);
   REG_reg_11_31_inst : DLH_X1 port map( G => n38, D => n1801, Q => 
                           REG_11_31_port);
   REG_reg_11_30_inst : DLH_X1 port map( G => n38, D => n1802, Q => 
                           REG_11_30_port);
   REG_reg_11_29_inst : DLH_X1 port map( G => n38, D => n1803, Q => 
                           REG_11_29_port);
   REG_reg_11_28_inst : DLH_X1 port map( G => n38, D => n1804, Q => 
                           REG_11_28_port);
   REG_reg_11_27_inst : DLH_X1 port map( G => n38, D => n1805, Q => 
                           REG_11_27_port);
   REG_reg_11_26_inst : DLH_X1 port map( G => n38, D => n1806, Q => 
                           REG_11_26_port);
   REG_reg_11_25_inst : DLH_X1 port map( G => n38, D => n1807, Q => 
                           REG_11_25_port);
   REG_reg_11_24_inst : DLH_X1 port map( G => n38, D => n1808, Q => 
                           REG_11_24_port);
   REG_reg_11_23_inst : DLH_X1 port map( G => n38, D => n1809, Q => 
                           REG_11_23_port);
   REG_reg_11_22_inst : DLH_X1 port map( G => n38, D => n1810, Q => 
                           REG_11_22_port);
   REG_reg_11_21_inst : DLH_X1 port map( G => n38, D => n1811, Q => 
                           REG_11_21_port);
   REG_reg_11_20_inst : DLH_X1 port map( G => n38, D => n1812, Q => 
                           REG_11_20_port);
   REG_reg_11_19_inst : DLH_X1 port map( G => n38, D => n1813, Q => 
                           REG_11_19_port);
   REG_reg_11_18_inst : DLH_X1 port map( G => n38, D => n1814, Q => 
                           REG_11_18_port);
   REG_reg_11_17_inst : DLH_X1 port map( G => n38, D => n1815, Q => 
                           REG_11_17_port);
   REG_reg_11_16_inst : DLH_X1 port map( G => n38, D => n1816, Q => 
                           REG_11_16_port);
   REG_reg_11_15_inst : DLH_X1 port map( G => n38, D => n1817, Q => 
                           REG_11_15_port);
   REG_reg_11_14_inst : DLH_X1 port map( G => n38, D => n1818, Q => 
                           REG_11_14_port);
   REG_reg_11_13_inst : DLH_X1 port map( G => n38, D => n1819, Q => 
                           REG_11_13_port);
   REG_reg_11_12_inst : DLH_X1 port map( G => n38, D => n1820, Q => 
                           REG_11_12_port);
   REG_reg_11_11_inst : DLH_X1 port map( G => n38, D => n1821, Q => 
                           REG_11_11_port);
   REG_reg_11_10_inst : DLH_X1 port map( G => n38, D => n1822, Q => 
                           REG_11_10_port);
   REG_reg_11_9_inst : DLH_X1 port map( G => n38, D => n1823, Q => 
                           REG_11_9_port);
   REG_reg_11_8_inst : DLH_X1 port map( G => n38, D => n1824, Q => 
                           REG_11_8_port);
   REG_reg_11_7_inst : DLH_X1 port map( G => n38, D => n1825, Q => 
                           REG_11_7_port);
   REG_reg_11_6_inst : DLH_X1 port map( G => n38, D => n1826, Q => 
                           REG_11_6_port);
   REG_reg_11_5_inst : DLH_X1 port map( G => n38, D => n1827, Q => 
                           REG_11_5_port);
   REG_reg_11_4_inst : DLH_X1 port map( G => n38, D => n1828, Q => 
                           REG_11_4_port);
   REG_reg_11_3_inst : DLH_X1 port map( G => n38, D => n1829, Q => 
                           REG_11_3_port);
   REG_reg_11_2_inst : DLH_X1 port map( G => n38, D => n1830, Q => 
                           REG_11_2_port);
   REG_reg_11_1_inst : DLH_X1 port map( G => n38, D => n1831, Q => 
                           REG_11_1_port);
   REG_reg_11_0_inst : DLH_X1 port map( G => n38, D => n1832, Q => 
                           REG_11_0_port);
   REG_reg_12_31_inst : DLH_X1 port map( G => n40, D => n1801, Q => 
                           REG_12_31_port);
   REG_reg_12_30_inst : DLH_X1 port map( G => n40, D => n1802, Q => 
                           REG_12_30_port);
   REG_reg_12_29_inst : DLH_X1 port map( G => n40, D => n1803, Q => 
                           REG_12_29_port);
   REG_reg_12_28_inst : DLH_X1 port map( G => n40, D => n1804, Q => 
                           REG_12_28_port);
   REG_reg_12_27_inst : DLH_X1 port map( G => n40, D => n1805, Q => 
                           REG_12_27_port);
   REG_reg_12_26_inst : DLH_X1 port map( G => n40, D => n1806, Q => 
                           REG_12_26_port);
   REG_reg_12_25_inst : DLH_X1 port map( G => n40, D => n1807, Q => 
                           REG_12_25_port);
   REG_reg_12_24_inst : DLH_X1 port map( G => n40, D => n1808, Q => 
                           REG_12_24_port);
   REG_reg_12_23_inst : DLH_X1 port map( G => n40, D => n1809, Q => 
                           REG_12_23_port);
   REG_reg_12_22_inst : DLH_X1 port map( G => n40, D => n1810, Q => 
                           REG_12_22_port);
   REG_reg_12_21_inst : DLH_X1 port map( G => n40, D => n1811, Q => 
                           REG_12_21_port);
   REG_reg_12_20_inst : DLH_X1 port map( G => n40, D => n1812, Q => 
                           REG_12_20_port);
   REG_reg_12_19_inst : DLH_X1 port map( G => n40, D => n1813, Q => 
                           REG_12_19_port);
   REG_reg_12_18_inst : DLH_X1 port map( G => n40, D => n1814, Q => 
                           REG_12_18_port);
   REG_reg_12_17_inst : DLH_X1 port map( G => n40, D => n1815, Q => 
                           REG_12_17_port);
   REG_reg_12_16_inst : DLH_X1 port map( G => n40, D => n1816, Q => 
                           REG_12_16_port);
   REG_reg_12_15_inst : DLH_X1 port map( G => n40, D => n1817, Q => 
                           REG_12_15_port);
   REG_reg_12_14_inst : DLH_X1 port map( G => n40, D => n1818, Q => 
                           REG_12_14_port);
   REG_reg_12_13_inst : DLH_X1 port map( G => n40, D => n1819, Q => 
                           REG_12_13_port);
   REG_reg_12_12_inst : DLH_X1 port map( G => n40, D => n1820, Q => 
                           REG_12_12_port);
   REG_reg_12_11_inst : DLH_X1 port map( G => n40, D => n1821, Q => 
                           REG_12_11_port);
   REG_reg_12_10_inst : DLH_X1 port map( G => n40, D => n1822, Q => 
                           REG_12_10_port);
   REG_reg_12_9_inst : DLH_X1 port map( G => n40, D => n1823, Q => 
                           REG_12_9_port);
   REG_reg_12_8_inst : DLH_X1 port map( G => n40, D => n1824, Q => 
                           REG_12_8_port);
   REG_reg_12_7_inst : DLH_X1 port map( G => n40, D => n1825, Q => 
                           REG_12_7_port);
   REG_reg_12_6_inst : DLH_X1 port map( G => n40, D => n1826, Q => 
                           REG_12_6_port);
   REG_reg_12_5_inst : DLH_X1 port map( G => n40, D => n1827, Q => 
                           REG_12_5_port);
   REG_reg_12_4_inst : DLH_X1 port map( G => n40, D => n1828, Q => 
                           REG_12_4_port);
   REG_reg_12_3_inst : DLH_X1 port map( G => n40, D => n1829, Q => 
                           REG_12_3_port);
   REG_reg_12_2_inst : DLH_X1 port map( G => n40, D => n1830, Q => 
                           REG_12_2_port);
   REG_reg_12_1_inst : DLH_X1 port map( G => n40, D => n1831, Q => 
                           REG_12_1_port);
   REG_reg_12_0_inst : DLH_X1 port map( G => n40, D => n1832, Q => 
                           REG_12_0_port);
   REG_reg_13_31_inst : DLH_X1 port map( G => n42, D => n1801, Q => 
                           REG_13_31_port);
   REG_reg_13_30_inst : DLH_X1 port map( G => n42, D => n1802, Q => 
                           REG_13_30_port);
   REG_reg_13_29_inst : DLH_X1 port map( G => n42, D => n1803, Q => 
                           REG_13_29_port);
   REG_reg_13_28_inst : DLH_X1 port map( G => n42, D => n1804, Q => 
                           REG_13_28_port);
   REG_reg_13_27_inst : DLH_X1 port map( G => n42, D => n1805, Q => 
                           REG_13_27_port);
   REG_reg_13_26_inst : DLH_X1 port map( G => n42, D => n1806, Q => 
                           REG_13_26_port);
   REG_reg_13_25_inst : DLH_X1 port map( G => n42, D => n1807, Q => 
                           REG_13_25_port);
   REG_reg_13_24_inst : DLH_X1 port map( G => n42, D => n1808, Q => 
                           REG_13_24_port);
   REG_reg_13_23_inst : DLH_X1 port map( G => n42, D => n1809, Q => 
                           REG_13_23_port);
   REG_reg_13_22_inst : DLH_X1 port map( G => n42, D => n1810, Q => 
                           REG_13_22_port);
   REG_reg_13_21_inst : DLH_X1 port map( G => n42, D => n1811, Q => 
                           REG_13_21_port);
   REG_reg_13_20_inst : DLH_X1 port map( G => n42, D => n1812, Q => 
                           REG_13_20_port);
   REG_reg_13_19_inst : DLH_X1 port map( G => n42, D => n1813, Q => 
                           REG_13_19_port);
   REG_reg_13_18_inst : DLH_X1 port map( G => n42, D => n1814, Q => 
                           REG_13_18_port);
   REG_reg_13_17_inst : DLH_X1 port map( G => n42, D => n1815, Q => 
                           REG_13_17_port);
   REG_reg_13_16_inst : DLH_X1 port map( G => n42, D => n1816, Q => 
                           REG_13_16_port);
   REG_reg_13_15_inst : DLH_X1 port map( G => n42, D => n1817, Q => 
                           REG_13_15_port);
   REG_reg_13_14_inst : DLH_X1 port map( G => n42, D => n1818, Q => 
                           REG_13_14_port);
   REG_reg_13_13_inst : DLH_X1 port map( G => n42, D => n1819, Q => 
                           REG_13_13_port);
   REG_reg_13_12_inst : DLH_X1 port map( G => n42, D => n1820, Q => 
                           REG_13_12_port);
   REG_reg_13_11_inst : DLH_X1 port map( G => n42, D => n1821, Q => 
                           REG_13_11_port);
   REG_reg_13_10_inst : DLH_X1 port map( G => n42, D => n1822, Q => 
                           REG_13_10_port);
   REG_reg_13_9_inst : DLH_X1 port map( G => n42, D => n1823, Q => 
                           REG_13_9_port);
   REG_reg_13_8_inst : DLH_X1 port map( G => n42, D => n1824, Q => 
                           REG_13_8_port);
   REG_reg_13_7_inst : DLH_X1 port map( G => n42, D => n1825, Q => 
                           REG_13_7_port);
   REG_reg_13_6_inst : DLH_X1 port map( G => n42, D => n1826, Q => 
                           REG_13_6_port);
   REG_reg_13_5_inst : DLH_X1 port map( G => n42, D => n1827, Q => 
                           REG_13_5_port);
   REG_reg_13_4_inst : DLH_X1 port map( G => n42, D => n1828, Q => 
                           REG_13_4_port);
   REG_reg_13_3_inst : DLH_X1 port map( G => n42, D => n1829, Q => 
                           REG_13_3_port);
   REG_reg_13_2_inst : DLH_X1 port map( G => n42, D => n1830, Q => 
                           REG_13_2_port);
   REG_reg_13_1_inst : DLH_X1 port map( G => n42, D => n1831, Q => 
                           REG_13_1_port);
   REG_reg_13_0_inst : DLH_X1 port map( G => n42, D => n1832, Q => 
                           REG_13_0_port);
   REG_reg_14_31_inst : DLH_X1 port map( G => n44, D => n1801, Q => 
                           REG_14_31_port);
   REG_reg_14_30_inst : DLH_X1 port map( G => n44, D => n1802, Q => 
                           REG_14_30_port);
   REG_reg_14_29_inst : DLH_X1 port map( G => n44, D => n1803, Q => 
                           REG_14_29_port);
   REG_reg_14_28_inst : DLH_X1 port map( G => n44, D => n1804, Q => 
                           REG_14_28_port);
   REG_reg_14_27_inst : DLH_X1 port map( G => n44, D => n1805, Q => 
                           REG_14_27_port);
   REG_reg_14_26_inst : DLH_X1 port map( G => n44, D => n1806, Q => 
                           REG_14_26_port);
   REG_reg_14_25_inst : DLH_X1 port map( G => n44, D => n1807, Q => 
                           REG_14_25_port);
   REG_reg_14_24_inst : DLH_X1 port map( G => n44, D => n1808, Q => 
                           REG_14_24_port);
   REG_reg_14_23_inst : DLH_X1 port map( G => n44, D => n1809, Q => 
                           REG_14_23_port);
   REG_reg_14_22_inst : DLH_X1 port map( G => n44, D => n1810, Q => 
                           REG_14_22_port);
   REG_reg_14_21_inst : DLH_X1 port map( G => n44, D => n1811, Q => 
                           REG_14_21_port);
   REG_reg_14_20_inst : DLH_X1 port map( G => n44, D => n1812, Q => 
                           REG_14_20_port);
   REG_reg_14_19_inst : DLH_X1 port map( G => n44, D => n1813, Q => 
                           REG_14_19_port);
   REG_reg_14_18_inst : DLH_X1 port map( G => n44, D => n1814, Q => 
                           REG_14_18_port);
   REG_reg_14_17_inst : DLH_X1 port map( G => n44, D => n1815, Q => 
                           REG_14_17_port);
   REG_reg_14_16_inst : DLH_X1 port map( G => n44, D => n1816, Q => 
                           REG_14_16_port);
   REG_reg_14_15_inst : DLH_X1 port map( G => n44, D => n1817, Q => 
                           REG_14_15_port);
   REG_reg_14_14_inst : DLH_X1 port map( G => n44, D => n1818, Q => 
                           REG_14_14_port);
   REG_reg_14_13_inst : DLH_X1 port map( G => n44, D => n1819, Q => 
                           REG_14_13_port);
   REG_reg_14_12_inst : DLH_X1 port map( G => n44, D => n1820, Q => 
                           REG_14_12_port);
   REG_reg_14_11_inst : DLH_X1 port map( G => n44, D => n1821, Q => 
                           REG_14_11_port);
   REG_reg_14_10_inst : DLH_X1 port map( G => n44, D => n1822, Q => 
                           REG_14_10_port);
   REG_reg_14_9_inst : DLH_X1 port map( G => n44, D => n1823, Q => 
                           REG_14_9_port);
   REG_reg_14_8_inst : DLH_X1 port map( G => n44, D => n1824, Q => 
                           REG_14_8_port);
   REG_reg_14_7_inst : DLH_X1 port map( G => n44, D => n1825, Q => 
                           REG_14_7_port);
   REG_reg_14_6_inst : DLH_X1 port map( G => n44, D => n1826, Q => 
                           REG_14_6_port);
   REG_reg_14_5_inst : DLH_X1 port map( G => n44, D => n1827, Q => 
                           REG_14_5_port);
   REG_reg_14_4_inst : DLH_X1 port map( G => n44, D => n1828, Q => 
                           REG_14_4_port);
   REG_reg_14_3_inst : DLH_X1 port map( G => n44, D => n1829, Q => 
                           REG_14_3_port);
   REG_reg_14_2_inst : DLH_X1 port map( G => n44, D => n1830, Q => 
                           REG_14_2_port);
   REG_reg_14_1_inst : DLH_X1 port map( G => n44, D => n1831, Q => 
                           REG_14_1_port);
   REG_reg_14_0_inst : DLH_X1 port map( G => n44, D => n1832, Q => 
                           REG_14_0_port);
   REG_reg_15_31_inst : DLH_X1 port map( G => n46, D => n1801, Q => 
                           REG_15_31_port);
   REG_reg_15_30_inst : DLH_X1 port map( G => n46, D => n1802, Q => 
                           REG_15_30_port);
   REG_reg_15_29_inst : DLH_X1 port map( G => n46, D => n1803, Q => 
                           REG_15_29_port);
   REG_reg_15_28_inst : DLH_X1 port map( G => n46, D => n1804, Q => 
                           REG_15_28_port);
   REG_reg_15_27_inst : DLH_X1 port map( G => n46, D => n1805, Q => 
                           REG_15_27_port);
   REG_reg_15_26_inst : DLH_X1 port map( G => n46, D => n1806, Q => 
                           REG_15_26_port);
   REG_reg_15_25_inst : DLH_X1 port map( G => n46, D => n1807, Q => 
                           REG_15_25_port);
   REG_reg_15_24_inst : DLH_X1 port map( G => n46, D => n1808, Q => 
                           REG_15_24_port);
   REG_reg_15_23_inst : DLH_X1 port map( G => n46, D => n1809, Q => 
                           REG_15_23_port);
   REG_reg_15_22_inst : DLH_X1 port map( G => n46, D => n1810, Q => 
                           REG_15_22_port);
   REG_reg_15_21_inst : DLH_X1 port map( G => n46, D => n1811, Q => 
                           REG_15_21_port);
   REG_reg_15_20_inst : DLH_X1 port map( G => n46, D => n1812, Q => 
                           REG_15_20_port);
   REG_reg_15_19_inst : DLH_X1 port map( G => n46, D => n1813, Q => 
                           REG_15_19_port);
   REG_reg_15_18_inst : DLH_X1 port map( G => n46, D => n1814, Q => 
                           REG_15_18_port);
   REG_reg_15_17_inst : DLH_X1 port map( G => n46, D => n1815, Q => 
                           REG_15_17_port);
   REG_reg_15_16_inst : DLH_X1 port map( G => n46, D => n1816, Q => 
                           REG_15_16_port);
   REG_reg_15_15_inst : DLH_X1 port map( G => n46, D => n1817, Q => 
                           REG_15_15_port);
   REG_reg_15_14_inst : DLH_X1 port map( G => n46, D => n1818, Q => 
                           REG_15_14_port);
   REG_reg_15_13_inst : DLH_X1 port map( G => n46, D => n1819, Q => 
                           REG_15_13_port);
   REG_reg_15_12_inst : DLH_X1 port map( G => n46, D => n1820, Q => 
                           REG_15_12_port);
   REG_reg_15_11_inst : DLH_X1 port map( G => n46, D => n1821, Q => 
                           REG_15_11_port);
   REG_reg_15_10_inst : DLH_X1 port map( G => n46, D => n1822, Q => 
                           REG_15_10_port);
   REG_reg_15_9_inst : DLH_X1 port map( G => n46, D => n1823, Q => 
                           REG_15_9_port);
   REG_reg_15_8_inst : DLH_X1 port map( G => n46, D => n1824, Q => 
                           REG_15_8_port);
   REG_reg_15_7_inst : DLH_X1 port map( G => n46, D => n1825, Q => 
                           REG_15_7_port);
   REG_reg_15_6_inst : DLH_X1 port map( G => n46, D => n1826, Q => 
                           REG_15_6_port);
   REG_reg_15_5_inst : DLH_X1 port map( G => n46, D => n1827, Q => 
                           REG_15_5_port);
   REG_reg_15_4_inst : DLH_X1 port map( G => n46, D => n1828, Q => 
                           REG_15_4_port);
   REG_reg_15_3_inst : DLH_X1 port map( G => n46, D => n1829, Q => 
                           REG_15_3_port);
   REG_reg_15_2_inst : DLH_X1 port map( G => n46, D => n1830, Q => 
                           REG_15_2_port);
   REG_reg_15_1_inst : DLH_X1 port map( G => n46, D => n1831, Q => 
                           REG_15_1_port);
   REG_reg_15_0_inst : DLH_X1 port map( G => n46, D => n1832, Q => 
                           REG_15_0_port);
   REG_reg_16_31_inst : DLH_X1 port map( G => n48, D => n1801, Q => 
                           REG_16_31_port);
   REG_reg_16_30_inst : DLH_X1 port map( G => n48, D => n1802, Q => 
                           REG_16_30_port);
   REG_reg_16_29_inst : DLH_X1 port map( G => n48, D => n1803, Q => 
                           REG_16_29_port);
   REG_reg_16_28_inst : DLH_X1 port map( G => n48, D => n1804, Q => 
                           REG_16_28_port);
   REG_reg_16_27_inst : DLH_X1 port map( G => n48, D => n1805, Q => 
                           REG_16_27_port);
   REG_reg_16_26_inst : DLH_X1 port map( G => n48, D => n1806, Q => 
                           REG_16_26_port);
   REG_reg_16_25_inst : DLH_X1 port map( G => n48, D => n1807, Q => 
                           REG_16_25_port);
   REG_reg_16_24_inst : DLH_X1 port map( G => n48, D => n1808, Q => 
                           REG_16_24_port);
   REG_reg_16_23_inst : DLH_X1 port map( G => n48, D => n1809, Q => 
                           REG_16_23_port);
   REG_reg_16_22_inst : DLH_X1 port map( G => n48, D => n1810, Q => 
                           REG_16_22_port);
   REG_reg_16_21_inst : DLH_X1 port map( G => n48, D => n1811, Q => 
                           REG_16_21_port);
   REG_reg_16_20_inst : DLH_X1 port map( G => n48, D => n1812, Q => 
                           REG_16_20_port);
   REG_reg_16_19_inst : DLH_X1 port map( G => n48, D => n1813, Q => 
                           REG_16_19_port);
   REG_reg_16_18_inst : DLH_X1 port map( G => n48, D => n1814, Q => 
                           REG_16_18_port);
   REG_reg_16_17_inst : DLH_X1 port map( G => n48, D => n1815, Q => 
                           REG_16_17_port);
   REG_reg_16_16_inst : DLH_X1 port map( G => n48, D => n1816, Q => 
                           REG_16_16_port);
   REG_reg_16_15_inst : DLH_X1 port map( G => n48, D => n1817, Q => 
                           REG_16_15_port);
   REG_reg_16_14_inst : DLH_X1 port map( G => n48, D => n1818, Q => 
                           REG_16_14_port);
   REG_reg_16_13_inst : DLH_X1 port map( G => n48, D => n1819, Q => 
                           REG_16_13_port);
   REG_reg_16_12_inst : DLH_X1 port map( G => n48, D => n1820, Q => 
                           REG_16_12_port);
   REG_reg_16_11_inst : DLH_X1 port map( G => n48, D => n1821, Q => 
                           REG_16_11_port);
   REG_reg_16_10_inst : DLH_X1 port map( G => n48, D => n1822, Q => 
                           REG_16_10_port);
   REG_reg_16_9_inst : DLH_X1 port map( G => n48, D => n1823, Q => 
                           REG_16_9_port);
   REG_reg_16_8_inst : DLH_X1 port map( G => n48, D => n1824, Q => 
                           REG_16_8_port);
   REG_reg_16_7_inst : DLH_X1 port map( G => n48, D => n1825, Q => 
                           REG_16_7_port);
   REG_reg_16_6_inst : DLH_X1 port map( G => n48, D => n1826, Q => 
                           REG_16_6_port);
   REG_reg_16_5_inst : DLH_X1 port map( G => n48, D => n1827, Q => 
                           REG_16_5_port);
   REG_reg_16_4_inst : DLH_X1 port map( G => n48, D => n1828, Q => 
                           REG_16_4_port);
   REG_reg_16_3_inst : DLH_X1 port map( G => n48, D => n1829, Q => 
                           REG_16_3_port);
   REG_reg_16_2_inst : DLH_X1 port map( G => n48, D => n1830, Q => 
                           REG_16_2_port);
   REG_reg_16_1_inst : DLH_X1 port map( G => n48, D => n1831, Q => 
                           REG_16_1_port);
   REG_reg_16_0_inst : DLH_X1 port map( G => n48, D => n1832, Q => 
                           REG_16_0_port);
   REG_reg_17_31_inst : DLH_X1 port map( G => n50, D => n1801, Q => 
                           REG_17_31_port);
   REG_reg_17_30_inst : DLH_X1 port map( G => n50, D => n1802, Q => 
                           REG_17_30_port);
   REG_reg_17_29_inst : DLH_X1 port map( G => n50, D => n1803, Q => 
                           REG_17_29_port);
   REG_reg_17_28_inst : DLH_X1 port map( G => n50, D => n1804, Q => 
                           REG_17_28_port);
   REG_reg_17_27_inst : DLH_X1 port map( G => n50, D => n1805, Q => 
                           REG_17_27_port);
   REG_reg_17_26_inst : DLH_X1 port map( G => n50, D => n1806, Q => 
                           REG_17_26_port);
   REG_reg_17_25_inst : DLH_X1 port map( G => n50, D => n1807, Q => 
                           REG_17_25_port);
   REG_reg_17_24_inst : DLH_X1 port map( G => n50, D => n1808, Q => 
                           REG_17_24_port);
   REG_reg_17_23_inst : DLH_X1 port map( G => n50, D => n1809, Q => 
                           REG_17_23_port);
   REG_reg_17_22_inst : DLH_X1 port map( G => n50, D => n1810, Q => 
                           REG_17_22_port);
   REG_reg_17_21_inst : DLH_X1 port map( G => n50, D => n1811, Q => 
                           REG_17_21_port);
   REG_reg_17_20_inst : DLH_X1 port map( G => n50, D => n1812, Q => 
                           REG_17_20_port);
   REG_reg_17_19_inst : DLH_X1 port map( G => n50, D => n1813, Q => 
                           REG_17_19_port);
   REG_reg_17_18_inst : DLH_X1 port map( G => n50, D => n1814, Q => 
                           REG_17_18_port);
   REG_reg_17_17_inst : DLH_X1 port map( G => n50, D => n1815, Q => 
                           REG_17_17_port);
   REG_reg_17_16_inst : DLH_X1 port map( G => n50, D => n1816, Q => 
                           REG_17_16_port);
   REG_reg_17_15_inst : DLH_X1 port map( G => n50, D => n1817, Q => 
                           REG_17_15_port);
   REG_reg_17_14_inst : DLH_X1 port map( G => n50, D => n1818, Q => 
                           REG_17_14_port);
   REG_reg_17_13_inst : DLH_X1 port map( G => n50, D => n1819, Q => 
                           REG_17_13_port);
   REG_reg_17_12_inst : DLH_X1 port map( G => n50, D => n1820, Q => 
                           REG_17_12_port);
   REG_reg_17_11_inst : DLH_X1 port map( G => n50, D => n1821, Q => 
                           REG_17_11_port);
   REG_reg_17_10_inst : DLH_X1 port map( G => n50, D => n1822, Q => 
                           REG_17_10_port);
   REG_reg_17_9_inst : DLH_X1 port map( G => n50, D => n1823, Q => 
                           REG_17_9_port);
   REG_reg_17_8_inst : DLH_X1 port map( G => n50, D => n1824, Q => 
                           REG_17_8_port);
   REG_reg_17_7_inst : DLH_X1 port map( G => n50, D => n1825, Q => 
                           REG_17_7_port);
   REG_reg_17_6_inst : DLH_X1 port map( G => n50, D => n1826, Q => 
                           REG_17_6_port);
   REG_reg_17_5_inst : DLH_X1 port map( G => n50, D => n1827, Q => 
                           REG_17_5_port);
   REG_reg_17_4_inst : DLH_X1 port map( G => n50, D => n1828, Q => 
                           REG_17_4_port);
   REG_reg_17_3_inst : DLH_X1 port map( G => n50, D => n1829, Q => 
                           REG_17_3_port);
   REG_reg_17_2_inst : DLH_X1 port map( G => n50, D => n1830, Q => 
                           REG_17_2_port);
   REG_reg_17_1_inst : DLH_X1 port map( G => n50, D => n1831, Q => 
                           REG_17_1_port);
   REG_reg_17_0_inst : DLH_X1 port map( G => n50, D => n1832, Q => 
                           REG_17_0_port);
   REG_reg_18_31_inst : DLH_X1 port map( G => n52, D => n1801, Q => 
                           REG_18_31_port);
   REG_reg_18_30_inst : DLH_X1 port map( G => n52, D => n1802, Q => 
                           REG_18_30_port);
   REG_reg_18_29_inst : DLH_X1 port map( G => n52, D => n1803, Q => 
                           REG_18_29_port);
   REG_reg_18_28_inst : DLH_X1 port map( G => n52, D => n1804, Q => 
                           REG_18_28_port);
   REG_reg_18_27_inst : DLH_X1 port map( G => n52, D => n1805, Q => 
                           REG_18_27_port);
   REG_reg_18_26_inst : DLH_X1 port map( G => n52, D => n1806, Q => 
                           REG_18_26_port);
   REG_reg_18_25_inst : DLH_X1 port map( G => n52, D => n1807, Q => 
                           REG_18_25_port);
   REG_reg_18_24_inst : DLH_X1 port map( G => n52, D => n1808, Q => 
                           REG_18_24_port);
   REG_reg_18_23_inst : DLH_X1 port map( G => n52, D => n1809, Q => 
                           REG_18_23_port);
   REG_reg_18_22_inst : DLH_X1 port map( G => n52, D => n1810, Q => 
                           REG_18_22_port);
   REG_reg_18_21_inst : DLH_X1 port map( G => n52, D => n1811, Q => 
                           REG_18_21_port);
   REG_reg_18_20_inst : DLH_X1 port map( G => n52, D => n1812, Q => 
                           REG_18_20_port);
   REG_reg_18_19_inst : DLH_X1 port map( G => n52, D => n1813, Q => 
                           REG_18_19_port);
   REG_reg_18_18_inst : DLH_X1 port map( G => n52, D => n1814, Q => 
                           REG_18_18_port);
   REG_reg_18_17_inst : DLH_X1 port map( G => n52, D => n1815, Q => 
                           REG_18_17_port);
   REG_reg_18_16_inst : DLH_X1 port map( G => n52, D => n1816, Q => 
                           REG_18_16_port);
   REG_reg_18_15_inst : DLH_X1 port map( G => n52, D => n1817, Q => 
                           REG_18_15_port);
   REG_reg_18_14_inst : DLH_X1 port map( G => n52, D => n1818, Q => 
                           REG_18_14_port);
   REG_reg_18_13_inst : DLH_X1 port map( G => n52, D => n1819, Q => 
                           REG_18_13_port);
   REG_reg_18_12_inst : DLH_X1 port map( G => n52, D => n1820, Q => 
                           REG_18_12_port);
   REG_reg_18_11_inst : DLH_X1 port map( G => n52, D => n1821, Q => 
                           REG_18_11_port);
   REG_reg_18_10_inst : DLH_X1 port map( G => n52, D => n1822, Q => 
                           REG_18_10_port);
   REG_reg_18_9_inst : DLH_X1 port map( G => n52, D => n1823, Q => 
                           REG_18_9_port);
   REG_reg_18_8_inst : DLH_X1 port map( G => n52, D => n1824, Q => 
                           REG_18_8_port);
   REG_reg_18_7_inst : DLH_X1 port map( G => n52, D => n1825, Q => 
                           REG_18_7_port);
   REG_reg_18_6_inst : DLH_X1 port map( G => n52, D => n1826, Q => 
                           REG_18_6_port);
   REG_reg_18_5_inst : DLH_X1 port map( G => n52, D => n1827, Q => 
                           REG_18_5_port);
   REG_reg_18_4_inst : DLH_X1 port map( G => n52, D => n1828, Q => 
                           REG_18_4_port);
   REG_reg_18_3_inst : DLH_X1 port map( G => n52, D => n1829, Q => 
                           REG_18_3_port);
   REG_reg_18_2_inst : DLH_X1 port map( G => n52, D => n1830, Q => 
                           REG_18_2_port);
   REG_reg_18_1_inst : DLH_X1 port map( G => n52, D => n1831, Q => 
                           REG_18_1_port);
   REG_reg_18_0_inst : DLH_X1 port map( G => n52, D => n1832, Q => 
                           REG_18_0_port);
   REG_reg_19_31_inst : DLH_X1 port map( G => n54, D => n1801, Q => 
                           REG_19_31_port);
   REG_reg_19_30_inst : DLH_X1 port map( G => n54, D => n1802, Q => 
                           REG_19_30_port);
   REG_reg_19_29_inst : DLH_X1 port map( G => n54, D => n1803, Q => 
                           REG_19_29_port);
   REG_reg_19_28_inst : DLH_X1 port map( G => n54, D => n1804, Q => 
                           REG_19_28_port);
   REG_reg_19_27_inst : DLH_X1 port map( G => n54, D => n1805, Q => 
                           REG_19_27_port);
   REG_reg_19_26_inst : DLH_X1 port map( G => n54, D => n1806, Q => 
                           REG_19_26_port);
   REG_reg_19_25_inst : DLH_X1 port map( G => n54, D => n1807, Q => 
                           REG_19_25_port);
   REG_reg_19_24_inst : DLH_X1 port map( G => n54, D => n1808, Q => 
                           REG_19_24_port);
   REG_reg_19_23_inst : DLH_X1 port map( G => n54, D => n1809, Q => 
                           REG_19_23_port);
   REG_reg_19_22_inst : DLH_X1 port map( G => n54, D => n1810, Q => 
                           REG_19_22_port);
   REG_reg_19_21_inst : DLH_X1 port map( G => n54, D => n1811, Q => 
                           REG_19_21_port);
   REG_reg_19_20_inst : DLH_X1 port map( G => n54, D => n1812, Q => 
                           REG_19_20_port);
   REG_reg_19_19_inst : DLH_X1 port map( G => n54, D => n1813, Q => 
                           REG_19_19_port);
   REG_reg_19_18_inst : DLH_X1 port map( G => n54, D => n1814, Q => 
                           REG_19_18_port);
   REG_reg_19_17_inst : DLH_X1 port map( G => n54, D => n1815, Q => 
                           REG_19_17_port);
   REG_reg_19_16_inst : DLH_X1 port map( G => n54, D => n1816, Q => 
                           REG_19_16_port);
   REG_reg_19_15_inst : DLH_X1 port map( G => n54, D => n1817, Q => 
                           REG_19_15_port);
   REG_reg_19_14_inst : DLH_X1 port map( G => n54, D => n1818, Q => 
                           REG_19_14_port);
   REG_reg_19_13_inst : DLH_X1 port map( G => n54, D => n1819, Q => 
                           REG_19_13_port);
   REG_reg_19_12_inst : DLH_X1 port map( G => n54, D => n1820, Q => 
                           REG_19_12_port);
   REG_reg_19_11_inst : DLH_X1 port map( G => n54, D => n1821, Q => 
                           REG_19_11_port);
   REG_reg_19_10_inst : DLH_X1 port map( G => n54, D => n1822, Q => 
                           REG_19_10_port);
   REG_reg_19_9_inst : DLH_X1 port map( G => n54, D => n1823, Q => 
                           REG_19_9_port);
   REG_reg_19_8_inst : DLH_X1 port map( G => n54, D => n1824, Q => 
                           REG_19_8_port);
   REG_reg_19_7_inst : DLH_X1 port map( G => n54, D => n1825, Q => 
                           REG_19_7_port);
   REG_reg_19_6_inst : DLH_X1 port map( G => n54, D => n1826, Q => 
                           REG_19_6_port);
   REG_reg_19_5_inst : DLH_X1 port map( G => n54, D => n1827, Q => 
                           REG_19_5_port);
   REG_reg_19_4_inst : DLH_X1 port map( G => n54, D => n1828, Q => 
                           REG_19_4_port);
   REG_reg_19_3_inst : DLH_X1 port map( G => n54, D => n1829, Q => 
                           REG_19_3_port);
   REG_reg_19_2_inst : DLH_X1 port map( G => n54, D => n1830, Q => 
                           REG_19_2_port);
   REG_reg_19_1_inst : DLH_X1 port map( G => n54, D => n1831, Q => 
                           REG_19_1_port);
   REG_reg_19_0_inst : DLH_X1 port map( G => n54, D => n1832, Q => 
                           REG_19_0_port);
   REG_reg_20_31_inst : DLH_X1 port map( G => n56, D => n1801, Q => 
                           REG_20_31_port);
   REG_reg_20_30_inst : DLH_X1 port map( G => n56, D => n1802, Q => 
                           REG_20_30_port);
   REG_reg_20_29_inst : DLH_X1 port map( G => n56, D => n1803, Q => 
                           REG_20_29_port);
   REG_reg_20_28_inst : DLH_X1 port map( G => n56, D => n1804, Q => 
                           REG_20_28_port);
   REG_reg_20_27_inst : DLH_X1 port map( G => n56, D => n1805, Q => 
                           REG_20_27_port);
   REG_reg_20_26_inst : DLH_X1 port map( G => n56, D => n1806, Q => 
                           REG_20_26_port);
   REG_reg_20_25_inst : DLH_X1 port map( G => n56, D => n1807, Q => 
                           REG_20_25_port);
   REG_reg_20_24_inst : DLH_X1 port map( G => n56, D => n1808, Q => 
                           REG_20_24_port);
   REG_reg_20_23_inst : DLH_X1 port map( G => n56, D => n1809, Q => 
                           REG_20_23_port);
   REG_reg_20_22_inst : DLH_X1 port map( G => n56, D => n1810, Q => 
                           REG_20_22_port);
   REG_reg_20_21_inst : DLH_X1 port map( G => n56, D => n1811, Q => 
                           REG_20_21_port);
   REG_reg_20_20_inst : DLH_X1 port map( G => n56, D => n1812, Q => 
                           REG_20_20_port);
   REG_reg_20_19_inst : DLH_X1 port map( G => n56, D => n1813, Q => 
                           REG_20_19_port);
   REG_reg_20_18_inst : DLH_X1 port map( G => n56, D => n1814, Q => 
                           REG_20_18_port);
   REG_reg_20_17_inst : DLH_X1 port map( G => n56, D => n1815, Q => 
                           REG_20_17_port);
   REG_reg_20_16_inst : DLH_X1 port map( G => n56, D => n1816, Q => 
                           REG_20_16_port);
   REG_reg_20_15_inst : DLH_X1 port map( G => n56, D => n1817, Q => 
                           REG_20_15_port);
   REG_reg_20_14_inst : DLH_X1 port map( G => n56, D => n1818, Q => 
                           REG_20_14_port);
   REG_reg_20_13_inst : DLH_X1 port map( G => n56, D => n1819, Q => 
                           REG_20_13_port);
   REG_reg_20_12_inst : DLH_X1 port map( G => n56, D => n1820, Q => 
                           REG_20_12_port);
   REG_reg_20_11_inst : DLH_X1 port map( G => n56, D => n1821, Q => 
                           REG_20_11_port);
   REG_reg_20_10_inst : DLH_X1 port map( G => n56, D => n1822, Q => 
                           REG_20_10_port);
   REG_reg_20_9_inst : DLH_X1 port map( G => n56, D => n1823, Q => 
                           REG_20_9_port);
   REG_reg_20_8_inst : DLH_X1 port map( G => n56, D => n1824, Q => 
                           REG_20_8_port);
   REG_reg_20_7_inst : DLH_X1 port map( G => n56, D => n1825, Q => 
                           REG_20_7_port);
   REG_reg_20_6_inst : DLH_X1 port map( G => n56, D => n1826, Q => 
                           REG_20_6_port);
   REG_reg_20_5_inst : DLH_X1 port map( G => n56, D => n1827, Q => 
                           REG_20_5_port);
   REG_reg_20_4_inst : DLH_X1 port map( G => n56, D => n1828, Q => 
                           REG_20_4_port);
   REG_reg_20_3_inst : DLH_X1 port map( G => n56, D => n1829, Q => 
                           REG_20_3_port);
   REG_reg_20_2_inst : DLH_X1 port map( G => n56, D => n1830, Q => 
                           REG_20_2_port);
   REG_reg_20_1_inst : DLH_X1 port map( G => n56, D => n1831, Q => 
                           REG_20_1_port);
   REG_reg_20_0_inst : DLH_X1 port map( G => n56, D => n1832, Q => 
                           REG_20_0_port);
   REG_reg_21_31_inst : DLH_X1 port map( G => n58, D => n1801, Q => 
                           REG_21_31_port);
   REG_reg_21_30_inst : DLH_X1 port map( G => n58, D => n1802, Q => 
                           REG_21_30_port);
   REG_reg_21_29_inst : DLH_X1 port map( G => n58, D => n1803, Q => 
                           REG_21_29_port);
   REG_reg_21_28_inst : DLH_X1 port map( G => n58, D => n1804, Q => 
                           REG_21_28_port);
   REG_reg_21_27_inst : DLH_X1 port map( G => n58, D => n1805, Q => 
                           REG_21_27_port);
   REG_reg_21_26_inst : DLH_X1 port map( G => n58, D => n1806, Q => 
                           REG_21_26_port);
   REG_reg_21_25_inst : DLH_X1 port map( G => n58, D => n1807, Q => 
                           REG_21_25_port);
   REG_reg_21_24_inst : DLH_X1 port map( G => n58, D => n1808, Q => 
                           REG_21_24_port);
   REG_reg_21_23_inst : DLH_X1 port map( G => n58, D => n1809, Q => 
                           REG_21_23_port);
   REG_reg_21_22_inst : DLH_X1 port map( G => n58, D => n1810, Q => 
                           REG_21_22_port);
   REG_reg_21_21_inst : DLH_X1 port map( G => n58, D => n1811, Q => 
                           REG_21_21_port);
   REG_reg_21_20_inst : DLH_X1 port map( G => n58, D => n1812, Q => 
                           REG_21_20_port);
   REG_reg_21_19_inst : DLH_X1 port map( G => n58, D => n1813, Q => 
                           REG_21_19_port);
   REG_reg_21_18_inst : DLH_X1 port map( G => n58, D => n1814, Q => 
                           REG_21_18_port);
   REG_reg_21_17_inst : DLH_X1 port map( G => n58, D => n1815, Q => 
                           REG_21_17_port);
   REG_reg_21_16_inst : DLH_X1 port map( G => n58, D => n1816, Q => 
                           REG_21_16_port);
   REG_reg_21_15_inst : DLH_X1 port map( G => n58, D => n1817, Q => 
                           REG_21_15_port);
   REG_reg_21_14_inst : DLH_X1 port map( G => n58, D => n1818, Q => 
                           REG_21_14_port);
   REG_reg_21_13_inst : DLH_X1 port map( G => n58, D => n1819, Q => 
                           REG_21_13_port);
   REG_reg_21_12_inst : DLH_X1 port map( G => n58, D => n1820, Q => 
                           REG_21_12_port);
   REG_reg_21_11_inst : DLH_X1 port map( G => n58, D => n1821, Q => 
                           REG_21_11_port);
   REG_reg_21_10_inst : DLH_X1 port map( G => n58, D => n1822, Q => 
                           REG_21_10_port);
   REG_reg_21_9_inst : DLH_X1 port map( G => n58, D => n1823, Q => 
                           REG_21_9_port);
   REG_reg_21_8_inst : DLH_X1 port map( G => n58, D => n1824, Q => 
                           REG_21_8_port);
   REG_reg_21_7_inst : DLH_X1 port map( G => n58, D => n1825, Q => 
                           REG_21_7_port);
   REG_reg_21_6_inst : DLH_X1 port map( G => n58, D => n1826, Q => 
                           REG_21_6_port);
   REG_reg_21_5_inst : DLH_X1 port map( G => n58, D => n1827, Q => 
                           REG_21_5_port);
   REG_reg_21_4_inst : DLH_X1 port map( G => n58, D => n1828, Q => 
                           REG_21_4_port);
   REG_reg_21_3_inst : DLH_X1 port map( G => n58, D => n1829, Q => 
                           REG_21_3_port);
   REG_reg_21_2_inst : DLH_X1 port map( G => n58, D => n1830, Q => 
                           REG_21_2_port);
   REG_reg_21_1_inst : DLH_X1 port map( G => n58, D => n1831, Q => 
                           REG_21_1_port);
   REG_reg_21_0_inst : DLH_X1 port map( G => n58, D => n1832, Q => 
                           REG_21_0_port);
   REG_reg_22_31_inst : DLH_X1 port map( G => n60, D => n1801, Q => 
                           REG_22_31_port);
   REG_reg_22_30_inst : DLH_X1 port map( G => n60, D => n1802, Q => 
                           REG_22_30_port);
   REG_reg_22_29_inst : DLH_X1 port map( G => n60, D => n1803, Q => 
                           REG_22_29_port);
   REG_reg_22_28_inst : DLH_X1 port map( G => n60, D => n1804, Q => 
                           REG_22_28_port);
   REG_reg_22_27_inst : DLH_X1 port map( G => n60, D => n1805, Q => 
                           REG_22_27_port);
   REG_reg_22_26_inst : DLH_X1 port map( G => n60, D => n1806, Q => 
                           REG_22_26_port);
   REG_reg_22_25_inst : DLH_X1 port map( G => n60, D => n1807, Q => 
                           REG_22_25_port);
   REG_reg_22_24_inst : DLH_X1 port map( G => n60, D => n1808, Q => 
                           REG_22_24_port);
   REG_reg_22_23_inst : DLH_X1 port map( G => n60, D => n1809, Q => 
                           REG_22_23_port);
   REG_reg_22_22_inst : DLH_X1 port map( G => n60, D => n1810, Q => 
                           REG_22_22_port);
   REG_reg_22_21_inst : DLH_X1 port map( G => n60, D => n1811, Q => 
                           REG_22_21_port);
   REG_reg_22_20_inst : DLH_X1 port map( G => n60, D => n1812, Q => 
                           REG_22_20_port);
   REG_reg_22_19_inst : DLH_X1 port map( G => n60, D => n1813, Q => 
                           REG_22_19_port);
   REG_reg_22_18_inst : DLH_X1 port map( G => n60, D => n1814, Q => 
                           REG_22_18_port);
   REG_reg_22_17_inst : DLH_X1 port map( G => n60, D => n1815, Q => 
                           REG_22_17_port);
   REG_reg_22_16_inst : DLH_X1 port map( G => n60, D => n1816, Q => 
                           REG_22_16_port);
   REG_reg_22_15_inst : DLH_X1 port map( G => n60, D => n1817, Q => 
                           REG_22_15_port);
   REG_reg_22_14_inst : DLH_X1 port map( G => n60, D => n1818, Q => 
                           REG_22_14_port);
   REG_reg_22_13_inst : DLH_X1 port map( G => n60, D => n1819, Q => 
                           REG_22_13_port);
   REG_reg_22_12_inst : DLH_X1 port map( G => n60, D => n1820, Q => 
                           REG_22_12_port);
   REG_reg_22_11_inst : DLH_X1 port map( G => n60, D => n1821, Q => 
                           REG_22_11_port);
   REG_reg_22_10_inst : DLH_X1 port map( G => n60, D => n1822, Q => 
                           REG_22_10_port);
   REG_reg_22_9_inst : DLH_X1 port map( G => n60, D => n1823, Q => 
                           REG_22_9_port);
   REG_reg_22_8_inst : DLH_X1 port map( G => n60, D => n1824, Q => 
                           REG_22_8_port);
   REG_reg_22_7_inst : DLH_X1 port map( G => n60, D => n1825, Q => 
                           REG_22_7_port);
   REG_reg_22_6_inst : DLH_X1 port map( G => n60, D => n1826, Q => 
                           REG_22_6_port);
   REG_reg_22_5_inst : DLH_X1 port map( G => n60, D => n1827, Q => 
                           REG_22_5_port);
   REG_reg_22_4_inst : DLH_X1 port map( G => n60, D => n1828, Q => 
                           REG_22_4_port);
   REG_reg_22_3_inst : DLH_X1 port map( G => n60, D => n1829, Q => 
                           REG_22_3_port);
   REG_reg_22_2_inst : DLH_X1 port map( G => n60, D => n1830, Q => 
                           REG_22_2_port);
   REG_reg_22_1_inst : DLH_X1 port map( G => n60, D => n1831, Q => 
                           REG_22_1_port);
   REG_reg_22_0_inst : DLH_X1 port map( G => n60, D => n1832, Q => 
                           REG_22_0_port);
   REG_reg_23_31_inst : DLH_X1 port map( G => n62, D => n1801, Q => 
                           REG_23_31_port);
   REG_reg_23_30_inst : DLH_X1 port map( G => n62, D => n1802, Q => 
                           REG_23_30_port);
   REG_reg_23_29_inst : DLH_X1 port map( G => n62, D => n1803, Q => 
                           REG_23_29_port);
   REG_reg_23_28_inst : DLH_X1 port map( G => n62, D => n1804, Q => 
                           REG_23_28_port);
   REG_reg_23_27_inst : DLH_X1 port map( G => n62, D => n1805, Q => 
                           REG_23_27_port);
   REG_reg_23_26_inst : DLH_X1 port map( G => n62, D => n1806, Q => 
                           REG_23_26_port);
   REG_reg_23_25_inst : DLH_X1 port map( G => n62, D => n1807, Q => 
                           REG_23_25_port);
   REG_reg_23_24_inst : DLH_X1 port map( G => n62, D => n1808, Q => 
                           REG_23_24_port);
   REG_reg_23_23_inst : DLH_X1 port map( G => n62, D => n1809, Q => 
                           REG_23_23_port);
   REG_reg_23_22_inst : DLH_X1 port map( G => n62, D => n1810, Q => 
                           REG_23_22_port);
   REG_reg_23_21_inst : DLH_X1 port map( G => n62, D => n1811, Q => 
                           REG_23_21_port);
   REG_reg_23_20_inst : DLH_X1 port map( G => n62, D => n1812, Q => 
                           REG_23_20_port);
   REG_reg_23_19_inst : DLH_X1 port map( G => n62, D => n1813, Q => 
                           REG_23_19_port);
   REG_reg_23_18_inst : DLH_X1 port map( G => n62, D => n1814, Q => 
                           REG_23_18_port);
   REG_reg_23_17_inst : DLH_X1 port map( G => n62, D => n1815, Q => 
                           REG_23_17_port);
   REG_reg_23_16_inst : DLH_X1 port map( G => n62, D => n1816, Q => 
                           REG_23_16_port);
   REG_reg_23_15_inst : DLH_X1 port map( G => n62, D => n1817, Q => 
                           REG_23_15_port);
   REG_reg_23_14_inst : DLH_X1 port map( G => n62, D => n1818, Q => 
                           REG_23_14_port);
   REG_reg_23_13_inst : DLH_X1 port map( G => n62, D => n1819, Q => 
                           REG_23_13_port);
   REG_reg_23_12_inst : DLH_X1 port map( G => n62, D => n1820, Q => 
                           REG_23_12_port);
   REG_reg_23_11_inst : DLH_X1 port map( G => n62, D => n1821, Q => 
                           REG_23_11_port);
   REG_reg_23_10_inst : DLH_X1 port map( G => n62, D => n1822, Q => 
                           REG_23_10_port);
   REG_reg_23_9_inst : DLH_X1 port map( G => n62, D => n1823, Q => 
                           REG_23_9_port);
   REG_reg_23_8_inst : DLH_X1 port map( G => n62, D => n1824, Q => 
                           REG_23_8_port);
   REG_reg_23_7_inst : DLH_X1 port map( G => n62, D => n1825, Q => 
                           REG_23_7_port);
   REG_reg_23_6_inst : DLH_X1 port map( G => n62, D => n1826, Q => 
                           REG_23_6_port);
   REG_reg_23_5_inst : DLH_X1 port map( G => n62, D => n1827, Q => 
                           REG_23_5_port);
   REG_reg_23_4_inst : DLH_X1 port map( G => n62, D => n1828, Q => 
                           REG_23_4_port);
   REG_reg_23_3_inst : DLH_X1 port map( G => n62, D => n1829, Q => 
                           REG_23_3_port);
   REG_reg_23_2_inst : DLH_X1 port map( G => n62, D => n1830, Q => 
                           REG_23_2_port);
   REG_reg_23_1_inst : DLH_X1 port map( G => n62, D => n1831, Q => 
                           REG_23_1_port);
   REG_reg_23_0_inst : DLH_X1 port map( G => n62, D => n1832, Q => 
                           REG_23_0_port);
   REG_reg_24_31_inst : DLH_X1 port map( G => n64, D => n1801, Q => 
                           REG_24_31_port);
   REG_reg_24_30_inst : DLH_X1 port map( G => n64, D => n1802, Q => 
                           REG_24_30_port);
   REG_reg_24_29_inst : DLH_X1 port map( G => n64, D => n1803, Q => 
                           REG_24_29_port);
   REG_reg_24_28_inst : DLH_X1 port map( G => n64, D => n1804, Q => 
                           REG_24_28_port);
   REG_reg_24_27_inst : DLH_X1 port map( G => n64, D => n1805, Q => 
                           REG_24_27_port);
   REG_reg_24_26_inst : DLH_X1 port map( G => n64, D => n1806, Q => 
                           REG_24_26_port);
   REG_reg_24_25_inst : DLH_X1 port map( G => n64, D => n1807, Q => 
                           REG_24_25_port);
   REG_reg_24_24_inst : DLH_X1 port map( G => n64, D => n1808, Q => 
                           REG_24_24_port);
   REG_reg_24_23_inst : DLH_X1 port map( G => n64, D => n1809, Q => 
                           REG_24_23_port);
   REG_reg_24_22_inst : DLH_X1 port map( G => n64, D => n1810, Q => 
                           REG_24_22_port);
   REG_reg_24_21_inst : DLH_X1 port map( G => n64, D => n1811, Q => 
                           REG_24_21_port);
   REG_reg_24_20_inst : DLH_X1 port map( G => n64, D => n1812, Q => 
                           REG_24_20_port);
   REG_reg_24_19_inst : DLH_X1 port map( G => n64, D => n1813, Q => 
                           REG_24_19_port);
   REG_reg_24_18_inst : DLH_X1 port map( G => n64, D => n1814, Q => 
                           REG_24_18_port);
   REG_reg_24_17_inst : DLH_X1 port map( G => n64, D => n1815, Q => 
                           REG_24_17_port);
   REG_reg_24_16_inst : DLH_X1 port map( G => n64, D => n1816, Q => 
                           REG_24_16_port);
   REG_reg_24_15_inst : DLH_X1 port map( G => n64, D => n1817, Q => 
                           REG_24_15_port);
   REG_reg_24_14_inst : DLH_X1 port map( G => n64, D => n1818, Q => 
                           REG_24_14_port);
   REG_reg_24_13_inst : DLH_X1 port map( G => n64, D => n1819, Q => 
                           REG_24_13_port);
   REG_reg_24_12_inst : DLH_X1 port map( G => n64, D => n1820, Q => 
                           REG_24_12_port);
   REG_reg_24_11_inst : DLH_X1 port map( G => n64, D => n1821, Q => 
                           REG_24_11_port);
   REG_reg_24_10_inst : DLH_X1 port map( G => n64, D => n1822, Q => 
                           REG_24_10_port);
   REG_reg_24_9_inst : DLH_X1 port map( G => n64, D => n1823, Q => 
                           REG_24_9_port);
   REG_reg_24_8_inst : DLH_X1 port map( G => n64, D => n1824, Q => 
                           REG_24_8_port);
   REG_reg_24_7_inst : DLH_X1 port map( G => n64, D => n1825, Q => 
                           REG_24_7_port);
   REG_reg_24_6_inst : DLH_X1 port map( G => n64, D => n1826, Q => 
                           REG_24_6_port);
   REG_reg_24_5_inst : DLH_X1 port map( G => n64, D => n1827, Q => 
                           REG_24_5_port);
   REG_reg_24_4_inst : DLH_X1 port map( G => n64, D => n1828, Q => 
                           REG_24_4_port);
   REG_reg_24_3_inst : DLH_X1 port map( G => n64, D => n1829, Q => 
                           REG_24_3_port);
   REG_reg_24_2_inst : DLH_X1 port map( G => n64, D => n1830, Q => 
                           REG_24_2_port);
   REG_reg_24_1_inst : DLH_X1 port map( G => n64, D => n1831, Q => 
                           REG_24_1_port);
   REG_reg_24_0_inst : DLH_X1 port map( G => n64, D => n1832, Q => 
                           REG_24_0_port);
   REG_reg_25_31_inst : DLH_X1 port map( G => n66, D => n1801, Q => 
                           REG_25_31_port);
   REG_reg_25_30_inst : DLH_X1 port map( G => n66, D => n1802, Q => 
                           REG_25_30_port);
   REG_reg_25_29_inst : DLH_X1 port map( G => n66, D => n1803, Q => 
                           REG_25_29_port);
   REG_reg_25_28_inst : DLH_X1 port map( G => n66, D => n1804, Q => 
                           REG_25_28_port);
   REG_reg_25_27_inst : DLH_X1 port map( G => n66, D => n1805, Q => 
                           REG_25_27_port);
   REG_reg_25_26_inst : DLH_X1 port map( G => n66, D => n1806, Q => 
                           REG_25_26_port);
   REG_reg_25_25_inst : DLH_X1 port map( G => n66, D => n1807, Q => 
                           REG_25_25_port);
   REG_reg_25_24_inst : DLH_X1 port map( G => n66, D => n1808, Q => 
                           REG_25_24_port);
   REG_reg_25_23_inst : DLH_X1 port map( G => n66, D => n1809, Q => 
                           REG_25_23_port);
   REG_reg_25_22_inst : DLH_X1 port map( G => n66, D => n1810, Q => 
                           REG_25_22_port);
   REG_reg_25_21_inst : DLH_X1 port map( G => n66, D => n1811, Q => 
                           REG_25_21_port);
   REG_reg_25_20_inst : DLH_X1 port map( G => n66, D => n1812, Q => 
                           REG_25_20_port);
   REG_reg_25_19_inst : DLH_X1 port map( G => n66, D => n1813, Q => 
                           REG_25_19_port);
   REG_reg_25_18_inst : DLH_X1 port map( G => n66, D => n1814, Q => 
                           REG_25_18_port);
   REG_reg_25_17_inst : DLH_X1 port map( G => n66, D => n1815, Q => 
                           REG_25_17_port);
   REG_reg_25_16_inst : DLH_X1 port map( G => n66, D => n1816, Q => 
                           REG_25_16_port);
   REG_reg_25_15_inst : DLH_X1 port map( G => n66, D => n1817, Q => 
                           REG_25_15_port);
   REG_reg_25_14_inst : DLH_X1 port map( G => n66, D => n1818, Q => 
                           REG_25_14_port);
   REG_reg_25_13_inst : DLH_X1 port map( G => n66, D => n1819, Q => 
                           REG_25_13_port);
   REG_reg_25_12_inst : DLH_X1 port map( G => n66, D => n1820, Q => 
                           REG_25_12_port);
   REG_reg_25_11_inst : DLH_X1 port map( G => n66, D => n1821, Q => 
                           REG_25_11_port);
   REG_reg_25_10_inst : DLH_X1 port map( G => n66, D => n1822, Q => 
                           REG_25_10_port);
   REG_reg_25_9_inst : DLH_X1 port map( G => n66, D => n1823, Q => 
                           REG_25_9_port);
   REG_reg_25_8_inst : DLH_X1 port map( G => n66, D => n1824, Q => 
                           REG_25_8_port);
   REG_reg_25_7_inst : DLH_X1 port map( G => n66, D => n1825, Q => 
                           REG_25_7_port);
   REG_reg_25_6_inst : DLH_X1 port map( G => n66, D => n1826, Q => 
                           REG_25_6_port);
   REG_reg_25_5_inst : DLH_X1 port map( G => n66, D => n1827, Q => 
                           REG_25_5_port);
   REG_reg_25_4_inst : DLH_X1 port map( G => n66, D => n1828, Q => 
                           REG_25_4_port);
   REG_reg_25_3_inst : DLH_X1 port map( G => n66, D => n1829, Q => 
                           REG_25_3_port);
   REG_reg_25_2_inst : DLH_X1 port map( G => n66, D => n1830, Q => 
                           REG_25_2_port);
   REG_reg_25_1_inst : DLH_X1 port map( G => n66, D => n1831, Q => 
                           REG_25_1_port);
   REG_reg_25_0_inst : DLH_X1 port map( G => n66, D => n1832, Q => 
                           REG_25_0_port);
   REG_reg_26_31_inst : DLH_X1 port map( G => n68, D => n1801, Q => 
                           REG_26_31_port);
   REG_reg_26_30_inst : DLH_X1 port map( G => n68, D => n1802, Q => 
                           REG_26_30_port);
   REG_reg_26_29_inst : DLH_X1 port map( G => n68, D => n1803, Q => 
                           REG_26_29_port);
   REG_reg_26_28_inst : DLH_X1 port map( G => n68, D => n1804, Q => 
                           REG_26_28_port);
   REG_reg_26_27_inst : DLH_X1 port map( G => n68, D => n1805, Q => 
                           REG_26_27_port);
   REG_reg_26_26_inst : DLH_X1 port map( G => n68, D => n1806, Q => 
                           REG_26_26_port);
   REG_reg_26_25_inst : DLH_X1 port map( G => n68, D => n1807, Q => 
                           REG_26_25_port);
   REG_reg_26_24_inst : DLH_X1 port map( G => n68, D => n1808, Q => 
                           REG_26_24_port);
   REG_reg_26_23_inst : DLH_X1 port map( G => n68, D => n1809, Q => 
                           REG_26_23_port);
   REG_reg_26_22_inst : DLH_X1 port map( G => n68, D => n1810, Q => 
                           REG_26_22_port);
   REG_reg_26_21_inst : DLH_X1 port map( G => n68, D => n1811, Q => 
                           REG_26_21_port);
   REG_reg_26_20_inst : DLH_X1 port map( G => n68, D => n1812, Q => 
                           REG_26_20_port);
   REG_reg_26_19_inst : DLH_X1 port map( G => n68, D => n1813, Q => 
                           REG_26_19_port);
   REG_reg_26_18_inst : DLH_X1 port map( G => n68, D => n1814, Q => 
                           REG_26_18_port);
   REG_reg_26_17_inst : DLH_X1 port map( G => n68, D => n1815, Q => 
                           REG_26_17_port);
   REG_reg_26_16_inst : DLH_X1 port map( G => n68, D => n1816, Q => 
                           REG_26_16_port);
   REG_reg_26_15_inst : DLH_X1 port map( G => n68, D => n1817, Q => 
                           REG_26_15_port);
   REG_reg_26_14_inst : DLH_X1 port map( G => n68, D => n1818, Q => 
                           REG_26_14_port);
   REG_reg_26_13_inst : DLH_X1 port map( G => n68, D => n1819, Q => 
                           REG_26_13_port);
   REG_reg_26_12_inst : DLH_X1 port map( G => n68, D => n1820, Q => 
                           REG_26_12_port);
   REG_reg_26_11_inst : DLH_X1 port map( G => n68, D => n1821, Q => 
                           REG_26_11_port);
   REG_reg_26_10_inst : DLH_X1 port map( G => n68, D => n1822, Q => 
                           REG_26_10_port);
   REG_reg_26_9_inst : DLH_X1 port map( G => n68, D => n1823, Q => 
                           REG_26_9_port);
   REG_reg_26_8_inst : DLH_X1 port map( G => n68, D => n1824, Q => 
                           REG_26_8_port);
   REG_reg_26_7_inst : DLH_X1 port map( G => n68, D => n1825, Q => 
                           REG_26_7_port);
   REG_reg_26_6_inst : DLH_X1 port map( G => n68, D => n1826, Q => 
                           REG_26_6_port);
   REG_reg_26_5_inst : DLH_X1 port map( G => n68, D => n1827, Q => 
                           REG_26_5_port);
   REG_reg_26_4_inst : DLH_X1 port map( G => n68, D => n1828, Q => 
                           REG_26_4_port);
   REG_reg_26_3_inst : DLH_X1 port map( G => n68, D => n1829, Q => 
                           REG_26_3_port);
   REG_reg_26_2_inst : DLH_X1 port map( G => n68, D => n1830, Q => 
                           REG_26_2_port);
   REG_reg_26_1_inst : DLH_X1 port map( G => n68, D => n1831, Q => 
                           REG_26_1_port);
   REG_reg_26_0_inst : DLH_X1 port map( G => n68, D => n1832, Q => 
                           REG_26_0_port);
   REG_reg_27_31_inst : DLH_X1 port map( G => n70, D => n1801, Q => 
                           REG_27_31_port);
   REG_reg_27_30_inst : DLH_X1 port map( G => n70, D => n1802, Q => 
                           REG_27_30_port);
   REG_reg_27_29_inst : DLH_X1 port map( G => n70, D => n1803, Q => 
                           REG_27_29_port);
   REG_reg_27_28_inst : DLH_X1 port map( G => n70, D => n1804, Q => 
                           REG_27_28_port);
   REG_reg_27_27_inst : DLH_X1 port map( G => n70, D => n1805, Q => 
                           REG_27_27_port);
   REG_reg_27_26_inst : DLH_X1 port map( G => n70, D => n1806, Q => 
                           REG_27_26_port);
   REG_reg_27_25_inst : DLH_X1 port map( G => n70, D => n1807, Q => 
                           REG_27_25_port);
   REG_reg_27_24_inst : DLH_X1 port map( G => n70, D => n1808, Q => 
                           REG_27_24_port);
   REG_reg_27_23_inst : DLH_X1 port map( G => n70, D => n1809, Q => 
                           REG_27_23_port);
   REG_reg_27_22_inst : DLH_X1 port map( G => n70, D => n1810, Q => 
                           REG_27_22_port);
   REG_reg_27_21_inst : DLH_X1 port map( G => n70, D => n1811, Q => 
                           REG_27_21_port);
   REG_reg_27_20_inst : DLH_X1 port map( G => n70, D => n1812, Q => 
                           REG_27_20_port);
   REG_reg_27_19_inst : DLH_X1 port map( G => n70, D => n1813, Q => 
                           REG_27_19_port);
   REG_reg_27_18_inst : DLH_X1 port map( G => n70, D => n1814, Q => 
                           REG_27_18_port);
   REG_reg_27_17_inst : DLH_X1 port map( G => n70, D => n1815, Q => 
                           REG_27_17_port);
   REG_reg_27_16_inst : DLH_X1 port map( G => n70, D => n1816, Q => 
                           REG_27_16_port);
   REG_reg_27_15_inst : DLH_X1 port map( G => n70, D => n1817, Q => 
                           REG_27_15_port);
   REG_reg_27_14_inst : DLH_X1 port map( G => n70, D => n1818, Q => 
                           REG_27_14_port);
   REG_reg_27_13_inst : DLH_X1 port map( G => n70, D => n1819, Q => 
                           REG_27_13_port);
   REG_reg_27_12_inst : DLH_X1 port map( G => n70, D => n1820, Q => 
                           REG_27_12_port);
   REG_reg_27_11_inst : DLH_X1 port map( G => n70, D => n1821, Q => 
                           REG_27_11_port);
   REG_reg_27_10_inst : DLH_X1 port map( G => n70, D => n1822, Q => 
                           REG_27_10_port);
   REG_reg_27_9_inst : DLH_X1 port map( G => n70, D => n1823, Q => 
                           REG_27_9_port);
   REG_reg_27_8_inst : DLH_X1 port map( G => n70, D => n1824, Q => 
                           REG_27_8_port);
   REG_reg_27_7_inst : DLH_X1 port map( G => n70, D => n1825, Q => 
                           REG_27_7_port);
   REG_reg_27_6_inst : DLH_X1 port map( G => n70, D => n1826, Q => 
                           REG_27_6_port);
   REG_reg_27_5_inst : DLH_X1 port map( G => n70, D => n1827, Q => 
                           REG_27_5_port);
   REG_reg_27_4_inst : DLH_X1 port map( G => n70, D => n1828, Q => 
                           REG_27_4_port);
   REG_reg_27_3_inst : DLH_X1 port map( G => n70, D => n1829, Q => 
                           REG_27_3_port);
   REG_reg_27_2_inst : DLH_X1 port map( G => n70, D => n1830, Q => 
                           REG_27_2_port);
   REG_reg_27_1_inst : DLH_X1 port map( G => n70, D => n1831, Q => 
                           REG_27_1_port);
   REG_reg_27_0_inst : DLH_X1 port map( G => n70, D => n1832, Q => 
                           REG_27_0_port);
   REG_reg_28_31_inst : DLH_X1 port map( G => n72, D => n1801, Q => 
                           REG_28_31_port);
   REG_reg_28_30_inst : DLH_X1 port map( G => n72, D => n1802, Q => 
                           REG_28_30_port);
   REG_reg_28_29_inst : DLH_X1 port map( G => n72, D => n1803, Q => 
                           REG_28_29_port);
   REG_reg_28_28_inst : DLH_X1 port map( G => n72, D => n1804, Q => 
                           REG_28_28_port);
   REG_reg_28_27_inst : DLH_X1 port map( G => n72, D => n1805, Q => 
                           REG_28_27_port);
   REG_reg_28_26_inst : DLH_X1 port map( G => n72, D => n1806, Q => 
                           REG_28_26_port);
   REG_reg_28_25_inst : DLH_X1 port map( G => n72, D => n1807, Q => 
                           REG_28_25_port);
   REG_reg_28_24_inst : DLH_X1 port map( G => n72, D => n1808, Q => 
                           REG_28_24_port);
   REG_reg_28_23_inst : DLH_X1 port map( G => n72, D => n1809, Q => 
                           REG_28_23_port);
   REG_reg_28_22_inst : DLH_X1 port map( G => n72, D => n1810, Q => 
                           REG_28_22_port);
   REG_reg_28_21_inst : DLH_X1 port map( G => n72, D => n1811, Q => 
                           REG_28_21_port);
   REG_reg_28_20_inst : DLH_X1 port map( G => n72, D => n1812, Q => 
                           REG_28_20_port);
   REG_reg_28_19_inst : DLH_X1 port map( G => n72, D => n1813, Q => 
                           REG_28_19_port);
   REG_reg_28_18_inst : DLH_X1 port map( G => n72, D => n1814, Q => 
                           REG_28_18_port);
   REG_reg_28_17_inst : DLH_X1 port map( G => n72, D => n1815, Q => 
                           REG_28_17_port);
   REG_reg_28_16_inst : DLH_X1 port map( G => n72, D => n1816, Q => 
                           REG_28_16_port);
   REG_reg_28_15_inst : DLH_X1 port map( G => n72, D => n1817, Q => 
                           REG_28_15_port);
   REG_reg_28_14_inst : DLH_X1 port map( G => n72, D => n1818, Q => 
                           REG_28_14_port);
   REG_reg_28_13_inst : DLH_X1 port map( G => n72, D => n1819, Q => 
                           REG_28_13_port);
   REG_reg_28_12_inst : DLH_X1 port map( G => n72, D => n1820, Q => 
                           REG_28_12_port);
   REG_reg_28_11_inst : DLH_X1 port map( G => n72, D => n1821, Q => 
                           REG_28_11_port);
   REG_reg_28_10_inst : DLH_X1 port map( G => n72, D => n1822, Q => 
                           REG_28_10_port);
   REG_reg_28_9_inst : DLH_X1 port map( G => n72, D => n1823, Q => 
                           REG_28_9_port);
   REG_reg_28_8_inst : DLH_X1 port map( G => n72, D => n1824, Q => 
                           REG_28_8_port);
   REG_reg_28_7_inst : DLH_X1 port map( G => n72, D => n1825, Q => 
                           REG_28_7_port);
   REG_reg_28_6_inst : DLH_X1 port map( G => n72, D => n1826, Q => 
                           REG_28_6_port);
   REG_reg_28_5_inst : DLH_X1 port map( G => n72, D => n1827, Q => 
                           REG_28_5_port);
   REG_reg_28_4_inst : DLH_X1 port map( G => n72, D => n1828, Q => 
                           REG_28_4_port);
   REG_reg_28_3_inst : DLH_X1 port map( G => n72, D => n1829, Q => 
                           REG_28_3_port);
   REG_reg_28_2_inst : DLH_X1 port map( G => n72, D => n1830, Q => 
                           REG_28_2_port);
   REG_reg_28_1_inst : DLH_X1 port map( G => n72, D => n1831, Q => 
                           REG_28_1_port);
   REG_reg_28_0_inst : DLH_X1 port map( G => n72, D => n1832, Q => 
                           REG_28_0_port);
   REG_reg_29_31_inst : DLH_X1 port map( G => n78, D => n1801, Q => 
                           REG_29_31_port);
   REG_reg_29_30_inst : DLH_X1 port map( G => n78, D => n1802, Q => 
                           REG_29_30_port);
   REG_reg_29_29_inst : DLH_X1 port map( G => n78, D => n1803, Q => 
                           REG_29_29_port);
   REG_reg_29_28_inst : DLH_X1 port map( G => n78, D => n1804, Q => 
                           REG_29_28_port);
   REG_reg_29_27_inst : DLH_X1 port map( G => n78, D => n1805, Q => 
                           REG_29_27_port);
   REG_reg_29_26_inst : DLH_X1 port map( G => n78, D => n1806, Q => 
                           REG_29_26_port);
   REG_reg_29_25_inst : DLH_X1 port map( G => n78, D => n1807, Q => 
                           REG_29_25_port);
   REG_reg_29_24_inst : DLH_X1 port map( G => n78, D => n1808, Q => 
                           REG_29_24_port);
   REG_reg_29_23_inst : DLH_X1 port map( G => n78, D => n1809, Q => 
                           REG_29_23_port);
   REG_reg_29_22_inst : DLH_X1 port map( G => n78, D => n1810, Q => 
                           REG_29_22_port);
   REG_reg_29_21_inst : DLH_X1 port map( G => n78, D => n1811, Q => 
                           REG_29_21_port);
   REG_reg_29_20_inst : DLH_X1 port map( G => n78, D => n1812, Q => 
                           REG_29_20_port);
   REG_reg_29_19_inst : DLH_X1 port map( G => n78, D => n1813, Q => 
                           REG_29_19_port);
   REG_reg_29_18_inst : DLH_X1 port map( G => n78, D => n1814, Q => 
                           REG_29_18_port);
   REG_reg_29_17_inst : DLH_X1 port map( G => n78, D => n1815, Q => 
                           REG_29_17_port);
   REG_reg_29_16_inst : DLH_X1 port map( G => n78, D => n1816, Q => 
                           REG_29_16_port);
   REG_reg_29_15_inst : DLH_X1 port map( G => n78, D => n1817, Q => 
                           REG_29_15_port);
   REG_reg_29_14_inst : DLH_X1 port map( G => n78, D => n1818, Q => 
                           REG_29_14_port);
   REG_reg_29_13_inst : DLH_X1 port map( G => n78, D => n1819, Q => 
                           REG_29_13_port);
   REG_reg_29_12_inst : DLH_X1 port map( G => n78, D => n1820, Q => 
                           REG_29_12_port);
   REG_reg_29_11_inst : DLH_X1 port map( G => n78, D => n1821, Q => 
                           REG_29_11_port);
   REG_reg_29_10_inst : DLH_X1 port map( G => n78, D => n1822, Q => 
                           REG_29_10_port);
   REG_reg_29_9_inst : DLH_X1 port map( G => n78, D => n1823, Q => 
                           REG_29_9_port);
   REG_reg_29_8_inst : DLH_X1 port map( G => n78, D => n1824, Q => 
                           REG_29_8_port);
   REG_reg_29_7_inst : DLH_X1 port map( G => n78, D => n1825, Q => 
                           REG_29_7_port);
   REG_reg_29_6_inst : DLH_X1 port map( G => n78, D => n1826, Q => 
                           REG_29_6_port);
   REG_reg_29_5_inst : DLH_X1 port map( G => n78, D => n1827, Q => 
                           REG_29_5_port);
   REG_reg_29_4_inst : DLH_X1 port map( G => n78, D => n1828, Q => 
                           REG_29_4_port);
   REG_reg_29_3_inst : DLH_X1 port map( G => n78, D => n1829, Q => 
                           REG_29_3_port);
   REG_reg_29_2_inst : DLH_X1 port map( G => n78, D => n1830, Q => 
                           REG_29_2_port);
   REG_reg_29_1_inst : DLH_X1 port map( G => n78, D => n1831, Q => 
                           REG_29_1_port);
   REG_reg_29_0_inst : DLH_X1 port map( G => n78, D => n1832, Q => 
                           REG_29_0_port);
   REG_reg_30_31_inst : DLH_X1 port map( G => n80, D => n1801, Q => 
                           REG_30_31_port);
   REG_reg_30_30_inst : DLH_X1 port map( G => n80, D => n1802, Q => 
                           REG_30_30_port);
   REG_reg_30_29_inst : DLH_X1 port map( G => n80, D => n1803, Q => 
                           REG_30_29_port);
   REG_reg_30_28_inst : DLH_X1 port map( G => n80, D => n1804, Q => 
                           REG_30_28_port);
   REG_reg_30_27_inst : DLH_X1 port map( G => n80, D => n1805, Q => 
                           REG_30_27_port);
   REG_reg_30_26_inst : DLH_X1 port map( G => n80, D => n1806, Q => 
                           REG_30_26_port);
   REG_reg_30_25_inst : DLH_X1 port map( G => n80, D => n1807, Q => 
                           REG_30_25_port);
   REG_reg_30_24_inst : DLH_X1 port map( G => n80, D => n1808, Q => 
                           REG_30_24_port);
   REG_reg_30_23_inst : DLH_X1 port map( G => n80, D => n1809, Q => 
                           REG_30_23_port);
   REG_reg_30_22_inst : DLH_X1 port map( G => n80, D => n1810, Q => 
                           REG_30_22_port);
   REG_reg_30_21_inst : DLH_X1 port map( G => n80, D => n1811, Q => 
                           REG_30_21_port);
   REG_reg_30_20_inst : DLH_X1 port map( G => n80, D => n1812, Q => 
                           REG_30_20_port);
   REG_reg_30_19_inst : DLH_X1 port map( G => n80, D => n1813, Q => 
                           REG_30_19_port);
   REG_reg_30_18_inst : DLH_X1 port map( G => n80, D => n1814, Q => 
                           REG_30_18_port);
   REG_reg_30_17_inst : DLH_X1 port map( G => n80, D => n1815, Q => 
                           REG_30_17_port);
   REG_reg_30_16_inst : DLH_X1 port map( G => n80, D => n1816, Q => 
                           REG_30_16_port);
   REG_reg_30_15_inst : DLH_X1 port map( G => n80, D => n1817, Q => 
                           REG_30_15_port);
   REG_reg_30_14_inst : DLH_X1 port map( G => n80, D => n1818, Q => 
                           REG_30_14_port);
   REG_reg_30_13_inst : DLH_X1 port map( G => n80, D => n1819, Q => 
                           REG_30_13_port);
   REG_reg_30_12_inst : DLH_X1 port map( G => n80, D => n1820, Q => 
                           REG_30_12_port);
   REG_reg_30_11_inst : DLH_X1 port map( G => n80, D => n1821, Q => 
                           REG_30_11_port);
   REG_reg_30_10_inst : DLH_X1 port map( G => n80, D => n1822, Q => 
                           REG_30_10_port);
   REG_reg_30_9_inst : DLH_X1 port map( G => n80, D => n1823, Q => 
                           REG_30_9_port);
   REG_reg_30_8_inst : DLH_X1 port map( G => n80, D => n1824, Q => 
                           REG_30_8_port);
   REG_reg_30_7_inst : DLH_X1 port map( G => n80, D => n1825, Q => 
                           REG_30_7_port);
   REG_reg_30_6_inst : DLH_X1 port map( G => n80, D => n1826, Q => 
                           REG_30_6_port);
   REG_reg_30_5_inst : DLH_X1 port map( G => n80, D => n1827, Q => 
                           REG_30_5_port);
   REG_reg_30_4_inst : DLH_X1 port map( G => n80, D => n1828, Q => 
                           REG_30_4_port);
   REG_reg_30_3_inst : DLH_X1 port map( G => n80, D => n1829, Q => 
                           REG_30_3_port);
   REG_reg_30_2_inst : DLH_X1 port map( G => n80, D => n1830, Q => 
                           REG_30_2_port);
   REG_reg_30_1_inst : DLH_X1 port map( G => n80, D => n1831, Q => 
                           REG_30_1_port);
   REG_reg_30_0_inst : DLH_X1 port map( G => n80, D => n1832, Q => 
                           REG_30_0_port);
   REG_reg_31_31_inst : DLH_X1 port map( G => n82, D => n1801, Q => 
                           REG_31_31_port);
   REG_reg_31_30_inst : DLH_X1 port map( G => n82, D => n1802, Q => 
                           REG_31_30_port);
   REG_reg_31_29_inst : DLH_X1 port map( G => n82, D => n1803, Q => 
                           REG_31_29_port);
   REG_reg_31_28_inst : DLH_X1 port map( G => n82, D => n1804, Q => 
                           REG_31_28_port);
   REG_reg_31_27_inst : DLH_X1 port map( G => n82, D => n1805, Q => 
                           REG_31_27_port);
   REG_reg_31_26_inst : DLH_X1 port map( G => n82, D => n1806, Q => 
                           REG_31_26_port);
   REG_reg_31_25_inst : DLH_X1 port map( G => n82, D => n1807, Q => 
                           REG_31_25_port);
   REG_reg_31_24_inst : DLH_X1 port map( G => n82, D => n1808, Q => 
                           REG_31_24_port);
   REG_reg_31_23_inst : DLH_X1 port map( G => n82, D => n1809, Q => 
                           REG_31_23_port);
   REG_reg_31_22_inst : DLH_X1 port map( G => n82, D => n1810, Q => 
                           REG_31_22_port);
   REG_reg_31_21_inst : DLH_X1 port map( G => n82, D => n1811, Q => 
                           REG_31_21_port);
   REG_reg_31_20_inst : DLH_X1 port map( G => n82, D => n1812, Q => 
                           REG_31_20_port);
   REG_reg_31_19_inst : DLH_X1 port map( G => n82, D => n1813, Q => 
                           REG_31_19_port);
   REG_reg_31_18_inst : DLH_X1 port map( G => n82, D => n1814, Q => 
                           REG_31_18_port);
   REG_reg_31_17_inst : DLH_X1 port map( G => n82, D => n1815, Q => 
                           REG_31_17_port);
   REG_reg_31_16_inst : DLH_X1 port map( G => n82, D => n1816, Q => 
                           REG_31_16_port);
   REG_reg_31_15_inst : DLH_X1 port map( G => n82, D => n1817, Q => 
                           REG_31_15_port);
   REG_reg_31_14_inst : DLH_X1 port map( G => n82, D => n1818, Q => 
                           REG_31_14_port);
   REG_reg_31_13_inst : DLH_X1 port map( G => n82, D => n1819, Q => 
                           REG_31_13_port);
   REG_reg_31_12_inst : DLH_X1 port map( G => n82, D => n1820, Q => 
                           REG_31_12_port);
   REG_reg_31_11_inst : DLH_X1 port map( G => n82, D => n1821, Q => 
                           REG_31_11_port);
   REG_reg_31_10_inst : DLH_X1 port map( G => n82, D => n1822, Q => 
                           REG_31_10_port);
   REG_reg_31_9_inst : DLH_X1 port map( G => n82, D => n1823, Q => 
                           REG_31_9_port);
   REG_reg_31_8_inst : DLH_X1 port map( G => n82, D => n1824, Q => 
                           REG_31_8_port);
   REG_reg_31_7_inst : DLH_X1 port map( G => n82, D => n1825, Q => 
                           REG_31_7_port);
   REG_reg_31_6_inst : DLH_X1 port map( G => n82, D => n1826, Q => 
                           REG_31_6_port);
   REG_reg_31_5_inst : DLH_X1 port map( G => n82, D => n1827, Q => 
                           REG_31_5_port);
   REG_reg_31_4_inst : DLH_X1 port map( G => n82, D => n1828, Q => 
                           REG_31_4_port);
   REG_reg_31_3_inst : DLH_X1 port map( G => n82, D => n1829, Q => 
                           REG_31_3_port);
   REG_reg_31_2_inst : DLH_X1 port map( G => n82, D => n1830, Q => 
                           REG_31_2_port);
   REG_reg_31_1_inst : DLH_X1 port map( G => n82, D => n1831, Q => 
                           REG_31_1_port);
   REG_reg_31_0_inst : DLH_X1 port map( G => n82, D => n1832, Q => 
                           REG_31_0_port);
   OUT2_reg_31_inst : DLH_X1 port map( G => N317, D => N284, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => N317, D => N285, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => N317, D => N286, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => N317, D => N287, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => N317, D => N288, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => N317, D => N289, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => N317, D => N290, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => N317, D => N291, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => N317, D => N292, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => N317, D => N293, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => N317, D => N294, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => N317, D => N295, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => N317, D => N296, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => N317, D => N297, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => N317, D => N298, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => N317, D => N299, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => N317, D => N300, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => N317, D => N301, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => N317, D => N302, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => N317, D => N303, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => N317, D => N304, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => N317, D => N305, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => N317, D => N306, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => N317, D => N307, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => N317, D => N308, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => N317, D => N309, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => N317, D => N310, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => N317, D => N311, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => N317, D => N312, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => N317, D => N313, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => N317, D => N314, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => N317, D => N315, Q => OUT2(0));
   OUT1_reg_31_inst : DLH_X1 port map( G => N316, D => N252, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => N316, D => N253, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => N316, D => N254, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => N316, D => N255, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => N316, D => N256, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => N316, D => N257, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => N316, D => N258, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => N316, D => N259, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => N316, D => N260, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => N316, D => N261, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => N316, D => N262, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => N316, D => N263, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => N316, D => N264, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => N316, D => N265, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => N316, D => N266, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => N316, D => N267, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => N316, D => N268, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => N316, D => N269, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => N316, D => N270, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => N316, D => N271, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => N316, D => N272, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => N316, D => N273, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => N316, D => N274, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => N316, D => N275, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => N316, D => N276, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => N316, D => N277, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => N316, D => N278, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => N316, D => N279, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => N316, D => N280, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => N316, D => N281, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => N316, D => N282, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => N316, D => N283, Q => OUT1(0));
   U3 : OR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n1);
   U4 : OR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n2);
   U5 : OR2_X1 port map( A1 => n1063, A2 => ADD_RD1(4), ZN => n3);
   U6 : OR2_X1 port map( A1 => n1745, A2 => ADD_RD2(4), ZN => n4);
   U7 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n1068, ZN => n5);
   U8 : AND2_X1 port map( A1 => n1067, A2 => ADD_RD2(0), ZN => n6);
   U9 : AND2_X1 port map( A1 => n1070, A2 => ADD_RD2(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n1069, A2 => ADD_RD2(0), ZN => n8);
   U11 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n386, ZN => n9);
   U12 : AND2_X1 port map( A1 => n386, A2 => n1066, ZN => n10);
   U13 : AND2_X1 port map( A1 => n1068, A2 => n1748, ZN => n11);
   U14 : AND2_X1 port map( A1 => n1069, A2 => n1748, ZN => n12);
   U15 : AND2_X1 port map( A1 => n385, A2 => ADD_RD1(0), ZN => n13);
   U16 : AND2_X1 port map( A1 => n388, A2 => ADD_RD1(0), ZN => n14);
   U17 : AND2_X1 port map( A1 => n387, A2 => ADD_RD1(0), ZN => n15);
   U18 : AND2_X1 port map( A1 => n385, A2 => n1066, ZN => n16);
   U19 : AND2_X1 port map( A1 => n388, A2 => n1066, ZN => n17);
   U20 : AND2_X1 port map( A1 => n387, A2 => n1066, ZN => n18);
   U21 : AND2_X1 port map( A1 => n1067, A2 => n1748, ZN => n19);
   U22 : AND2_X1 port map( A1 => n1070, A2 => n1748, ZN => n20);
   U23 : INV_X1 port map( A => N214, ZN => n21);
   U24 : INV_X1 port map( A => n21, ZN => n22);
   U25 : INV_X1 port map( A => N213, ZN => n23);
   U26 : INV_X1 port map( A => n23, ZN => n24);
   U27 : INV_X1 port map( A => N212, ZN => n25);
   U28 : INV_X1 port map( A => n25, ZN => n26);
   U29 : INV_X1 port map( A => N211, ZN => n27);
   U30 : INV_X1 port map( A => n27, ZN => n28);
   U31 : INV_X1 port map( A => N210, ZN => n29);
   U32 : INV_X1 port map( A => n29, ZN => n30);
   U33 : INV_X1 port map( A => N209, ZN => n31);
   U34 : INV_X1 port map( A => n31, ZN => n32);
   U35 : INV_X1 port map( A => N215, ZN => n33);
   U36 : INV_X1 port map( A => n33, ZN => n34);
   U37 : INV_X1 port map( A => N208, ZN => n35);
   U38 : INV_X1 port map( A => n35, ZN => n36);
   U39 : INV_X1 port map( A => N207, ZN => n37);
   U40 : INV_X1 port map( A => n37, ZN => n38);
   U41 : INV_X1 port map( A => N206, ZN => n39);
   U42 : INV_X1 port map( A => n39, ZN => n40);
   U43 : INV_X1 port map( A => N205, ZN => n41);
   U44 : INV_X1 port map( A => n41, ZN => n42);
   U45 : INV_X1 port map( A => N204, ZN => n43);
   U46 : INV_X1 port map( A => n43, ZN => n44);
   U47 : INV_X1 port map( A => N203, ZN => n45);
   U48 : INV_X1 port map( A => n45, ZN => n46);
   U49 : INV_X1 port map( A => N202, ZN => n47);
   U50 : INV_X1 port map( A => n47, ZN => n48);
   U51 : INV_X1 port map( A => N201, ZN => n49);
   U52 : INV_X1 port map( A => n49, ZN => n50);
   U53 : INV_X1 port map( A => N200, ZN => n51);
   U54 : INV_X1 port map( A => n51, ZN => n52);
   U55 : INV_X1 port map( A => N199, ZN => n53);
   U56 : INV_X1 port map( A => n53, ZN => n54);
   U57 : INV_X1 port map( A => N198, ZN => n55);
   U58 : INV_X1 port map( A => n55, ZN => n56);
   U59 : INV_X1 port map( A => N197, ZN => n57);
   U60 : INV_X1 port map( A => n57, ZN => n58);
   U61 : INV_X1 port map( A => N196, ZN => n59);
   U62 : INV_X1 port map( A => n59, ZN => n60);
   U63 : INV_X1 port map( A => N195, ZN => n61);
   U64 : INV_X1 port map( A => n61, ZN => n62);
   U65 : INV_X1 port map( A => N194, ZN => n63);
   U66 : INV_X1 port map( A => n63, ZN => n64);
   U67 : INV_X1 port map( A => N193, ZN => n65);
   U68 : INV_X1 port map( A => n65, ZN => n66);
   U69 : INV_X1 port map( A => N192, ZN => n67);
   U70 : INV_X1 port map( A => n67, ZN => n68);
   U71 : INV_X1 port map( A => N191, ZN => n69);
   U72 : INV_X1 port map( A => n69, ZN => n70);
   U73 : INV_X1 port map( A => N190, ZN => n71);
   U74 : INV_X1 port map( A => n71, ZN => n72);
   U75 : INV_X1 port map( A => N217, ZN => n73);
   U76 : INV_X1 port map( A => n73, ZN => n74);
   U77 : INV_X1 port map( A => N216, ZN => n75);
   U78 : INV_X1 port map( A => n75, ZN => n76);
   U79 : INV_X1 port map( A => N189, ZN => n77);
   U80 : INV_X1 port map( A => n77, ZN => n78);
   U81 : INV_X1 port map( A => N188, ZN => n79);
   U82 : INV_X1 port map( A => n79, ZN => n80);
   U83 : INV_X1 port map( A => N155, ZN => n81);
   U84 : INV_X1 port map( A => n81, ZN => n82);
   U85 : INV_X2 port map( A => n3, ZN => n83);
   U86 : INV_X2 port map( A => n4, ZN => n84);
   U87 : INV_X2 port map( A => n1, ZN => n85);
   U88 : INV_X2 port map( A => n2, ZN => n86);
   U89 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n1741);
   U90 : NAND2_X2 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n1059);
   U91 : OAI21_X4 port map( B1 => n1782, B2 => n1781, A => n379, ZN => N218);
   U92 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => n1745, ZN => n1743);
   U93 : NAND2_X2 port map( A1 => ADD_RD1(4), A2 => n1063, ZN => n1061);
   U94 : OR3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(4), A3 => n1783, ZN => 
                           n1781);
   U95 : INV_X2 port map( A => n1781, ZN => n87);
   U96 : BUF_X1 port map( A => n374, Z => n373);
   U97 : BUF_X1 port map( A => n356, Z => n355);
   U98 : BUF_X1 port map( A => n374, Z => n372);
   U99 : BUF_X1 port map( A => n356, Z => n354);
   U100 : BUF_X1 port map( A => n374, Z => n371);
   U101 : BUF_X1 port map( A => n356, Z => n353);
   U102 : BUF_X1 port map( A => n338, Z => n337);
   U103 : BUF_X1 port map( A => n320, Z => n319);
   U104 : BUF_X1 port map( A => n338, Z => n336);
   U105 : BUF_X1 port map( A => n320, Z => n318);
   U106 : BUF_X1 port map( A => n338, Z => n335);
   U107 : BUF_X1 port map( A => n320, Z => n317_port);
   U108 : BUF_X1 port map( A => n12, Z => n374);
   U109 : BUF_X1 port map( A => n20, Z => n356);
   U110 : BUF_X1 port map( A => n19, Z => n338);
   U111 : BUF_X1 port map( A => n11, Z => n320);
   U112 : BUF_X1 port map( A => n376, Z => n383);
   U113 : BUF_X1 port map( A => n376, Z => n384);
   U114 : BUF_X1 port map( A => n230_port, Z => n229_port);
   U115 : BUF_X1 port map( A => n212_port, Z => n211_port);
   U116 : BUF_X1 port map( A => n230_port, Z => n228_port);
   U117 : BUF_X1 port map( A => n212_port, Z => n210_port);
   U118 : BUF_X1 port map( A => n230_port, Z => n227_port);
   U119 : BUF_X1 port map( A => n212_port, Z => n209_port);
   U120 : BUF_X1 port map( A => n194_port, Z => n193_port);
   U121 : BUF_X1 port map( A => n176, Z => n175);
   U122 : BUF_X1 port map( A => n194_port, Z => n192_port);
   U123 : BUF_X1 port map( A => n176, Z => n174);
   U124 : BUF_X1 port map( A => n194_port, Z => n191_port);
   U125 : BUF_X1 port map( A => n176, Z => n173);
   U126 : BUF_X1 port map( A => n302_port, Z => n301_port);
   U127 : BUF_X1 port map( A => n284_port, Z => n283_port);
   U128 : BUF_X1 port map( A => n266_port, Z => n265_port);
   U129 : BUF_X1 port map( A => n248_port, Z => n247_port);
   U130 : BUF_X1 port map( A => n302_port, Z => n300_port);
   U131 : BUF_X1 port map( A => n284_port, Z => n282_port);
   U132 : BUF_X1 port map( A => n266_port, Z => n264_port);
   U133 : BUF_X1 port map( A => n248_port, Z => n246_port);
   U134 : BUF_X1 port map( A => n302_port, Z => n299_port);
   U135 : BUF_X1 port map( A => n284_port, Z => n281_port);
   U136 : BUF_X1 port map( A => n266_port, Z => n263_port);
   U137 : BUF_X1 port map( A => n248_port, Z => n245_port);
   U138 : BUF_X1 port map( A => n375, Z => n370);
   U139 : BUF_X1 port map( A => n357, Z => n352);
   U140 : BUF_X1 port map( A => n339, Z => n334);
   U141 : BUF_X1 port map( A => n321, Z => n316_port);
   U142 : BUF_X1 port map( A => n8, Z => n302_port);
   U143 : BUF_X1 port map( A => n7, Z => n284_port);
   U144 : BUF_X1 port map( A => n6, Z => n266_port);
   U145 : BUF_X1 port map( A => n5, Z => n248_port);
   U146 : BUF_X1 port map( A => n18, Z => n230_port);
   U147 : BUF_X1 port map( A => n17, Z => n212_port);
   U148 : BUF_X1 port map( A => n16, Z => n194_port);
   U149 : BUF_X1 port map( A => n10, Z => n176);
   U150 : BUF_X1 port map( A => n158, Z => n157);
   U151 : BUF_X1 port map( A => n140, Z => n139);
   U152 : BUF_X1 port map( A => n122, Z => n121);
   U153 : BUF_X1 port map( A => n104, Z => n103);
   U154 : BUF_X1 port map( A => n158, Z => n156);
   U155 : BUF_X1 port map( A => n140, Z => n138);
   U156 : BUF_X1 port map( A => n122, Z => n120);
   U157 : BUF_X1 port map( A => n104, Z => n102);
   U158 : BUF_X1 port map( A => n158, Z => n155_port);
   U159 : BUF_X1 port map( A => n140, Z => n137);
   U160 : BUF_X1 port map( A => n122, Z => n119);
   U161 : BUF_X1 port map( A => n104, Z => n101);
   U162 : BUF_X1 port map( A => n231_port, Z => n226_port);
   U163 : BUF_X1 port map( A => n213_port, Z => n208_port);
   U164 : BUF_X1 port map( A => n195_port, Z => n190_port);
   U165 : BUF_X1 port map( A => n177, Z => n172);
   U166 : BUF_X1 port map( A => n303_port, Z => n298_port);
   U167 : BUF_X1 port map( A => n285_port, Z => n280_port);
   U168 : BUF_X1 port map( A => n267_port, Z => n262_port);
   U169 : BUF_X1 port map( A => n249_port, Z => n244_port);
   U170 : BUF_X1 port map( A => n9, Z => n104);
   U171 : BUF_X1 port map( A => n15, Z => n158);
   U172 : BUF_X1 port map( A => n14, Z => n140);
   U173 : BUF_X1 port map( A => n13, Z => n122);
   U174 : BUF_X1 port map( A => n159, Z => n154);
   U175 : BUF_X1 port map( A => n141, Z => n136);
   U176 : BUF_X1 port map( A => n123, Z => n118);
   U177 : BUF_X1 port map( A => n105, Z => n100);
   U178 : BUF_X1 port map( A => n373, Z => n358);
   U179 : BUF_X1 port map( A => n372, Z => n361);
   U180 : BUF_X1 port map( A => n372, Z => n362);
   U181 : BUF_X1 port map( A => n371, Z => n365);
   U182 : BUF_X1 port map( A => n371, Z => n366);
   U183 : BUF_X1 port map( A => n337, Z => n322);
   U184 : BUF_X1 port map( A => n373, Z => n359);
   U185 : BUF_X1 port map( A => n337, Z => n323);
   U186 : BUF_X1 port map( A => n373, Z => n360);
   U187 : BUF_X1 port map( A => n337, Z => n324);
   U188 : BUF_X1 port map( A => n336, Z => n325);
   U189 : BUF_X1 port map( A => n336, Z => n326);
   U190 : BUF_X1 port map( A => n372, Z => n363);
   U191 : BUF_X1 port map( A => n336, Z => n327);
   U192 : BUF_X1 port map( A => n371, Z => n364);
   U193 : BUF_X1 port map( A => n335, Z => n328);
   U194 : BUF_X1 port map( A => n335, Z => n329);
   U195 : BUF_X1 port map( A => n335, Z => n330);
   U196 : BUF_X1 port map( A => n355, Z => n340);
   U197 : BUF_X1 port map( A => n354, Z => n343);
   U198 : BUF_X1 port map( A => n354, Z => n344);
   U199 : BUF_X1 port map( A => n353, Z => n347);
   U200 : BUF_X1 port map( A => n353, Z => n348);
   U201 : BUF_X1 port map( A => n319, Z => n304_port);
   U202 : BUF_X1 port map( A => n355, Z => n341);
   U203 : BUF_X1 port map( A => n319, Z => n305_port);
   U204 : BUF_X1 port map( A => n355, Z => n342);
   U205 : BUF_X1 port map( A => n319, Z => n306_port);
   U206 : BUF_X1 port map( A => n318, Z => n307_port);
   U207 : BUF_X1 port map( A => n318, Z => n308_port);
   U208 : BUF_X1 port map( A => n354, Z => n345);
   U209 : BUF_X1 port map( A => n318, Z => n309_port);
   U210 : BUF_X1 port map( A => n353, Z => n346);
   U211 : BUF_X1 port map( A => n317_port, Z => n310_port);
   U212 : BUF_X1 port map( A => n317_port, Z => n311_port);
   U213 : BUF_X1 port map( A => n317_port, Z => n312_port);
   U214 : BUF_X1 port map( A => n229_port, Z => n214_port);
   U215 : BUF_X1 port map( A => n228_port, Z => n217_port);
   U216 : BUF_X1 port map( A => n228_port, Z => n218_port);
   U217 : BUF_X1 port map( A => n227_port, Z => n221_port);
   U218 : BUF_X1 port map( A => n227_port, Z => n222_port);
   U219 : BUF_X1 port map( A => n193_port, Z => n178);
   U220 : BUF_X1 port map( A => n229_port, Z => n215_port);
   U221 : BUF_X1 port map( A => n193_port, Z => n179);
   U222 : BUF_X1 port map( A => n229_port, Z => n216_port);
   U223 : BUF_X1 port map( A => n193_port, Z => n180);
   U224 : BUF_X1 port map( A => n192_port, Z => n181);
   U225 : BUF_X1 port map( A => n192_port, Z => n182);
   U226 : BUF_X1 port map( A => n228_port, Z => n219_port);
   U227 : BUF_X1 port map( A => n192_port, Z => n183);
   U228 : BUF_X1 port map( A => n227_port, Z => n220_port);
   U229 : BUF_X1 port map( A => n191_port, Z => n184);
   U230 : BUF_X1 port map( A => n191_port, Z => n185);
   U231 : BUF_X1 port map( A => n191_port, Z => n186);
   U232 : BUF_X1 port map( A => n301_port, Z => n286_port);
   U233 : BUF_X1 port map( A => n265_port, Z => n250_port);
   U234 : BUF_X1 port map( A => n301_port, Z => n287_port);
   U235 : BUF_X1 port map( A => n265_port, Z => n251);
   U236 : BUF_X1 port map( A => n301_port, Z => n288_port);
   U237 : BUF_X1 port map( A => n265_port, Z => n252_port);
   U238 : BUF_X1 port map( A => n300_port, Z => n289_port);
   U239 : BUF_X1 port map( A => n264_port, Z => n253_port);
   U240 : BUF_X1 port map( A => n300_port, Z => n290_port);
   U241 : BUF_X1 port map( A => n264_port, Z => n254_port);
   U242 : BUF_X1 port map( A => n300_port, Z => n291_port);
   U243 : BUF_X1 port map( A => n264_port, Z => n255_port);
   U244 : BUF_X1 port map( A => n299_port, Z => n292_port);
   U245 : BUF_X1 port map( A => n263_port, Z => n256_port);
   U246 : BUF_X1 port map( A => n299_port, Z => n293_port);
   U247 : BUF_X1 port map( A => n263_port, Z => n257_port);
   U248 : BUF_X1 port map( A => n299_port, Z => n294_port);
   U249 : BUF_X1 port map( A => n263_port, Z => n258_port);
   U250 : BUF_X1 port map( A => n370, Z => n367);
   U251 : BUF_X1 port map( A => n334, Z => n331);
   U252 : BUF_X1 port map( A => n370, Z => n368);
   U253 : BUF_X1 port map( A => n334, Z => n332);
   U254 : BUF_X1 port map( A => n384, Z => n377);
   U255 : BUF_X1 port map( A => n384, Z => n378);
   U256 : BUF_X1 port map( A => n384, Z => n379);
   U257 : BUF_X1 port map( A => n383, Z => n380);
   U258 : BUF_X1 port map( A => n383, Z => n381);
   U259 : BUF_X1 port map( A => n211_port, Z => n196_port);
   U260 : BUF_X1 port map( A => n210_port, Z => n199_port);
   U261 : BUF_X1 port map( A => n210_port, Z => n200_port);
   U262 : BUF_X1 port map( A => n209_port, Z => n203_port);
   U263 : BUF_X1 port map( A => n209_port, Z => n204_port);
   U264 : BUF_X1 port map( A => n175, Z => n160);
   U265 : BUF_X1 port map( A => n211_port, Z => n197_port);
   U266 : BUF_X1 port map( A => n175, Z => n161);
   U267 : BUF_X1 port map( A => n211_port, Z => n198_port);
   U268 : BUF_X1 port map( A => n175, Z => n162);
   U269 : BUF_X1 port map( A => n174, Z => n163);
   U270 : BUF_X1 port map( A => n174, Z => n164);
   U271 : BUF_X1 port map( A => n210_port, Z => n201_port);
   U272 : BUF_X1 port map( A => n174, Z => n165);
   U273 : BUF_X1 port map( A => n209_port, Z => n202_port);
   U274 : BUF_X1 port map( A => n173, Z => n166);
   U275 : BUF_X1 port map( A => n173, Z => n167);
   U276 : BUF_X1 port map( A => n173, Z => n168);
   U277 : BUF_X1 port map( A => n283_port, Z => n268_port);
   U278 : BUF_X1 port map( A => n247_port, Z => n232_port);
   U279 : BUF_X1 port map( A => n283_port, Z => n269_port);
   U280 : BUF_X1 port map( A => n247_port, Z => n233_port);
   U281 : BUF_X1 port map( A => n283_port, Z => n270_port);
   U282 : BUF_X1 port map( A => n247_port, Z => n234_port);
   U283 : BUF_X1 port map( A => n282_port, Z => n271_port);
   U284 : BUF_X1 port map( A => n246_port, Z => n235_port);
   U285 : BUF_X1 port map( A => n282_port, Z => n272_port);
   U286 : BUF_X1 port map( A => n246_port, Z => n236_port);
   U287 : BUF_X1 port map( A => n282_port, Z => n273_port);
   U288 : BUF_X1 port map( A => n246_port, Z => n237_port);
   U289 : BUF_X1 port map( A => n281_port, Z => n274_port);
   U290 : BUF_X1 port map( A => n245_port, Z => n238_port);
   U291 : BUF_X1 port map( A => n281_port, Z => n275_port);
   U292 : BUF_X1 port map( A => n245_port, Z => n239_port);
   U293 : BUF_X1 port map( A => n281_port, Z => n276_port);
   U294 : BUF_X1 port map( A => n245_port, Z => n240_port);
   U295 : BUF_X1 port map( A => n352, Z => n349);
   U296 : BUF_X1 port map( A => n316_port, Z => n313_port);
   U297 : BUF_X1 port map( A => n352, Z => n350);
   U298 : BUF_X1 port map( A => n316_port, Z => n314_port);
   U299 : BUF_X1 port map( A => n383, Z => n382);
   U300 : BUF_X1 port map( A => n370, Z => n369);
   U301 : BUF_X1 port map( A => n334, Z => n333);
   U302 : BUF_X1 port map( A => n352, Z => n351);
   U303 : BUF_X1 port map( A => n316_port, Z => n315_port);
   U304 : BUF_X1 port map( A => n12, Z => n375);
   U305 : BUF_X1 port map( A => n20, Z => n357);
   U306 : BUF_X1 port map( A => n19, Z => n339);
   U307 : BUF_X1 port map( A => n11, Z => n321);
   U308 : BUF_X1 port map( A => n157, Z => n142);
   U309 : BUF_X1 port map( A => n121, Z => n106);
   U310 : BUF_X1 port map( A => n157, Z => n143);
   U311 : BUF_X1 port map( A => n121, Z => n107);
   U312 : BUF_X1 port map( A => n157, Z => n144);
   U313 : BUF_X1 port map( A => n121, Z => n108);
   U314 : BUF_X1 port map( A => n156, Z => n145);
   U315 : BUF_X1 port map( A => n120, Z => n109);
   U316 : BUF_X1 port map( A => n156, Z => n146);
   U317 : BUF_X1 port map( A => n120, Z => n110);
   U318 : BUF_X1 port map( A => n156, Z => n147);
   U319 : BUF_X1 port map( A => n120, Z => n111);
   U320 : BUF_X1 port map( A => n155_port, Z => n148);
   U321 : BUF_X1 port map( A => n119, Z => n112);
   U322 : BUF_X1 port map( A => n155_port, Z => n149);
   U323 : BUF_X1 port map( A => n119, Z => n113);
   U324 : BUF_X1 port map( A => n155_port, Z => n150);
   U325 : BUF_X1 port map( A => n119, Z => n114);
   U326 : BUF_X1 port map( A => n226_port, Z => n223_port);
   U327 : BUF_X1 port map( A => n190_port, Z => n187);
   U328 : BUF_X1 port map( A => n226_port, Z => n224_port);
   U329 : BUF_X1 port map( A => n190_port, Z => n188_port);
   U330 : BUF_X1 port map( A => n298_port, Z => n295_port);
   U331 : BUF_X1 port map( A => n262_port, Z => n259_port);
   U332 : BUF_X1 port map( A => n298_port, Z => n296_port);
   U333 : BUF_X1 port map( A => n262_port, Z => n260_port);
   U334 : BUF_X1 port map( A => n139, Z => n124);
   U335 : BUF_X1 port map( A => n103, Z => n88);
   U336 : BUF_X1 port map( A => n139, Z => n125);
   U337 : BUF_X1 port map( A => n103, Z => n89);
   U338 : BUF_X1 port map( A => n139, Z => n126);
   U339 : BUF_X1 port map( A => n103, Z => n90);
   U340 : BUF_X1 port map( A => n138, Z => n127);
   U341 : BUF_X1 port map( A => n102, Z => n91);
   U342 : BUF_X1 port map( A => n138, Z => n128);
   U343 : BUF_X1 port map( A => n102, Z => n92);
   U344 : BUF_X1 port map( A => n138, Z => n129);
   U345 : BUF_X1 port map( A => n102, Z => n93);
   U346 : BUF_X1 port map( A => n137, Z => n130);
   U347 : BUF_X1 port map( A => n101, Z => n94);
   U348 : BUF_X1 port map( A => n137, Z => n131);
   U349 : BUF_X1 port map( A => n101, Z => n95);
   U350 : BUF_X1 port map( A => n137, Z => n132);
   U351 : BUF_X1 port map( A => n101, Z => n96);
   U352 : BUF_X1 port map( A => n208_port, Z => n205_port);
   U353 : BUF_X1 port map( A => n172, Z => n169);
   U354 : BUF_X1 port map( A => n208_port, Z => n206_port);
   U355 : BUF_X1 port map( A => n172, Z => n170);
   U356 : BUF_X1 port map( A => n280_port, Z => n277_port);
   U357 : BUF_X1 port map( A => n244_port, Z => n241_port);
   U358 : BUF_X1 port map( A => n280_port, Z => n278_port);
   U359 : BUF_X1 port map( A => n244_port, Z => n242_port);
   U360 : BUF_X1 port map( A => n226_port, Z => n225_port);
   U361 : BUF_X1 port map( A => n190_port, Z => n189_port);
   U362 : BUF_X1 port map( A => n298_port, Z => n297_port);
   U363 : BUF_X1 port map( A => n262_port, Z => n261_port);
   U364 : BUF_X1 port map( A => n208_port, Z => n207_port);
   U365 : BUF_X1 port map( A => n172, Z => n171);
   U366 : BUF_X1 port map( A => n280_port, Z => n279_port);
   U367 : BUF_X1 port map( A => n244_port, Z => n243_port);
   U368 : BUF_X1 port map( A => n18, Z => n231_port);
   U369 : BUF_X1 port map( A => n17, Z => n213_port);
   U370 : BUF_X1 port map( A => n16, Z => n195_port);
   U371 : BUF_X1 port map( A => n10, Z => n177);
   U372 : BUF_X1 port map( A => n8, Z => n303_port);
   U373 : BUF_X1 port map( A => n7, Z => n285_port);
   U374 : BUF_X1 port map( A => n6, Z => n267_port);
   U375 : BUF_X1 port map( A => n5, Z => n249_port);
   U376 : BUF_X1 port map( A => RST, Z => n376);
   U377 : BUF_X1 port map( A => n154, Z => n151);
   U378 : BUF_X1 port map( A => n118, Z => n115);
   U379 : BUF_X1 port map( A => n154, Z => n152);
   U380 : BUF_X1 port map( A => n118, Z => n116);
   U381 : BUF_X1 port map( A => n136, Z => n133);
   U382 : BUF_X1 port map( A => n100, Z => n97);
   U383 : BUF_X1 port map( A => n136, Z => n134);
   U384 : BUF_X1 port map( A => n100, Z => n98);
   U385 : BUF_X1 port map( A => n154, Z => n153);
   U386 : BUF_X1 port map( A => n118, Z => n117);
   U387 : BUF_X1 port map( A => n136, Z => n135);
   U388 : BUF_X1 port map( A => n100, Z => n99);
   U389 : INV_X1 port map( A => ADD_RD2(0), ZN => n1748);
   U390 : INV_X1 port map( A => ADD_RD2(1), ZN => n1747);
   U391 : INV_X1 port map( A => ADD_RD2(3), ZN => n1745);
   U392 : INV_X1 port map( A => ADD_RD2(2), ZN => n1746);
   U393 : BUF_X1 port map( A => n15, Z => n159);
   U394 : BUF_X1 port map( A => n14, Z => n141);
   U395 : BUF_X1 port map( A => n13, Z => n123);
   U396 : BUF_X1 port map( A => n9, Z => n105);
   U397 : INV_X1 port map( A => ADD_RD1(0), ZN => n1066);
   U398 : INV_X1 port map( A => ADD_RD1(2), ZN => n1064);
   U399 : INV_X1 port map( A => ADD_RD1(3), ZN => n1063);
   U400 : INV_X1 port map( A => ADD_RD1(1), ZN => n1065);
   U401 : NOR2_X1 port map( A1 => n1064, A2 => ADD_RD1(1), ZN => n385);
   U402 : NOR2_X1 port map( A1 => n1064, A2 => n1065, ZN => n386);
   U403 : AOI22_X1 port map( A1 => REG_21_0_port, A2 => n106, B1 => 
                           REG_23_0_port, B2 => n88, ZN => n392);
   U404 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n387);
   U405 : NOR2_X1 port map( A1 => n1065, A2 => ADD_RD1(2), ZN => n388);
   U406 : AOI22_X1 port map( A1 => REG_17_0_port, A2 => n142, B1 => 
                           REG_19_0_port, B2 => n124, ZN => n391);
   U407 : AOI22_X1 port map( A1 => REG_20_0_port, A2 => n178, B1 => 
                           REG_22_0_port, B2 => n160, ZN => n390);
   U408 : AOI22_X1 port map( A1 => REG_16_0_port, A2 => n214_port, B1 => 
                           REG_18_0_port, B2 => n196_port, ZN => n389);
   U409 : AND4_X1 port map( A1 => n392, A2 => n391, A3 => n390, A4 => n389, ZN 
                           => n409);
   U410 : AOI22_X1 port map( A1 => REG_29_0_port, A2 => n106, B1 => 
                           REG_31_0_port, B2 => n88, ZN => n396);
   U411 : AOI22_X1 port map( A1 => REG_25_0_port, A2 => n142, B1 => 
                           REG_27_0_port, B2 => n124, ZN => n395);
   U412 : AOI22_X1 port map( A1 => REG_28_0_port, A2 => n178, B1 => 
                           REG_30_0_port, B2 => n160, ZN => n394);
   U413 : AOI22_X1 port map( A1 => REG_24_0_port, A2 => n214_port, B1 => 
                           REG_26_0_port, B2 => n196_port, ZN => n393);
   U414 : AND4_X1 port map( A1 => n396, A2 => n395, A3 => n394, A4 => n393, ZN 
                           => n408);
   U415 : AOI22_X1 port map( A1 => REG_5_0_port, A2 => n106, B1 => REG_7_0_port
                           , B2 => n88, ZN => n400);
   U416 : AOI22_X1 port map( A1 => REG_1_0_port, A2 => n142, B1 => REG_3_0_port
                           , B2 => n124, ZN => n399);
   U417 : AOI22_X1 port map( A1 => REG_4_0_port, A2 => n178, B1 => REG_6_0_port
                           , B2 => n160, ZN => n398);
   U418 : AOI22_X1 port map( A1 => REG_0_0_port, A2 => n214_port, B1 => 
                           REG_2_0_port, B2 => n196_port, ZN => n397);
   U419 : NAND4_X1 port map( A1 => n400, A2 => n399, A3 => n398, A4 => n397, ZN
                           => n406);
   U420 : AOI22_X1 port map( A1 => REG_13_0_port, A2 => n106, B1 => 
                           REG_15_0_port, B2 => n88, ZN => n404);
   U421 : AOI22_X1 port map( A1 => REG_9_0_port, A2 => n142, B1 => 
                           REG_11_0_port, B2 => n124, ZN => n403);
   U422 : AOI22_X1 port map( A1 => REG_12_0_port, A2 => n178, B1 => 
                           REG_14_0_port, B2 => n160, ZN => n402);
   U423 : AOI22_X1 port map( A1 => REG_8_0_port, A2 => n214_port, B1 => 
                           REG_10_0_port, B2 => n196_port, ZN => n401);
   U424 : NAND4_X1 port map( A1 => n404, A2 => n403, A3 => n402, A4 => n401, ZN
                           => n405);
   U425 : AOI22_X1 port map( A1 => n406, A2 => n85, B1 => n405, B2 => n83, ZN 
                           => n407);
   U426 : OAI221_X1 port map( B1 => n1061, B2 => n409, C1 => n1059, C2 => n408,
                           A => n407, ZN => N283);
   U427 : AOI22_X1 port map( A1 => REG_21_1_port, A2 => n106, B1 => 
                           REG_23_1_port, B2 => n88, ZN => n413);
   U428 : AOI22_X1 port map( A1 => REG_17_1_port, A2 => n142, B1 => 
                           REG_19_1_port, B2 => n124, ZN => n412);
   U429 : AOI22_X1 port map( A1 => REG_20_1_port, A2 => n178, B1 => 
                           REG_22_1_port, B2 => n160, ZN => n411);
   U430 : AOI22_X1 port map( A1 => REG_16_1_port, A2 => n214_port, B1 => 
                           REG_18_1_port, B2 => n196_port, ZN => n410);
   U431 : AND4_X1 port map( A1 => n413, A2 => n412, A3 => n411, A4 => n410, ZN 
                           => n430);
   U432 : AOI22_X1 port map( A1 => REG_29_1_port, A2 => n106, B1 => 
                           REG_31_1_port, B2 => n88, ZN => n417);
   U433 : AOI22_X1 port map( A1 => REG_25_1_port, A2 => n142, B1 => 
                           REG_27_1_port, B2 => n124, ZN => n416);
   U434 : AOI22_X1 port map( A1 => REG_28_1_port, A2 => n178, B1 => 
                           REG_30_1_port, B2 => n160, ZN => n415);
   U435 : AOI22_X1 port map( A1 => REG_24_1_port, A2 => n214_port, B1 => 
                           REG_26_1_port, B2 => n196_port, ZN => n414);
   U436 : AND4_X1 port map( A1 => n417, A2 => n416, A3 => n415, A4 => n414, ZN 
                           => n429);
   U437 : AOI22_X1 port map( A1 => REG_5_1_port, A2 => n106, B1 => REG_7_1_port
                           , B2 => n88, ZN => n421);
   U438 : AOI22_X1 port map( A1 => REG_1_1_port, A2 => n142, B1 => REG_3_1_port
                           , B2 => n124, ZN => n420);
   U439 : AOI22_X1 port map( A1 => REG_4_1_port, A2 => n178, B1 => REG_6_1_port
                           , B2 => n160, ZN => n419);
   U440 : AOI22_X1 port map( A1 => REG_0_1_port, A2 => n214_port, B1 => 
                           REG_2_1_port, B2 => n196_port, ZN => n418);
   U441 : NAND4_X1 port map( A1 => n421, A2 => n420, A3 => n419, A4 => n418, ZN
                           => n427);
   U442 : AOI22_X1 port map( A1 => REG_13_1_port, A2 => n106, B1 => 
                           REG_15_1_port, B2 => n88, ZN => n425);
   U443 : AOI22_X1 port map( A1 => REG_9_1_port, A2 => n142, B1 => 
                           REG_11_1_port, B2 => n124, ZN => n424);
   U444 : AOI22_X1 port map( A1 => REG_12_1_port, A2 => n178, B1 => 
                           REG_14_1_port, B2 => n160, ZN => n423);
   U445 : AOI22_X1 port map( A1 => REG_8_1_port, A2 => n214_port, B1 => 
                           REG_10_1_port, B2 => n196_port, ZN => n422);
   U446 : NAND4_X1 port map( A1 => n425, A2 => n424, A3 => n423, A4 => n422, ZN
                           => n426);
   U447 : AOI22_X1 port map( A1 => n427, A2 => n85, B1 => n426, B2 => n83, ZN 
                           => n428);
   U448 : OAI221_X1 port map( B1 => n1061, B2 => n430, C1 => n1059, C2 => n429,
                           A => n428, ZN => N282);
   U449 : AOI22_X1 port map( A1 => REG_21_2_port, A2 => n106, B1 => 
                           REG_23_2_port, B2 => n88, ZN => n434);
   U450 : AOI22_X1 port map( A1 => REG_17_2_port, A2 => n142, B1 => 
                           REG_19_2_port, B2 => n124, ZN => n433);
   U451 : AOI22_X1 port map( A1 => REG_20_2_port, A2 => n178, B1 => 
                           REG_22_2_port, B2 => n160, ZN => n432);
   U452 : AOI22_X1 port map( A1 => REG_16_2_port, A2 => n214_port, B1 => 
                           REG_18_2_port, B2 => n196_port, ZN => n431);
   U453 : AND4_X1 port map( A1 => n434, A2 => n433, A3 => n432, A4 => n431, ZN 
                           => n451);
   U454 : AOI22_X1 port map( A1 => REG_29_2_port, A2 => n106, B1 => 
                           REG_31_2_port, B2 => n88, ZN => n438);
   U455 : AOI22_X1 port map( A1 => REG_25_2_port, A2 => n142, B1 => 
                           REG_27_2_port, B2 => n124, ZN => n437);
   U456 : AOI22_X1 port map( A1 => REG_28_2_port, A2 => n178, B1 => 
                           REG_30_2_port, B2 => n160, ZN => n436);
   U457 : AOI22_X1 port map( A1 => REG_24_2_port, A2 => n214_port, B1 => 
                           REG_26_2_port, B2 => n196_port, ZN => n435);
   U458 : AND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN 
                           => n450);
   U459 : AOI22_X1 port map( A1 => REG_5_2_port, A2 => n106, B1 => REG_7_2_port
                           , B2 => n88, ZN => n442);
   U460 : AOI22_X1 port map( A1 => REG_1_2_port, A2 => n142, B1 => REG_3_2_port
                           , B2 => n124, ZN => n441);
   U461 : AOI22_X1 port map( A1 => REG_4_2_port, A2 => n178, B1 => REG_6_2_port
                           , B2 => n160, ZN => n440);
   U462 : AOI22_X1 port map( A1 => REG_0_2_port, A2 => n214_port, B1 => 
                           REG_2_2_port, B2 => n196_port, ZN => n439);
   U463 : NAND4_X1 port map( A1 => n442, A2 => n441, A3 => n440, A4 => n439, ZN
                           => n448);
   U464 : AOI22_X1 port map( A1 => REG_13_2_port, A2 => n107, B1 => 
                           REG_15_2_port, B2 => n89, ZN => n446);
   U465 : AOI22_X1 port map( A1 => REG_9_2_port, A2 => n143, B1 => 
                           REG_11_2_port, B2 => n125, ZN => n445);
   U466 : AOI22_X1 port map( A1 => REG_12_2_port, A2 => n179, B1 => 
                           REG_14_2_port, B2 => n161, ZN => n444);
   U467 : AOI22_X1 port map( A1 => REG_8_2_port, A2 => n215_port, B1 => 
                           REG_10_2_port, B2 => n197_port, ZN => n443);
   U468 : NAND4_X1 port map( A1 => n446, A2 => n445, A3 => n444, A4 => n443, ZN
                           => n447);
   U469 : AOI22_X1 port map( A1 => n448, A2 => n85, B1 => n447, B2 => n83, ZN 
                           => n449);
   U470 : OAI221_X1 port map( B1 => n1061, B2 => n451, C1 => n1059, C2 => n450,
                           A => n449, ZN => N281);
   U471 : AOI22_X1 port map( A1 => REG_21_3_port, A2 => n107, B1 => 
                           REG_23_3_port, B2 => n89, ZN => n455);
   U472 : AOI22_X1 port map( A1 => REG_17_3_port, A2 => n143, B1 => 
                           REG_19_3_port, B2 => n125, ZN => n454);
   U473 : AOI22_X1 port map( A1 => REG_20_3_port, A2 => n179, B1 => 
                           REG_22_3_port, B2 => n161, ZN => n453);
   U474 : AOI22_X1 port map( A1 => REG_16_3_port, A2 => n215_port, B1 => 
                           REG_18_3_port, B2 => n197_port, ZN => n452);
   U475 : AND4_X1 port map( A1 => n455, A2 => n454, A3 => n453, A4 => n452, ZN 
                           => n472);
   U476 : AOI22_X1 port map( A1 => REG_29_3_port, A2 => n107, B1 => 
                           REG_31_3_port, B2 => n89, ZN => n459);
   U477 : AOI22_X1 port map( A1 => REG_25_3_port, A2 => n143, B1 => 
                           REG_27_3_port, B2 => n125, ZN => n458);
   U478 : AOI22_X1 port map( A1 => REG_28_3_port, A2 => n179, B1 => 
                           REG_30_3_port, B2 => n161, ZN => n457);
   U479 : AOI22_X1 port map( A1 => REG_24_3_port, A2 => n215_port, B1 => 
                           REG_26_3_port, B2 => n197_port, ZN => n456);
   U480 : AND4_X1 port map( A1 => n459, A2 => n458, A3 => n457, A4 => n456, ZN 
                           => n471);
   U481 : AOI22_X1 port map( A1 => REG_5_3_port, A2 => n107, B1 => REG_7_3_port
                           , B2 => n89, ZN => n463);
   U482 : AOI22_X1 port map( A1 => REG_1_3_port, A2 => n143, B1 => REG_3_3_port
                           , B2 => n125, ZN => n462);
   U483 : AOI22_X1 port map( A1 => REG_4_3_port, A2 => n179, B1 => REG_6_3_port
                           , B2 => n161, ZN => n461);
   U484 : AOI22_X1 port map( A1 => REG_0_3_port, A2 => n215_port, B1 => 
                           REG_2_3_port, B2 => n197_port, ZN => n460);
   U485 : NAND4_X1 port map( A1 => n463, A2 => n462, A3 => n461, A4 => n460, ZN
                           => n469);
   U486 : AOI22_X1 port map( A1 => REG_13_3_port, A2 => n107, B1 => 
                           REG_15_3_port, B2 => n89, ZN => n467);
   U487 : AOI22_X1 port map( A1 => REG_9_3_port, A2 => n143, B1 => 
                           REG_11_3_port, B2 => n125, ZN => n466);
   U488 : AOI22_X1 port map( A1 => REG_12_3_port, A2 => n179, B1 => 
                           REG_14_3_port, B2 => n161, ZN => n465);
   U489 : AOI22_X1 port map( A1 => REG_8_3_port, A2 => n215_port, B1 => 
                           REG_10_3_port, B2 => n197_port, ZN => n464);
   U490 : NAND4_X1 port map( A1 => n467, A2 => n466, A3 => n465, A4 => n464, ZN
                           => n468);
   U491 : AOI22_X1 port map( A1 => n469, A2 => n85, B1 => n468, B2 => n83, ZN 
                           => n470);
   U492 : OAI221_X1 port map( B1 => n1061, B2 => n472, C1 => n1059, C2 => n471,
                           A => n470, ZN => N280);
   U493 : AOI22_X1 port map( A1 => REG_21_4_port, A2 => n107, B1 => 
                           REG_23_4_port, B2 => n89, ZN => n476);
   U494 : AOI22_X1 port map( A1 => REG_17_4_port, A2 => n143, B1 => 
                           REG_19_4_port, B2 => n125, ZN => n475);
   U495 : AOI22_X1 port map( A1 => REG_20_4_port, A2 => n179, B1 => 
                           REG_22_4_port, B2 => n161, ZN => n474);
   U496 : AOI22_X1 port map( A1 => REG_16_4_port, A2 => n215_port, B1 => 
                           REG_18_4_port, B2 => n197_port, ZN => n473);
   U497 : AND4_X1 port map( A1 => n476, A2 => n475, A3 => n474, A4 => n473, ZN 
                           => n493);
   U498 : AOI22_X1 port map( A1 => REG_29_4_port, A2 => n107, B1 => 
                           REG_31_4_port, B2 => n89, ZN => n480);
   U499 : AOI22_X1 port map( A1 => REG_25_4_port, A2 => n143, B1 => 
                           REG_27_4_port, B2 => n125, ZN => n479);
   U500 : AOI22_X1 port map( A1 => REG_28_4_port, A2 => n179, B1 => 
                           REG_30_4_port, B2 => n161, ZN => n478);
   U501 : AOI22_X1 port map( A1 => REG_24_4_port, A2 => n215_port, B1 => 
                           REG_26_4_port, B2 => n197_port, ZN => n477);
   U502 : AND4_X1 port map( A1 => n480, A2 => n479, A3 => n478, A4 => n477, ZN 
                           => n492);
   U503 : AOI22_X1 port map( A1 => REG_5_4_port, A2 => n107, B1 => REG_7_4_port
                           , B2 => n89, ZN => n484);
   U504 : AOI22_X1 port map( A1 => REG_1_4_port, A2 => n143, B1 => REG_3_4_port
                           , B2 => n125, ZN => n483);
   U505 : AOI22_X1 port map( A1 => REG_4_4_port, A2 => n179, B1 => REG_6_4_port
                           , B2 => n161, ZN => n482);
   U506 : AOI22_X1 port map( A1 => REG_0_4_port, A2 => n215_port, B1 => 
                           REG_2_4_port, B2 => n197_port, ZN => n481);
   U507 : NAND4_X1 port map( A1 => n484, A2 => n483, A3 => n482, A4 => n481, ZN
                           => n490);
   U508 : AOI22_X1 port map( A1 => REG_13_4_port, A2 => n107, B1 => 
                           REG_15_4_port, B2 => n89, ZN => n488);
   U509 : AOI22_X1 port map( A1 => REG_9_4_port, A2 => n143, B1 => 
                           REG_11_4_port, B2 => n125, ZN => n487);
   U510 : AOI22_X1 port map( A1 => REG_12_4_port, A2 => n179, B1 => 
                           REG_14_4_port, B2 => n161, ZN => n486);
   U511 : AOI22_X1 port map( A1 => REG_8_4_port, A2 => n215_port, B1 => 
                           REG_10_4_port, B2 => n197_port, ZN => n485);
   U512 : NAND4_X1 port map( A1 => n488, A2 => n487, A3 => n486, A4 => n485, ZN
                           => n489);
   U513 : AOI22_X1 port map( A1 => n490, A2 => n85, B1 => n489, B2 => n83, ZN 
                           => n491);
   U514 : OAI221_X1 port map( B1 => n1061, B2 => n493, C1 => n1059, C2 => n492,
                           A => n491, ZN => N279);
   U515 : AOI22_X1 port map( A1 => REG_21_5_port, A2 => n107, B1 => 
                           REG_23_5_port, B2 => n89, ZN => n497);
   U516 : AOI22_X1 port map( A1 => REG_17_5_port, A2 => n143, B1 => 
                           REG_19_5_port, B2 => n125, ZN => n496);
   U517 : AOI22_X1 port map( A1 => REG_20_5_port, A2 => n179, B1 => 
                           REG_22_5_port, B2 => n161, ZN => n495);
   U518 : AOI22_X1 port map( A1 => REG_16_5_port, A2 => n215_port, B1 => 
                           REG_18_5_port, B2 => n197_port, ZN => n494);
   U519 : AND4_X1 port map( A1 => n497, A2 => n496, A3 => n495, A4 => n494, ZN 
                           => n514);
   U520 : AOI22_X1 port map( A1 => REG_29_5_port, A2 => n107, B1 => 
                           REG_31_5_port, B2 => n89, ZN => n501);
   U521 : AOI22_X1 port map( A1 => REG_25_5_port, A2 => n143, B1 => 
                           REG_27_5_port, B2 => n125, ZN => n500);
   U522 : AOI22_X1 port map( A1 => REG_28_5_port, A2 => n179, B1 => 
                           REG_30_5_port, B2 => n161, ZN => n499);
   U523 : AOI22_X1 port map( A1 => REG_24_5_port, A2 => n215_port, B1 => 
                           REG_26_5_port, B2 => n197_port, ZN => n498);
   U524 : AND4_X1 port map( A1 => n501, A2 => n500, A3 => n499, A4 => n498, ZN 
                           => n513);
   U525 : AOI22_X1 port map( A1 => REG_5_5_port, A2 => n108, B1 => REG_7_5_port
                           , B2 => n90, ZN => n505);
   U526 : AOI22_X1 port map( A1 => REG_1_5_port, A2 => n144, B1 => REG_3_5_port
                           , B2 => n126, ZN => n504);
   U527 : AOI22_X1 port map( A1 => REG_4_5_port, A2 => n180, B1 => REG_6_5_port
                           , B2 => n162, ZN => n503);
   U528 : AOI22_X1 port map( A1 => REG_0_5_port, A2 => n216_port, B1 => 
                           REG_2_5_port, B2 => n198_port, ZN => n502);
   U529 : NAND4_X1 port map( A1 => n505, A2 => n504, A3 => n503, A4 => n502, ZN
                           => n511);
   U530 : AOI22_X1 port map( A1 => REG_13_5_port, A2 => n108, B1 => 
                           REG_15_5_port, B2 => n90, ZN => n509);
   U531 : AOI22_X1 port map( A1 => REG_9_5_port, A2 => n144, B1 => 
                           REG_11_5_port, B2 => n126, ZN => n508);
   U532 : AOI22_X1 port map( A1 => REG_12_5_port, A2 => n180, B1 => 
                           REG_14_5_port, B2 => n162, ZN => n507);
   U533 : AOI22_X1 port map( A1 => REG_8_5_port, A2 => n216_port, B1 => 
                           REG_10_5_port, B2 => n198_port, ZN => n506);
   U534 : NAND4_X1 port map( A1 => n509, A2 => n508, A3 => n507, A4 => n506, ZN
                           => n510);
   U535 : AOI22_X1 port map( A1 => n511, A2 => n85, B1 => n510, B2 => n83, ZN 
                           => n512);
   U536 : OAI221_X1 port map( B1 => n1061, B2 => n514, C1 => n1059, C2 => n513,
                           A => n512, ZN => N278);
   U537 : AOI22_X1 port map( A1 => REG_21_6_port, A2 => n108, B1 => 
                           REG_23_6_port, B2 => n90, ZN => n518);
   U538 : AOI22_X1 port map( A1 => REG_17_6_port, A2 => n144, B1 => 
                           REG_19_6_port, B2 => n126, ZN => n517);
   U539 : AOI22_X1 port map( A1 => REG_20_6_port, A2 => n180, B1 => 
                           REG_22_6_port, B2 => n162, ZN => n516);
   U540 : AOI22_X1 port map( A1 => REG_16_6_port, A2 => n216_port, B1 => 
                           REG_18_6_port, B2 => n198_port, ZN => n515);
   U541 : AND4_X1 port map( A1 => n518, A2 => n517, A3 => n516, A4 => n515, ZN 
                           => n535);
   U542 : AOI22_X1 port map( A1 => REG_29_6_port, A2 => n108, B1 => 
                           REG_31_6_port, B2 => n90, ZN => n522);
   U543 : AOI22_X1 port map( A1 => REG_25_6_port, A2 => n144, B1 => 
                           REG_27_6_port, B2 => n126, ZN => n521);
   U544 : AOI22_X1 port map( A1 => REG_28_6_port, A2 => n180, B1 => 
                           REG_30_6_port, B2 => n162, ZN => n520);
   U545 : AOI22_X1 port map( A1 => REG_24_6_port, A2 => n216_port, B1 => 
                           REG_26_6_port, B2 => n198_port, ZN => n519);
   U546 : AND4_X1 port map( A1 => n522, A2 => n521, A3 => n520, A4 => n519, ZN 
                           => n534);
   U547 : AOI22_X1 port map( A1 => REG_5_6_port, A2 => n108, B1 => REG_7_6_port
                           , B2 => n90, ZN => n526);
   U548 : AOI22_X1 port map( A1 => REG_1_6_port, A2 => n144, B1 => REG_3_6_port
                           , B2 => n126, ZN => n525);
   U549 : AOI22_X1 port map( A1 => REG_4_6_port, A2 => n180, B1 => REG_6_6_port
                           , B2 => n162, ZN => n524);
   U550 : AOI22_X1 port map( A1 => REG_0_6_port, A2 => n216_port, B1 => 
                           REG_2_6_port, B2 => n198_port, ZN => n523);
   U551 : NAND4_X1 port map( A1 => n526, A2 => n525, A3 => n524, A4 => n523, ZN
                           => n532);
   U552 : AOI22_X1 port map( A1 => REG_13_6_port, A2 => n108, B1 => 
                           REG_15_6_port, B2 => n90, ZN => n530);
   U553 : AOI22_X1 port map( A1 => REG_9_6_port, A2 => n144, B1 => 
                           REG_11_6_port, B2 => n126, ZN => n529);
   U554 : AOI22_X1 port map( A1 => REG_12_6_port, A2 => n180, B1 => 
                           REG_14_6_port, B2 => n162, ZN => n528);
   U555 : AOI22_X1 port map( A1 => REG_8_6_port, A2 => n216_port, B1 => 
                           REG_10_6_port, B2 => n198_port, ZN => n527);
   U556 : NAND4_X1 port map( A1 => n530, A2 => n529, A3 => n528, A4 => n527, ZN
                           => n531);
   U557 : AOI22_X1 port map( A1 => n532, A2 => n85, B1 => n531, B2 => n83, ZN 
                           => n533);
   U558 : OAI221_X1 port map( B1 => n1061, B2 => n535, C1 => n1059, C2 => n534,
                           A => n533, ZN => N277);
   U559 : AOI22_X1 port map( A1 => REG_21_7_port, A2 => n108, B1 => 
                           REG_23_7_port, B2 => n90, ZN => n539);
   U560 : AOI22_X1 port map( A1 => REG_17_7_port, A2 => n144, B1 => 
                           REG_19_7_port, B2 => n126, ZN => n538);
   U561 : AOI22_X1 port map( A1 => REG_20_7_port, A2 => n180, B1 => 
                           REG_22_7_port, B2 => n162, ZN => n537);
   U562 : AOI22_X1 port map( A1 => REG_16_7_port, A2 => n216_port, B1 => 
                           REG_18_7_port, B2 => n198_port, ZN => n536);
   U563 : AND4_X1 port map( A1 => n539, A2 => n538, A3 => n537, A4 => n536, ZN 
                           => n556);
   U564 : AOI22_X1 port map( A1 => REG_29_7_port, A2 => n108, B1 => 
                           REG_31_7_port, B2 => n90, ZN => n543);
   U565 : AOI22_X1 port map( A1 => REG_25_7_port, A2 => n144, B1 => 
                           REG_27_7_port, B2 => n126, ZN => n542);
   U566 : AOI22_X1 port map( A1 => REG_28_7_port, A2 => n180, B1 => 
                           REG_30_7_port, B2 => n162, ZN => n541);
   U567 : AOI22_X1 port map( A1 => REG_24_7_port, A2 => n216_port, B1 => 
                           REG_26_7_port, B2 => n198_port, ZN => n540);
   U568 : AND4_X1 port map( A1 => n543, A2 => n542, A3 => n541, A4 => n540, ZN 
                           => n555);
   U569 : AOI22_X1 port map( A1 => REG_5_7_port, A2 => n108, B1 => REG_7_7_port
                           , B2 => n90, ZN => n547);
   U570 : AOI22_X1 port map( A1 => REG_1_7_port, A2 => n144, B1 => REG_3_7_port
                           , B2 => n126, ZN => n546);
   U571 : AOI22_X1 port map( A1 => REG_4_7_port, A2 => n180, B1 => REG_6_7_port
                           , B2 => n162, ZN => n545);
   U572 : AOI22_X1 port map( A1 => REG_0_7_port, A2 => n216_port, B1 => 
                           REG_2_7_port, B2 => n198_port, ZN => n544);
   U573 : NAND4_X1 port map( A1 => n547, A2 => n546, A3 => n545, A4 => n544, ZN
                           => n553);
   U574 : AOI22_X1 port map( A1 => REG_13_7_port, A2 => n108, B1 => 
                           REG_15_7_port, B2 => n90, ZN => n551);
   U575 : AOI22_X1 port map( A1 => REG_9_7_port, A2 => n144, B1 => 
                           REG_11_7_port, B2 => n126, ZN => n550);
   U576 : AOI22_X1 port map( A1 => REG_12_7_port, A2 => n180, B1 => 
                           REG_14_7_port, B2 => n162, ZN => n549);
   U577 : AOI22_X1 port map( A1 => REG_8_7_port, A2 => n216_port, B1 => 
                           REG_10_7_port, B2 => n198_port, ZN => n548);
   U578 : NAND4_X1 port map( A1 => n551, A2 => n550, A3 => n549, A4 => n548, ZN
                           => n552);
   U579 : AOI22_X1 port map( A1 => n553, A2 => n85, B1 => n552, B2 => n83, ZN 
                           => n554);
   U580 : OAI221_X1 port map( B1 => n1061, B2 => n556, C1 => n1059, C2 => n555,
                           A => n554, ZN => N276);
   U581 : AOI22_X1 port map( A1 => REG_21_8_port, A2 => n108, B1 => 
                           REG_23_8_port, B2 => n90, ZN => n560);
   U582 : AOI22_X1 port map( A1 => REG_17_8_port, A2 => n144, B1 => 
                           REG_19_8_port, B2 => n126, ZN => n559);
   U583 : AOI22_X1 port map( A1 => REG_20_8_port, A2 => n180, B1 => 
                           REG_22_8_port, B2 => n162, ZN => n558);
   U584 : AOI22_X1 port map( A1 => REG_16_8_port, A2 => n216_port, B1 => 
                           REG_18_8_port, B2 => n198_port, ZN => n557);
   U585 : AND4_X1 port map( A1 => n560, A2 => n559, A3 => n558, A4 => n557, ZN 
                           => n577);
   U586 : AOI22_X1 port map( A1 => REG_29_8_port, A2 => n109, B1 => 
                           REG_31_8_port, B2 => n91, ZN => n564);
   U587 : AOI22_X1 port map( A1 => REG_25_8_port, A2 => n145, B1 => 
                           REG_27_8_port, B2 => n127, ZN => n563);
   U588 : AOI22_X1 port map( A1 => REG_28_8_port, A2 => n181, B1 => 
                           REG_30_8_port, B2 => n163, ZN => n562);
   U589 : AOI22_X1 port map( A1 => REG_24_8_port, A2 => n217_port, B1 => 
                           REG_26_8_port, B2 => n199_port, ZN => n561);
   U590 : AND4_X1 port map( A1 => n564, A2 => n563, A3 => n562, A4 => n561, ZN 
                           => n576);
   U591 : AOI22_X1 port map( A1 => REG_5_8_port, A2 => n109, B1 => REG_7_8_port
                           , B2 => n91, ZN => n568);
   U592 : AOI22_X1 port map( A1 => REG_1_8_port, A2 => n145, B1 => REG_3_8_port
                           , B2 => n127, ZN => n567);
   U593 : AOI22_X1 port map( A1 => REG_4_8_port, A2 => n181, B1 => REG_6_8_port
                           , B2 => n163, ZN => n566);
   U594 : AOI22_X1 port map( A1 => REG_0_8_port, A2 => n217_port, B1 => 
                           REG_2_8_port, B2 => n199_port, ZN => n565);
   U595 : NAND4_X1 port map( A1 => n568, A2 => n567, A3 => n566, A4 => n565, ZN
                           => n574);
   U596 : AOI22_X1 port map( A1 => REG_13_8_port, A2 => n109, B1 => 
                           REG_15_8_port, B2 => n91, ZN => n572);
   U597 : AOI22_X1 port map( A1 => REG_9_8_port, A2 => n145, B1 => 
                           REG_11_8_port, B2 => n127, ZN => n571);
   U598 : AOI22_X1 port map( A1 => REG_12_8_port, A2 => n181, B1 => 
                           REG_14_8_port, B2 => n163, ZN => n570);
   U599 : AOI22_X1 port map( A1 => REG_8_8_port, A2 => n217_port, B1 => 
                           REG_10_8_port, B2 => n199_port, ZN => n569);
   U600 : NAND4_X1 port map( A1 => n572, A2 => n571, A3 => n570, A4 => n569, ZN
                           => n573);
   U601 : AOI22_X1 port map( A1 => n574, A2 => n85, B1 => n573, B2 => n83, ZN 
                           => n575);
   U602 : OAI221_X1 port map( B1 => n1061, B2 => n577, C1 => n1059, C2 => n576,
                           A => n575, ZN => N275);
   U603 : AOI22_X1 port map( A1 => REG_21_9_port, A2 => n109, B1 => 
                           REG_23_9_port, B2 => n91, ZN => n581);
   U604 : AOI22_X1 port map( A1 => REG_17_9_port, A2 => n145, B1 => 
                           REG_19_9_port, B2 => n127, ZN => n580);
   U605 : AOI22_X1 port map( A1 => REG_20_9_port, A2 => n181, B1 => 
                           REG_22_9_port, B2 => n163, ZN => n579);
   U606 : AOI22_X1 port map( A1 => REG_16_9_port, A2 => n217_port, B1 => 
                           REG_18_9_port, B2 => n199_port, ZN => n578);
   U607 : AND4_X1 port map( A1 => n581, A2 => n580, A3 => n579, A4 => n578, ZN 
                           => n598);
   U608 : AOI22_X1 port map( A1 => REG_29_9_port, A2 => n109, B1 => 
                           REG_31_9_port, B2 => n91, ZN => n585);
   U609 : AOI22_X1 port map( A1 => REG_25_9_port, A2 => n145, B1 => 
                           REG_27_9_port, B2 => n127, ZN => n584);
   U610 : AOI22_X1 port map( A1 => REG_28_9_port, A2 => n181, B1 => 
                           REG_30_9_port, B2 => n163, ZN => n583);
   U611 : AOI22_X1 port map( A1 => REG_24_9_port, A2 => n217_port, B1 => 
                           REG_26_9_port, B2 => n199_port, ZN => n582);
   U612 : AND4_X1 port map( A1 => n585, A2 => n584, A3 => n583, A4 => n582, ZN 
                           => n597);
   U613 : AOI22_X1 port map( A1 => REG_5_9_port, A2 => n109, B1 => REG_7_9_port
                           , B2 => n91, ZN => n589);
   U614 : AOI22_X1 port map( A1 => REG_1_9_port, A2 => n145, B1 => REG_3_9_port
                           , B2 => n127, ZN => n588);
   U615 : AOI22_X1 port map( A1 => REG_4_9_port, A2 => n181, B1 => REG_6_9_port
                           , B2 => n163, ZN => n587);
   U616 : AOI22_X1 port map( A1 => REG_0_9_port, A2 => n217_port, B1 => 
                           REG_2_9_port, B2 => n199_port, ZN => n586);
   U617 : NAND4_X1 port map( A1 => n589, A2 => n588, A3 => n587, A4 => n586, ZN
                           => n595);
   U618 : AOI22_X1 port map( A1 => REG_13_9_port, A2 => n109, B1 => 
                           REG_15_9_port, B2 => n91, ZN => n593);
   U619 : AOI22_X1 port map( A1 => REG_9_9_port, A2 => n145, B1 => 
                           REG_11_9_port, B2 => n127, ZN => n592);
   U620 : AOI22_X1 port map( A1 => REG_12_9_port, A2 => n181, B1 => 
                           REG_14_9_port, B2 => n163, ZN => n591);
   U621 : AOI22_X1 port map( A1 => REG_8_9_port, A2 => n217_port, B1 => 
                           REG_10_9_port, B2 => n199_port, ZN => n590);
   U622 : NAND4_X1 port map( A1 => n593, A2 => n592, A3 => n591, A4 => n590, ZN
                           => n594);
   U623 : AOI22_X1 port map( A1 => n595, A2 => n85, B1 => n594, B2 => n83, ZN 
                           => n596);
   U624 : OAI221_X1 port map( B1 => n1061, B2 => n598, C1 => n1059, C2 => n597,
                           A => n596, ZN => N274);
   U625 : AOI22_X1 port map( A1 => REG_21_10_port, A2 => n109, B1 => 
                           REG_23_10_port, B2 => n91, ZN => n602);
   U626 : AOI22_X1 port map( A1 => REG_17_10_port, A2 => n145, B1 => 
                           REG_19_10_port, B2 => n127, ZN => n601);
   U627 : AOI22_X1 port map( A1 => REG_20_10_port, A2 => n181, B1 => 
                           REG_22_10_port, B2 => n163, ZN => n600);
   U628 : AOI22_X1 port map( A1 => REG_16_10_port, A2 => n217_port, B1 => 
                           REG_18_10_port, B2 => n199_port, ZN => n599);
   U629 : AND4_X1 port map( A1 => n602, A2 => n601, A3 => n600, A4 => n599, ZN 
                           => n619);
   U630 : AOI22_X1 port map( A1 => REG_29_10_port, A2 => n109, B1 => 
                           REG_31_10_port, B2 => n91, ZN => n606);
   U631 : AOI22_X1 port map( A1 => REG_25_10_port, A2 => n145, B1 => 
                           REG_27_10_port, B2 => n127, ZN => n605);
   U632 : AOI22_X1 port map( A1 => REG_28_10_port, A2 => n181, B1 => 
                           REG_30_10_port, B2 => n163, ZN => n604);
   U633 : AOI22_X1 port map( A1 => REG_24_10_port, A2 => n217_port, B1 => 
                           REG_26_10_port, B2 => n199_port, ZN => n603);
   U634 : AND4_X1 port map( A1 => n606, A2 => n605, A3 => n604, A4 => n603, ZN 
                           => n618);
   U635 : AOI22_X1 port map( A1 => REG_5_10_port, A2 => n109, B1 => 
                           REG_7_10_port, B2 => n91, ZN => n610);
   U636 : AOI22_X1 port map( A1 => REG_1_10_port, A2 => n145, B1 => 
                           REG_3_10_port, B2 => n127, ZN => n609);
   U637 : AOI22_X1 port map( A1 => REG_4_10_port, A2 => n181, B1 => 
                           REG_6_10_port, B2 => n163, ZN => n608);
   U638 : AOI22_X1 port map( A1 => REG_0_10_port, A2 => n217_port, B1 => 
                           REG_2_10_port, B2 => n199_port, ZN => n607);
   U639 : NAND4_X1 port map( A1 => n610, A2 => n609, A3 => n608, A4 => n607, ZN
                           => n616);
   U640 : AOI22_X1 port map( A1 => REG_13_10_port, A2 => n109, B1 => 
                           REG_15_10_port, B2 => n91, ZN => n614);
   U641 : AOI22_X1 port map( A1 => REG_9_10_port, A2 => n145, B1 => 
                           REG_11_10_port, B2 => n127, ZN => n613);
   U642 : AOI22_X1 port map( A1 => REG_12_10_port, A2 => n181, B1 => 
                           REG_14_10_port, B2 => n163, ZN => n612);
   U643 : AOI22_X1 port map( A1 => REG_8_10_port, A2 => n217_port, B1 => 
                           REG_10_10_port, B2 => n199_port, ZN => n611);
   U644 : NAND4_X1 port map( A1 => n614, A2 => n613, A3 => n612, A4 => n611, ZN
                           => n615);
   U645 : AOI22_X1 port map( A1 => n616, A2 => n85, B1 => n615, B2 => n83, ZN 
                           => n617);
   U646 : OAI221_X1 port map( B1 => n1061, B2 => n619, C1 => n1059, C2 => n618,
                           A => n617, ZN => N273);
   U647 : AOI22_X1 port map( A1 => REG_21_11_port, A2 => n110, B1 => 
                           REG_23_11_port, B2 => n92, ZN => n623);
   U648 : AOI22_X1 port map( A1 => REG_17_11_port, A2 => n146, B1 => 
                           REG_19_11_port, B2 => n128, ZN => n622);
   U649 : AOI22_X1 port map( A1 => REG_20_11_port, A2 => n182, B1 => 
                           REG_22_11_port, B2 => n164, ZN => n621);
   U650 : AOI22_X1 port map( A1 => REG_16_11_port, A2 => n218_port, B1 => 
                           REG_18_11_port, B2 => n200_port, ZN => n620);
   U651 : AND4_X1 port map( A1 => n623, A2 => n622, A3 => n621, A4 => n620, ZN 
                           => n640);
   U652 : AOI22_X1 port map( A1 => REG_29_11_port, A2 => n110, B1 => 
                           REG_31_11_port, B2 => n92, ZN => n627);
   U653 : AOI22_X1 port map( A1 => REG_25_11_port, A2 => n146, B1 => 
                           REG_27_11_port, B2 => n128, ZN => n626);
   U654 : AOI22_X1 port map( A1 => REG_28_11_port, A2 => n182, B1 => 
                           REG_30_11_port, B2 => n164, ZN => n625);
   U655 : AOI22_X1 port map( A1 => REG_24_11_port, A2 => n218_port, B1 => 
                           REG_26_11_port, B2 => n200_port, ZN => n624);
   U656 : AND4_X1 port map( A1 => n627, A2 => n626, A3 => n625, A4 => n624, ZN 
                           => n639);
   U657 : AOI22_X1 port map( A1 => REG_5_11_port, A2 => n110, B1 => 
                           REG_7_11_port, B2 => n92, ZN => n631);
   U658 : AOI22_X1 port map( A1 => REG_1_11_port, A2 => n146, B1 => 
                           REG_3_11_port, B2 => n128, ZN => n630);
   U659 : AOI22_X1 port map( A1 => REG_4_11_port, A2 => n182, B1 => 
                           REG_6_11_port, B2 => n164, ZN => n629);
   U660 : AOI22_X1 port map( A1 => REG_0_11_port, A2 => n218_port, B1 => 
                           REG_2_11_port, B2 => n200_port, ZN => n628);
   U661 : NAND4_X1 port map( A1 => n631, A2 => n630, A3 => n629, A4 => n628, ZN
                           => n637);
   U662 : AOI22_X1 port map( A1 => REG_13_11_port, A2 => n110, B1 => 
                           REG_15_11_port, B2 => n92, ZN => n635);
   U663 : AOI22_X1 port map( A1 => REG_9_11_port, A2 => n146, B1 => 
                           REG_11_11_port, B2 => n128, ZN => n634);
   U664 : AOI22_X1 port map( A1 => REG_12_11_port, A2 => n182, B1 => 
                           REG_14_11_port, B2 => n164, ZN => n633);
   U665 : AOI22_X1 port map( A1 => REG_8_11_port, A2 => n218_port, B1 => 
                           REG_10_11_port, B2 => n200_port, ZN => n632);
   U666 : NAND4_X1 port map( A1 => n635, A2 => n634, A3 => n633, A4 => n632, ZN
                           => n636);
   U667 : AOI22_X1 port map( A1 => n637, A2 => n85, B1 => n636, B2 => n83, ZN 
                           => n638);
   U668 : OAI221_X1 port map( B1 => n1061, B2 => n640, C1 => n1059, C2 => n639,
                           A => n638, ZN => N272);
   U669 : AOI22_X1 port map( A1 => REG_21_12_port, A2 => n110, B1 => 
                           REG_23_12_port, B2 => n92, ZN => n644);
   U670 : AOI22_X1 port map( A1 => REG_17_12_port, A2 => n146, B1 => 
                           REG_19_12_port, B2 => n128, ZN => n643);
   U671 : AOI22_X1 port map( A1 => REG_20_12_port, A2 => n182, B1 => 
                           REG_22_12_port, B2 => n164, ZN => n642);
   U672 : AOI22_X1 port map( A1 => REG_16_12_port, A2 => n218_port, B1 => 
                           REG_18_12_port, B2 => n200_port, ZN => n641);
   U673 : AND4_X1 port map( A1 => n644, A2 => n643, A3 => n642, A4 => n641, ZN 
                           => n661);
   U674 : AOI22_X1 port map( A1 => REG_29_12_port, A2 => n110, B1 => 
                           REG_31_12_port, B2 => n92, ZN => n648);
   U675 : AOI22_X1 port map( A1 => REG_25_12_port, A2 => n146, B1 => 
                           REG_27_12_port, B2 => n128, ZN => n647);
   U676 : AOI22_X1 port map( A1 => REG_28_12_port, A2 => n182, B1 => 
                           REG_30_12_port, B2 => n164, ZN => n646);
   U677 : AOI22_X1 port map( A1 => REG_24_12_port, A2 => n218_port, B1 => 
                           REG_26_12_port, B2 => n200_port, ZN => n645);
   U678 : AND4_X1 port map( A1 => n648, A2 => n647, A3 => n646, A4 => n645, ZN 
                           => n660);
   U679 : AOI22_X1 port map( A1 => REG_5_12_port, A2 => n110, B1 => 
                           REG_7_12_port, B2 => n92, ZN => n652);
   U680 : AOI22_X1 port map( A1 => REG_1_12_port, A2 => n146, B1 => 
                           REG_3_12_port, B2 => n128, ZN => n651);
   U681 : AOI22_X1 port map( A1 => REG_4_12_port, A2 => n182, B1 => 
                           REG_6_12_port, B2 => n164, ZN => n650);
   U682 : AOI22_X1 port map( A1 => REG_0_12_port, A2 => n218_port, B1 => 
                           REG_2_12_port, B2 => n200_port, ZN => n649);
   U683 : NAND4_X1 port map( A1 => n652, A2 => n651, A3 => n650, A4 => n649, ZN
                           => n658);
   U684 : AOI22_X1 port map( A1 => REG_13_12_port, A2 => n110, B1 => 
                           REG_15_12_port, B2 => n92, ZN => n656);
   U685 : AOI22_X1 port map( A1 => REG_9_12_port, A2 => n146, B1 => 
                           REG_11_12_port, B2 => n128, ZN => n655);
   U686 : AOI22_X1 port map( A1 => REG_12_12_port, A2 => n182, B1 => 
                           REG_14_12_port, B2 => n164, ZN => n654);
   U687 : AOI22_X1 port map( A1 => REG_8_12_port, A2 => n218_port, B1 => 
                           REG_10_12_port, B2 => n200_port, ZN => n653);
   U688 : NAND4_X1 port map( A1 => n656, A2 => n655, A3 => n654, A4 => n653, ZN
                           => n657);
   U689 : AOI22_X1 port map( A1 => n658, A2 => n85, B1 => n657, B2 => n83, ZN 
                           => n659);
   U690 : OAI221_X1 port map( B1 => n1061, B2 => n661, C1 => n1059, C2 => n660,
                           A => n659, ZN => N271);
   U691 : AOI22_X1 port map( A1 => REG_21_13_port, A2 => n110, B1 => 
                           REG_23_13_port, B2 => n92, ZN => n665);
   U692 : AOI22_X1 port map( A1 => REG_17_13_port, A2 => n146, B1 => 
                           REG_19_13_port, B2 => n128, ZN => n664);
   U693 : AOI22_X1 port map( A1 => REG_20_13_port, A2 => n182, B1 => 
                           REG_22_13_port, B2 => n164, ZN => n663);
   U694 : AOI22_X1 port map( A1 => REG_16_13_port, A2 => n218_port, B1 => 
                           REG_18_13_port, B2 => n200_port, ZN => n662);
   U695 : AND4_X1 port map( A1 => n665, A2 => n664, A3 => n663, A4 => n662, ZN 
                           => n682);
   U696 : AOI22_X1 port map( A1 => REG_29_13_port, A2 => n110, B1 => 
                           REG_31_13_port, B2 => n92, ZN => n669);
   U697 : AOI22_X1 port map( A1 => REG_25_13_port, A2 => n146, B1 => 
                           REG_27_13_port, B2 => n128, ZN => n668);
   U698 : AOI22_X1 port map( A1 => REG_28_13_port, A2 => n182, B1 => 
                           REG_30_13_port, B2 => n164, ZN => n667);
   U699 : AOI22_X1 port map( A1 => REG_24_13_port, A2 => n218_port, B1 => 
                           REG_26_13_port, B2 => n200_port, ZN => n666);
   U700 : AND4_X1 port map( A1 => n669, A2 => n668, A3 => n667, A4 => n666, ZN 
                           => n681);
   U701 : AOI22_X1 port map( A1 => REG_5_13_port, A2 => n110, B1 => 
                           REG_7_13_port, B2 => n92, ZN => n673);
   U702 : AOI22_X1 port map( A1 => REG_1_13_port, A2 => n146, B1 => 
                           REG_3_13_port, B2 => n128, ZN => n672);
   U703 : AOI22_X1 port map( A1 => REG_4_13_port, A2 => n182, B1 => 
                           REG_6_13_port, B2 => n164, ZN => n671);
   U704 : AOI22_X1 port map( A1 => REG_0_13_port, A2 => n218_port, B1 => 
                           REG_2_13_port, B2 => n200_port, ZN => n670);
   U705 : NAND4_X1 port map( A1 => n673, A2 => n672, A3 => n671, A4 => n670, ZN
                           => n679);
   U706 : AOI22_X1 port map( A1 => REG_13_13_port, A2 => n111, B1 => 
                           REG_15_13_port, B2 => n93, ZN => n677);
   U707 : AOI22_X1 port map( A1 => REG_9_13_port, A2 => n147, B1 => 
                           REG_11_13_port, B2 => n129, ZN => n676);
   U708 : AOI22_X1 port map( A1 => REG_12_13_port, A2 => n183, B1 => 
                           REG_14_13_port, B2 => n165, ZN => n675);
   U709 : AOI22_X1 port map( A1 => REG_8_13_port, A2 => n219_port, B1 => 
                           REG_10_13_port, B2 => n201_port, ZN => n674);
   U710 : NAND4_X1 port map( A1 => n677, A2 => n676, A3 => n675, A4 => n674, ZN
                           => n678);
   U711 : AOI22_X1 port map( A1 => n679, A2 => n85, B1 => n678, B2 => n83, ZN 
                           => n680);
   U712 : OAI221_X1 port map( B1 => n1061, B2 => n682, C1 => n1059, C2 => n681,
                           A => n680, ZN => N270);
   U713 : AOI22_X1 port map( A1 => REG_21_14_port, A2 => n111, B1 => 
                           REG_23_14_port, B2 => n93, ZN => n686);
   U714 : AOI22_X1 port map( A1 => REG_17_14_port, A2 => n147, B1 => 
                           REG_19_14_port, B2 => n129, ZN => n685);
   U715 : AOI22_X1 port map( A1 => REG_20_14_port, A2 => n183, B1 => 
                           REG_22_14_port, B2 => n165, ZN => n684);
   U716 : AOI22_X1 port map( A1 => REG_16_14_port, A2 => n219_port, B1 => 
                           REG_18_14_port, B2 => n201_port, ZN => n683);
   U717 : AND4_X1 port map( A1 => n686, A2 => n685, A3 => n684, A4 => n683, ZN 
                           => n703);
   U718 : AOI22_X1 port map( A1 => REG_29_14_port, A2 => n111, B1 => 
                           REG_31_14_port, B2 => n93, ZN => n690);
   U719 : AOI22_X1 port map( A1 => REG_25_14_port, A2 => n147, B1 => 
                           REG_27_14_port, B2 => n129, ZN => n689);
   U720 : AOI22_X1 port map( A1 => REG_28_14_port, A2 => n183, B1 => 
                           REG_30_14_port, B2 => n165, ZN => n688);
   U721 : AOI22_X1 port map( A1 => REG_24_14_port, A2 => n219_port, B1 => 
                           REG_26_14_port, B2 => n201_port, ZN => n687);
   U722 : AND4_X1 port map( A1 => n690, A2 => n689, A3 => n688, A4 => n687, ZN 
                           => n702);
   U723 : AOI22_X1 port map( A1 => REG_5_14_port, A2 => n111, B1 => 
                           REG_7_14_port, B2 => n93, ZN => n694);
   U724 : AOI22_X1 port map( A1 => REG_1_14_port, A2 => n147, B1 => 
                           REG_3_14_port, B2 => n129, ZN => n693);
   U725 : AOI22_X1 port map( A1 => REG_4_14_port, A2 => n183, B1 => 
                           REG_6_14_port, B2 => n165, ZN => n692);
   U726 : AOI22_X1 port map( A1 => REG_0_14_port, A2 => n219_port, B1 => 
                           REG_2_14_port, B2 => n201_port, ZN => n691);
   U727 : NAND4_X1 port map( A1 => n694, A2 => n693, A3 => n692, A4 => n691, ZN
                           => n700);
   U728 : AOI22_X1 port map( A1 => REG_13_14_port, A2 => n111, B1 => 
                           REG_15_14_port, B2 => n93, ZN => n698);
   U729 : AOI22_X1 port map( A1 => REG_9_14_port, A2 => n147, B1 => 
                           REG_11_14_port, B2 => n129, ZN => n697);
   U730 : AOI22_X1 port map( A1 => REG_12_14_port, A2 => n183, B1 => 
                           REG_14_14_port, B2 => n165, ZN => n696);
   U731 : AOI22_X1 port map( A1 => REG_8_14_port, A2 => n219_port, B1 => 
                           REG_10_14_port, B2 => n201_port, ZN => n695);
   U732 : NAND4_X1 port map( A1 => n698, A2 => n697, A3 => n696, A4 => n695, ZN
                           => n699);
   U733 : AOI22_X1 port map( A1 => n700, A2 => n85, B1 => n699, B2 => n83, ZN 
                           => n701);
   U734 : OAI221_X1 port map( B1 => n1061, B2 => n703, C1 => n1059, C2 => n702,
                           A => n701, ZN => N269);
   U735 : AOI22_X1 port map( A1 => REG_21_15_port, A2 => n111, B1 => 
                           REG_23_15_port, B2 => n93, ZN => n707);
   U736 : AOI22_X1 port map( A1 => REG_17_15_port, A2 => n147, B1 => 
                           REG_19_15_port, B2 => n129, ZN => n706);
   U737 : AOI22_X1 port map( A1 => REG_20_15_port, A2 => n183, B1 => 
                           REG_22_15_port, B2 => n165, ZN => n705);
   U738 : AOI22_X1 port map( A1 => REG_16_15_port, A2 => n219_port, B1 => 
                           REG_18_15_port, B2 => n201_port, ZN => n704);
   U739 : AND4_X1 port map( A1 => n707, A2 => n706, A3 => n705, A4 => n704, ZN 
                           => n724);
   U740 : AOI22_X1 port map( A1 => REG_29_15_port, A2 => n111, B1 => 
                           REG_31_15_port, B2 => n93, ZN => n711);
   U741 : AOI22_X1 port map( A1 => REG_25_15_port, A2 => n147, B1 => 
                           REG_27_15_port, B2 => n129, ZN => n710);
   U742 : AOI22_X1 port map( A1 => REG_28_15_port, A2 => n183, B1 => 
                           REG_30_15_port, B2 => n165, ZN => n709);
   U743 : AOI22_X1 port map( A1 => REG_24_15_port, A2 => n219_port, B1 => 
                           REG_26_15_port, B2 => n201_port, ZN => n708);
   U744 : AND4_X1 port map( A1 => n711, A2 => n710, A3 => n709, A4 => n708, ZN 
                           => n723);
   U745 : AOI22_X1 port map( A1 => REG_5_15_port, A2 => n111, B1 => 
                           REG_7_15_port, B2 => n93, ZN => n715);
   U746 : AOI22_X1 port map( A1 => REG_1_15_port, A2 => n147, B1 => 
                           REG_3_15_port, B2 => n129, ZN => n714);
   U747 : AOI22_X1 port map( A1 => REG_4_15_port, A2 => n183, B1 => 
                           REG_6_15_port, B2 => n165, ZN => n713);
   U748 : AOI22_X1 port map( A1 => REG_0_15_port, A2 => n219_port, B1 => 
                           REG_2_15_port, B2 => n201_port, ZN => n712);
   U749 : NAND4_X1 port map( A1 => n715, A2 => n714, A3 => n713, A4 => n712, ZN
                           => n721);
   U750 : AOI22_X1 port map( A1 => REG_13_15_port, A2 => n111, B1 => 
                           REG_15_15_port, B2 => n93, ZN => n719);
   U751 : AOI22_X1 port map( A1 => REG_9_15_port, A2 => n147, B1 => 
                           REG_11_15_port, B2 => n129, ZN => n718);
   U752 : AOI22_X1 port map( A1 => REG_12_15_port, A2 => n183, B1 => 
                           REG_14_15_port, B2 => n165, ZN => n717);
   U753 : AOI22_X1 port map( A1 => REG_8_15_port, A2 => n219_port, B1 => 
                           REG_10_15_port, B2 => n201_port, ZN => n716);
   U754 : NAND4_X1 port map( A1 => n719, A2 => n718, A3 => n717, A4 => n716, ZN
                           => n720);
   U755 : AOI22_X1 port map( A1 => n721, A2 => n85, B1 => n720, B2 => n83, ZN 
                           => n722);
   U756 : OAI221_X1 port map( B1 => n1061, B2 => n724, C1 => n1059, C2 => n723,
                           A => n722, ZN => N268);
   U757 : AOI22_X1 port map( A1 => REG_21_16_port, A2 => n111, B1 => 
                           REG_23_16_port, B2 => n93, ZN => n728);
   U758 : AOI22_X1 port map( A1 => REG_17_16_port, A2 => n147, B1 => 
                           REG_19_16_port, B2 => n129, ZN => n727);
   U759 : AOI22_X1 port map( A1 => REG_20_16_port, A2 => n183, B1 => 
                           REG_22_16_port, B2 => n165, ZN => n726);
   U760 : AOI22_X1 port map( A1 => REG_16_16_port, A2 => n219_port, B1 => 
                           REG_18_16_port, B2 => n201_port, ZN => n725);
   U761 : AND4_X1 port map( A1 => n728, A2 => n727, A3 => n726, A4 => n725, ZN 
                           => n745);
   U762 : AOI22_X1 port map( A1 => REG_29_16_port, A2 => n111, B1 => 
                           REG_31_16_port, B2 => n93, ZN => n732);
   U763 : AOI22_X1 port map( A1 => REG_25_16_port, A2 => n147, B1 => 
                           REG_27_16_port, B2 => n129, ZN => n731);
   U764 : AOI22_X1 port map( A1 => REG_28_16_port, A2 => n183, B1 => 
                           REG_30_16_port, B2 => n165, ZN => n730);
   U765 : AOI22_X1 port map( A1 => REG_24_16_port, A2 => n219_port, B1 => 
                           REG_26_16_port, B2 => n201_port, ZN => n729);
   U766 : AND4_X1 port map( A1 => n732, A2 => n731, A3 => n730, A4 => n729, ZN 
                           => n744);
   U767 : AOI22_X1 port map( A1 => REG_5_16_port, A2 => n112, B1 => 
                           REG_7_16_port, B2 => n94, ZN => n736);
   U768 : AOI22_X1 port map( A1 => REG_1_16_port, A2 => n148, B1 => 
                           REG_3_16_port, B2 => n130, ZN => n735);
   U769 : AOI22_X1 port map( A1 => REG_4_16_port, A2 => n184, B1 => 
                           REG_6_16_port, B2 => n166, ZN => n734);
   U770 : AOI22_X1 port map( A1 => REG_0_16_port, A2 => n220_port, B1 => 
                           REG_2_16_port, B2 => n202_port, ZN => n733);
   U771 : NAND4_X1 port map( A1 => n736, A2 => n735, A3 => n734, A4 => n733, ZN
                           => n742);
   U772 : AOI22_X1 port map( A1 => REG_13_16_port, A2 => n112, B1 => 
                           REG_15_16_port, B2 => n94, ZN => n740);
   U773 : AOI22_X1 port map( A1 => REG_9_16_port, A2 => n148, B1 => 
                           REG_11_16_port, B2 => n130, ZN => n739);
   U774 : AOI22_X1 port map( A1 => REG_12_16_port, A2 => n184, B1 => 
                           REG_14_16_port, B2 => n166, ZN => n738);
   U775 : AOI22_X1 port map( A1 => REG_8_16_port, A2 => n220_port, B1 => 
                           REG_10_16_port, B2 => n202_port, ZN => n737);
   U776 : NAND4_X1 port map( A1 => n740, A2 => n739, A3 => n738, A4 => n737, ZN
                           => n741);
   U777 : AOI22_X1 port map( A1 => n742, A2 => n85, B1 => n741, B2 => n83, ZN 
                           => n743);
   U778 : OAI221_X1 port map( B1 => n1061, B2 => n745, C1 => n1059, C2 => n744,
                           A => n743, ZN => N267);
   U779 : AOI22_X1 port map( A1 => REG_21_17_port, A2 => n112, B1 => 
                           REG_23_17_port, B2 => n94, ZN => n749);
   U780 : AOI22_X1 port map( A1 => REG_17_17_port, A2 => n148, B1 => 
                           REG_19_17_port, B2 => n130, ZN => n748);
   U781 : AOI22_X1 port map( A1 => REG_20_17_port, A2 => n184, B1 => 
                           REG_22_17_port, B2 => n166, ZN => n747);
   U782 : AOI22_X1 port map( A1 => REG_16_17_port, A2 => n220_port, B1 => 
                           REG_18_17_port, B2 => n202_port, ZN => n746);
   U783 : AND4_X1 port map( A1 => n749, A2 => n748, A3 => n747, A4 => n746, ZN 
                           => n766);
   U784 : AOI22_X1 port map( A1 => REG_29_17_port, A2 => n112, B1 => 
                           REG_31_17_port, B2 => n94, ZN => n753);
   U785 : AOI22_X1 port map( A1 => REG_25_17_port, A2 => n148, B1 => 
                           REG_27_17_port, B2 => n130, ZN => n752);
   U786 : AOI22_X1 port map( A1 => REG_28_17_port, A2 => n184, B1 => 
                           REG_30_17_port, B2 => n166, ZN => n751);
   U787 : AOI22_X1 port map( A1 => REG_24_17_port, A2 => n220_port, B1 => 
                           REG_26_17_port, B2 => n202_port, ZN => n750);
   U788 : AND4_X1 port map( A1 => n753, A2 => n752, A3 => n751, A4 => n750, ZN 
                           => n765);
   U789 : AOI22_X1 port map( A1 => REG_5_17_port, A2 => n112, B1 => 
                           REG_7_17_port, B2 => n94, ZN => n757);
   U790 : AOI22_X1 port map( A1 => REG_1_17_port, A2 => n148, B1 => 
                           REG_3_17_port, B2 => n130, ZN => n756);
   U791 : AOI22_X1 port map( A1 => REG_4_17_port, A2 => n184, B1 => 
                           REG_6_17_port, B2 => n166, ZN => n755);
   U792 : AOI22_X1 port map( A1 => REG_0_17_port, A2 => n220_port, B1 => 
                           REG_2_17_port, B2 => n202_port, ZN => n754);
   U793 : NAND4_X1 port map( A1 => n757, A2 => n756, A3 => n755, A4 => n754, ZN
                           => n763);
   U794 : AOI22_X1 port map( A1 => REG_13_17_port, A2 => n112, B1 => 
                           REG_15_17_port, B2 => n94, ZN => n761);
   U795 : AOI22_X1 port map( A1 => REG_9_17_port, A2 => n148, B1 => 
                           REG_11_17_port, B2 => n130, ZN => n760);
   U796 : AOI22_X1 port map( A1 => REG_12_17_port, A2 => n184, B1 => 
                           REG_14_17_port, B2 => n166, ZN => n759);
   U797 : AOI22_X1 port map( A1 => REG_8_17_port, A2 => n220_port, B1 => 
                           REG_10_17_port, B2 => n202_port, ZN => n758);
   U798 : NAND4_X1 port map( A1 => n761, A2 => n760, A3 => n759, A4 => n758, ZN
                           => n762);
   U799 : AOI22_X1 port map( A1 => n763, A2 => n85, B1 => n762, B2 => n83, ZN 
                           => n764);
   U800 : OAI221_X1 port map( B1 => n1061, B2 => n766, C1 => n1059, C2 => n765,
                           A => n764, ZN => N266);
   U801 : AOI22_X1 port map( A1 => REG_21_18_port, A2 => n112, B1 => 
                           REG_23_18_port, B2 => n94, ZN => n770);
   U802 : AOI22_X1 port map( A1 => REG_17_18_port, A2 => n148, B1 => 
                           REG_19_18_port, B2 => n130, ZN => n769);
   U803 : AOI22_X1 port map( A1 => REG_20_18_port, A2 => n184, B1 => 
                           REG_22_18_port, B2 => n166, ZN => n768);
   U804 : AOI22_X1 port map( A1 => REG_16_18_port, A2 => n220_port, B1 => 
                           REG_18_18_port, B2 => n202_port, ZN => n767);
   U805 : AND4_X1 port map( A1 => n770, A2 => n769, A3 => n768, A4 => n767, ZN 
                           => n787);
   U806 : AOI22_X1 port map( A1 => REG_29_18_port, A2 => n112, B1 => 
                           REG_31_18_port, B2 => n94, ZN => n774);
   U807 : AOI22_X1 port map( A1 => REG_25_18_port, A2 => n148, B1 => 
                           REG_27_18_port, B2 => n130, ZN => n773);
   U808 : AOI22_X1 port map( A1 => REG_28_18_port, A2 => n184, B1 => 
                           REG_30_18_port, B2 => n166, ZN => n772);
   U809 : AOI22_X1 port map( A1 => REG_24_18_port, A2 => n220_port, B1 => 
                           REG_26_18_port, B2 => n202_port, ZN => n771);
   U810 : AND4_X1 port map( A1 => n774, A2 => n773, A3 => n772, A4 => n771, ZN 
                           => n786);
   U811 : AOI22_X1 port map( A1 => REG_5_18_port, A2 => n112, B1 => 
                           REG_7_18_port, B2 => n94, ZN => n778);
   U812 : AOI22_X1 port map( A1 => REG_1_18_port, A2 => n148, B1 => 
                           REG_3_18_port, B2 => n130, ZN => n777);
   U813 : AOI22_X1 port map( A1 => REG_4_18_port, A2 => n184, B1 => 
                           REG_6_18_port, B2 => n166, ZN => n776);
   U814 : AOI22_X1 port map( A1 => REG_0_18_port, A2 => n220_port, B1 => 
                           REG_2_18_port, B2 => n202_port, ZN => n775);
   U815 : NAND4_X1 port map( A1 => n778, A2 => n777, A3 => n776, A4 => n775, ZN
                           => n784);
   U816 : AOI22_X1 port map( A1 => REG_13_18_port, A2 => n112, B1 => 
                           REG_15_18_port, B2 => n94, ZN => n782);
   U817 : AOI22_X1 port map( A1 => REG_9_18_port, A2 => n148, B1 => 
                           REG_11_18_port, B2 => n130, ZN => n781);
   U818 : AOI22_X1 port map( A1 => REG_12_18_port, A2 => n184, B1 => 
                           REG_14_18_port, B2 => n166, ZN => n780);
   U819 : AOI22_X1 port map( A1 => REG_8_18_port, A2 => n220_port, B1 => 
                           REG_10_18_port, B2 => n202_port, ZN => n779);
   U820 : NAND4_X1 port map( A1 => n782, A2 => n781, A3 => n780, A4 => n779, ZN
                           => n783);
   U821 : AOI22_X1 port map( A1 => n784, A2 => n85, B1 => n783, B2 => n83, ZN 
                           => n785);
   U822 : OAI221_X1 port map( B1 => n1061, B2 => n787, C1 => n1059, C2 => n786,
                           A => n785, ZN => N265);
   U823 : AOI22_X1 port map( A1 => REG_21_19_port, A2 => n112, B1 => 
                           REG_23_19_port, B2 => n94, ZN => n791);
   U824 : AOI22_X1 port map( A1 => REG_17_19_port, A2 => n148, B1 => 
                           REG_19_19_port, B2 => n130, ZN => n790);
   U825 : AOI22_X1 port map( A1 => REG_20_19_port, A2 => n184, B1 => 
                           REG_22_19_port, B2 => n166, ZN => n789);
   U826 : AOI22_X1 port map( A1 => REG_16_19_port, A2 => n220_port, B1 => 
                           REG_18_19_port, B2 => n202_port, ZN => n788);
   U827 : AND4_X1 port map( A1 => n791, A2 => n790, A3 => n789, A4 => n788, ZN 
                           => n808);
   U828 : AOI22_X1 port map( A1 => REG_29_19_port, A2 => n113, B1 => 
                           REG_31_19_port, B2 => n95, ZN => n795);
   U829 : AOI22_X1 port map( A1 => REG_25_19_port, A2 => n149, B1 => 
                           REG_27_19_port, B2 => n131, ZN => n794);
   U830 : AOI22_X1 port map( A1 => REG_28_19_port, A2 => n185, B1 => 
                           REG_30_19_port, B2 => n167, ZN => n793);
   U831 : AOI22_X1 port map( A1 => REG_24_19_port, A2 => n221_port, B1 => 
                           REG_26_19_port, B2 => n203_port, ZN => n792);
   U832 : AND4_X1 port map( A1 => n795, A2 => n794, A3 => n793, A4 => n792, ZN 
                           => n807);
   U833 : AOI22_X1 port map( A1 => REG_5_19_port, A2 => n113, B1 => 
                           REG_7_19_port, B2 => n95, ZN => n799);
   U834 : AOI22_X1 port map( A1 => REG_1_19_port, A2 => n149, B1 => 
                           REG_3_19_port, B2 => n131, ZN => n798);
   U835 : AOI22_X1 port map( A1 => REG_4_19_port, A2 => n185, B1 => 
                           REG_6_19_port, B2 => n167, ZN => n797);
   U836 : AOI22_X1 port map( A1 => REG_0_19_port, A2 => n221_port, B1 => 
                           REG_2_19_port, B2 => n203_port, ZN => n796);
   U837 : NAND4_X1 port map( A1 => n799, A2 => n798, A3 => n797, A4 => n796, ZN
                           => n805);
   U838 : AOI22_X1 port map( A1 => REG_13_19_port, A2 => n113, B1 => 
                           REG_15_19_port, B2 => n95, ZN => n803);
   U839 : AOI22_X1 port map( A1 => REG_9_19_port, A2 => n149, B1 => 
                           REG_11_19_port, B2 => n131, ZN => n802);
   U840 : AOI22_X1 port map( A1 => REG_12_19_port, A2 => n185, B1 => 
                           REG_14_19_port, B2 => n167, ZN => n801);
   U841 : AOI22_X1 port map( A1 => REG_8_19_port, A2 => n221_port, B1 => 
                           REG_10_19_port, B2 => n203_port, ZN => n800);
   U842 : NAND4_X1 port map( A1 => n803, A2 => n802, A3 => n801, A4 => n800, ZN
                           => n804);
   U843 : AOI22_X1 port map( A1 => n805, A2 => n85, B1 => n804, B2 => n83, ZN 
                           => n806);
   U844 : OAI221_X1 port map( B1 => n1061, B2 => n808, C1 => n1059, C2 => n807,
                           A => n806, ZN => N264);
   U845 : AOI22_X1 port map( A1 => REG_21_20_port, A2 => n113, B1 => 
                           REG_23_20_port, B2 => n95, ZN => n812);
   U846 : AOI22_X1 port map( A1 => REG_17_20_port, A2 => n149, B1 => 
                           REG_19_20_port, B2 => n131, ZN => n811);
   U847 : AOI22_X1 port map( A1 => REG_20_20_port, A2 => n185, B1 => 
                           REG_22_20_port, B2 => n167, ZN => n810);
   U848 : AOI22_X1 port map( A1 => REG_16_20_port, A2 => n221_port, B1 => 
                           REG_18_20_port, B2 => n203_port, ZN => n809);
   U849 : AND4_X1 port map( A1 => n812, A2 => n811, A3 => n810, A4 => n809, ZN 
                           => n829);
   U850 : AOI22_X1 port map( A1 => REG_29_20_port, A2 => n113, B1 => 
                           REG_31_20_port, B2 => n95, ZN => n816);
   U851 : AOI22_X1 port map( A1 => REG_25_20_port, A2 => n149, B1 => 
                           REG_27_20_port, B2 => n131, ZN => n815);
   U852 : AOI22_X1 port map( A1 => REG_28_20_port, A2 => n185, B1 => 
                           REG_30_20_port, B2 => n167, ZN => n814);
   U853 : AOI22_X1 port map( A1 => REG_24_20_port, A2 => n221_port, B1 => 
                           REG_26_20_port, B2 => n203_port, ZN => n813);
   U854 : AND4_X1 port map( A1 => n816, A2 => n815, A3 => n814, A4 => n813, ZN 
                           => n828);
   U855 : AOI22_X1 port map( A1 => REG_5_20_port, A2 => n113, B1 => 
                           REG_7_20_port, B2 => n95, ZN => n820);
   U856 : AOI22_X1 port map( A1 => REG_1_20_port, A2 => n149, B1 => 
                           REG_3_20_port, B2 => n131, ZN => n819);
   U857 : AOI22_X1 port map( A1 => REG_4_20_port, A2 => n185, B1 => 
                           REG_6_20_port, B2 => n167, ZN => n818);
   U858 : AOI22_X1 port map( A1 => REG_0_20_port, A2 => n221_port, B1 => 
                           REG_2_20_port, B2 => n203_port, ZN => n817);
   U859 : NAND4_X1 port map( A1 => n820, A2 => n819, A3 => n818, A4 => n817, ZN
                           => n826);
   U860 : AOI22_X1 port map( A1 => REG_13_20_port, A2 => n113, B1 => 
                           REG_15_20_port, B2 => n95, ZN => n824);
   U861 : AOI22_X1 port map( A1 => REG_9_20_port, A2 => n149, B1 => 
                           REG_11_20_port, B2 => n131, ZN => n823);
   U862 : AOI22_X1 port map( A1 => REG_12_20_port, A2 => n185, B1 => 
                           REG_14_20_port, B2 => n167, ZN => n822);
   U863 : AOI22_X1 port map( A1 => REG_8_20_port, A2 => n221_port, B1 => 
                           REG_10_20_port, B2 => n203_port, ZN => n821);
   U864 : NAND4_X1 port map( A1 => n824, A2 => n823, A3 => n822, A4 => n821, ZN
                           => n825);
   U865 : AOI22_X1 port map( A1 => n826, A2 => n85, B1 => n825, B2 => n83, ZN 
                           => n827);
   U866 : OAI221_X1 port map( B1 => n1061, B2 => n829, C1 => n1059, C2 => n828,
                           A => n827, ZN => N263);
   U867 : AOI22_X1 port map( A1 => REG_21_21_port, A2 => n113, B1 => 
                           REG_23_21_port, B2 => n95, ZN => n833);
   U868 : AOI22_X1 port map( A1 => REG_17_21_port, A2 => n149, B1 => 
                           REG_19_21_port, B2 => n131, ZN => n832);
   U869 : AOI22_X1 port map( A1 => REG_20_21_port, A2 => n185, B1 => 
                           REG_22_21_port, B2 => n167, ZN => n831);
   U870 : AOI22_X1 port map( A1 => REG_16_21_port, A2 => n221_port, B1 => 
                           REG_18_21_port, B2 => n203_port, ZN => n830);
   U871 : AND4_X1 port map( A1 => n833, A2 => n832, A3 => n831, A4 => n830, ZN 
                           => n850);
   U872 : AOI22_X1 port map( A1 => REG_29_21_port, A2 => n113, B1 => 
                           REG_31_21_port, B2 => n95, ZN => n837);
   U873 : AOI22_X1 port map( A1 => REG_25_21_port, A2 => n149, B1 => 
                           REG_27_21_port, B2 => n131, ZN => n836);
   U874 : AOI22_X1 port map( A1 => REG_28_21_port, A2 => n185, B1 => 
                           REG_30_21_port, B2 => n167, ZN => n835);
   U875 : AOI22_X1 port map( A1 => REG_24_21_port, A2 => n221_port, B1 => 
                           REG_26_21_port, B2 => n203_port, ZN => n834);
   U876 : AND4_X1 port map( A1 => n837, A2 => n836, A3 => n835, A4 => n834, ZN 
                           => n849);
   U877 : AOI22_X1 port map( A1 => REG_5_21_port, A2 => n113, B1 => 
                           REG_7_21_port, B2 => n95, ZN => n841);
   U878 : AOI22_X1 port map( A1 => REG_1_21_port, A2 => n149, B1 => 
                           REG_3_21_port, B2 => n131, ZN => n840);
   U879 : AOI22_X1 port map( A1 => REG_4_21_port, A2 => n185, B1 => 
                           REG_6_21_port, B2 => n167, ZN => n839);
   U880 : AOI22_X1 port map( A1 => REG_0_21_port, A2 => n221_port, B1 => 
                           REG_2_21_port, B2 => n203_port, ZN => n838);
   U881 : NAND4_X1 port map( A1 => n841, A2 => n840, A3 => n839, A4 => n838, ZN
                           => n847);
   U882 : AOI22_X1 port map( A1 => REG_13_21_port, A2 => n113, B1 => 
                           REG_15_21_port, B2 => n95, ZN => n845);
   U883 : AOI22_X1 port map( A1 => REG_9_21_port, A2 => n149, B1 => 
                           REG_11_21_port, B2 => n131, ZN => n844);
   U884 : AOI22_X1 port map( A1 => REG_12_21_port, A2 => n185, B1 => 
                           REG_14_21_port, B2 => n167, ZN => n843);
   U885 : AOI22_X1 port map( A1 => REG_8_21_port, A2 => n221_port, B1 => 
                           REG_10_21_port, B2 => n203_port, ZN => n842);
   U886 : NAND4_X1 port map( A1 => n845, A2 => n844, A3 => n843, A4 => n842, ZN
                           => n846);
   U887 : AOI22_X1 port map( A1 => n847, A2 => n85, B1 => n846, B2 => n83, ZN 
                           => n848);
   U888 : OAI221_X1 port map( B1 => n1061, B2 => n850, C1 => n1059, C2 => n849,
                           A => n848, ZN => N262);
   U889 : AOI22_X1 port map( A1 => REG_21_22_port, A2 => n114, B1 => 
                           REG_23_22_port, B2 => n96, ZN => n854);
   U890 : AOI22_X1 port map( A1 => REG_17_22_port, A2 => n150, B1 => 
                           REG_19_22_port, B2 => n132, ZN => n853);
   U891 : AOI22_X1 port map( A1 => REG_20_22_port, A2 => n186, B1 => 
                           REG_22_22_port, B2 => n168, ZN => n852);
   U892 : AOI22_X1 port map( A1 => REG_16_22_port, A2 => n222_port, B1 => 
                           REG_18_22_port, B2 => n204_port, ZN => n851);
   U893 : AND4_X1 port map( A1 => n854, A2 => n853, A3 => n852, A4 => n851, ZN 
                           => n871);
   U894 : AOI22_X1 port map( A1 => REG_29_22_port, A2 => n114, B1 => 
                           REG_31_22_port, B2 => n96, ZN => n858);
   U895 : AOI22_X1 port map( A1 => REG_25_22_port, A2 => n150, B1 => 
                           REG_27_22_port, B2 => n132, ZN => n857);
   U896 : AOI22_X1 port map( A1 => REG_28_22_port, A2 => n186, B1 => 
                           REG_30_22_port, B2 => n168, ZN => n856);
   U897 : AOI22_X1 port map( A1 => REG_24_22_port, A2 => n222_port, B1 => 
                           REG_26_22_port, B2 => n204_port, ZN => n855);
   U898 : AND4_X1 port map( A1 => n858, A2 => n857, A3 => n856, A4 => n855, ZN 
                           => n870);
   U899 : AOI22_X1 port map( A1 => REG_5_22_port, A2 => n114, B1 => 
                           REG_7_22_port, B2 => n96, ZN => n862);
   U900 : AOI22_X1 port map( A1 => REG_1_22_port, A2 => n150, B1 => 
                           REG_3_22_port, B2 => n132, ZN => n861);
   U901 : AOI22_X1 port map( A1 => REG_4_22_port, A2 => n186, B1 => 
                           REG_6_22_port, B2 => n168, ZN => n860);
   U902 : AOI22_X1 port map( A1 => REG_0_22_port, A2 => n222_port, B1 => 
                           REG_2_22_port, B2 => n204_port, ZN => n859);
   U903 : NAND4_X1 port map( A1 => n862, A2 => n861, A3 => n860, A4 => n859, ZN
                           => n868);
   U904 : AOI22_X1 port map( A1 => REG_13_22_port, A2 => n114, B1 => 
                           REG_15_22_port, B2 => n96, ZN => n866);
   U905 : AOI22_X1 port map( A1 => REG_9_22_port, A2 => n150, B1 => 
                           REG_11_22_port, B2 => n132, ZN => n865);
   U906 : AOI22_X1 port map( A1 => REG_12_22_port, A2 => n186, B1 => 
                           REG_14_22_port, B2 => n168, ZN => n864);
   U907 : AOI22_X1 port map( A1 => REG_8_22_port, A2 => n222_port, B1 => 
                           REG_10_22_port, B2 => n204_port, ZN => n863);
   U908 : NAND4_X1 port map( A1 => n866, A2 => n865, A3 => n864, A4 => n863, ZN
                           => n867);
   U909 : AOI22_X1 port map( A1 => n868, A2 => n85, B1 => n867, B2 => n83, ZN 
                           => n869);
   U910 : OAI221_X1 port map( B1 => n1061, B2 => n871, C1 => n1059, C2 => n870,
                           A => n869, ZN => N261);
   U911 : AOI22_X1 port map( A1 => REG_21_23_port, A2 => n114, B1 => 
                           REG_23_23_port, B2 => n96, ZN => n875);
   U912 : AOI22_X1 port map( A1 => REG_17_23_port, A2 => n150, B1 => 
                           REG_19_23_port, B2 => n132, ZN => n874);
   U913 : AOI22_X1 port map( A1 => REG_20_23_port, A2 => n186, B1 => 
                           REG_22_23_port, B2 => n168, ZN => n873);
   U914 : AOI22_X1 port map( A1 => REG_16_23_port, A2 => n222_port, B1 => 
                           REG_18_23_port, B2 => n204_port, ZN => n872);
   U915 : AND4_X1 port map( A1 => n875, A2 => n874, A3 => n873, A4 => n872, ZN 
                           => n892);
   U916 : AOI22_X1 port map( A1 => REG_29_23_port, A2 => n114, B1 => 
                           REG_31_23_port, B2 => n96, ZN => n879);
   U917 : AOI22_X1 port map( A1 => REG_25_23_port, A2 => n150, B1 => 
                           REG_27_23_port, B2 => n132, ZN => n878);
   U918 : AOI22_X1 port map( A1 => REG_28_23_port, A2 => n186, B1 => 
                           REG_30_23_port, B2 => n168, ZN => n877);
   U919 : AOI22_X1 port map( A1 => REG_24_23_port, A2 => n222_port, B1 => 
                           REG_26_23_port, B2 => n204_port, ZN => n876);
   U920 : AND4_X1 port map( A1 => n879, A2 => n878, A3 => n877, A4 => n876, ZN 
                           => n891);
   U921 : AOI22_X1 port map( A1 => REG_5_23_port, A2 => n114, B1 => 
                           REG_7_23_port, B2 => n96, ZN => n883);
   U922 : AOI22_X1 port map( A1 => REG_1_23_port, A2 => n150, B1 => 
                           REG_3_23_port, B2 => n132, ZN => n882);
   U923 : AOI22_X1 port map( A1 => REG_4_23_port, A2 => n186, B1 => 
                           REG_6_23_port, B2 => n168, ZN => n881);
   U924 : AOI22_X1 port map( A1 => REG_0_23_port, A2 => n222_port, B1 => 
                           REG_2_23_port, B2 => n204_port, ZN => n880);
   U925 : NAND4_X1 port map( A1 => n883, A2 => n882, A3 => n881, A4 => n880, ZN
                           => n889);
   U926 : AOI22_X1 port map( A1 => REG_13_23_port, A2 => n114, B1 => 
                           REG_15_23_port, B2 => n96, ZN => n887);
   U927 : AOI22_X1 port map( A1 => REG_9_23_port, A2 => n150, B1 => 
                           REG_11_23_port, B2 => n132, ZN => n886);
   U928 : AOI22_X1 port map( A1 => REG_12_23_port, A2 => n186, B1 => 
                           REG_14_23_port, B2 => n168, ZN => n885);
   U929 : AOI22_X1 port map( A1 => REG_8_23_port, A2 => n222_port, B1 => 
                           REG_10_23_port, B2 => n204_port, ZN => n884);
   U930 : NAND4_X1 port map( A1 => n887, A2 => n886, A3 => n885, A4 => n884, ZN
                           => n888);
   U931 : AOI22_X1 port map( A1 => n889, A2 => n85, B1 => n888, B2 => n83, ZN 
                           => n890);
   U932 : OAI221_X1 port map( B1 => n1061, B2 => n892, C1 => n1059, C2 => n891,
                           A => n890, ZN => N260);
   U933 : AOI22_X1 port map( A1 => REG_21_24_port, A2 => n114, B1 => 
                           REG_23_24_port, B2 => n96, ZN => n896);
   U934 : AOI22_X1 port map( A1 => REG_17_24_port, A2 => n150, B1 => 
                           REG_19_24_port, B2 => n132, ZN => n895);
   U935 : AOI22_X1 port map( A1 => REG_20_24_port, A2 => n186, B1 => 
                           REG_22_24_port, B2 => n168, ZN => n894);
   U936 : AOI22_X1 port map( A1 => REG_16_24_port, A2 => n222_port, B1 => 
                           REG_18_24_port, B2 => n204_port, ZN => n893);
   U937 : AND4_X1 port map( A1 => n896, A2 => n895, A3 => n894, A4 => n893, ZN 
                           => n913);
   U938 : AOI22_X1 port map( A1 => REG_29_24_port, A2 => n114, B1 => 
                           REG_31_24_port, B2 => n96, ZN => n900);
   U939 : AOI22_X1 port map( A1 => REG_25_24_port, A2 => n150, B1 => 
                           REG_27_24_port, B2 => n132, ZN => n899);
   U940 : AOI22_X1 port map( A1 => REG_28_24_port, A2 => n186, B1 => 
                           REG_30_24_port, B2 => n168, ZN => n898);
   U941 : AOI22_X1 port map( A1 => REG_24_24_port, A2 => n222_port, B1 => 
                           REG_26_24_port, B2 => n204_port, ZN => n897);
   U942 : AND4_X1 port map( A1 => n900, A2 => n899, A3 => n898, A4 => n897, ZN 
                           => n912);
   U943 : AOI22_X1 port map( A1 => REG_5_24_port, A2 => n114, B1 => 
                           REG_7_24_port, B2 => n96, ZN => n904);
   U944 : AOI22_X1 port map( A1 => REG_1_24_port, A2 => n150, B1 => 
                           REG_3_24_port, B2 => n132, ZN => n903);
   U945 : AOI22_X1 port map( A1 => REG_4_24_port, A2 => n186, B1 => 
                           REG_6_24_port, B2 => n168, ZN => n902);
   U946 : AOI22_X1 port map( A1 => REG_0_24_port, A2 => n222_port, B1 => 
                           REG_2_24_port, B2 => n204_port, ZN => n901);
   U947 : NAND4_X1 port map( A1 => n904, A2 => n903, A3 => n902, A4 => n901, ZN
                           => n910);
   U948 : AOI22_X1 port map( A1 => REG_13_24_port, A2 => n115, B1 => 
                           REG_15_24_port, B2 => n97, ZN => n908);
   U949 : AOI22_X1 port map( A1 => REG_9_24_port, A2 => n151, B1 => 
                           REG_11_24_port, B2 => n133, ZN => n907);
   U950 : AOI22_X1 port map( A1 => REG_12_24_port, A2 => n187, B1 => 
                           REG_14_24_port, B2 => n169, ZN => n906);
   U951 : AOI22_X1 port map( A1 => REG_8_24_port, A2 => n223_port, B1 => 
                           REG_10_24_port, B2 => n205_port, ZN => n905);
   U952 : NAND4_X1 port map( A1 => n908, A2 => n907, A3 => n906, A4 => n905, ZN
                           => n909);
   U953 : AOI22_X1 port map( A1 => n910, A2 => n85, B1 => n909, B2 => n83, ZN 
                           => n911);
   U954 : OAI221_X1 port map( B1 => n1061, B2 => n913, C1 => n1059, C2 => n912,
                           A => n911, ZN => N259);
   U955 : AOI22_X1 port map( A1 => REG_21_25_port, A2 => n115, B1 => 
                           REG_23_25_port, B2 => n97, ZN => n917);
   U956 : AOI22_X1 port map( A1 => REG_17_25_port, A2 => n151, B1 => 
                           REG_19_25_port, B2 => n133, ZN => n916);
   U957 : AOI22_X1 port map( A1 => REG_20_25_port, A2 => n187, B1 => 
                           REG_22_25_port, B2 => n169, ZN => n915);
   U958 : AOI22_X1 port map( A1 => REG_16_25_port, A2 => n223_port, B1 => 
                           REG_18_25_port, B2 => n205_port, ZN => n914);
   U959 : AND4_X1 port map( A1 => n917, A2 => n916, A3 => n915, A4 => n914, ZN 
                           => n934);
   U960 : AOI22_X1 port map( A1 => REG_29_25_port, A2 => n115, B1 => 
                           REG_31_25_port, B2 => n97, ZN => n921);
   U961 : AOI22_X1 port map( A1 => REG_25_25_port, A2 => n151, B1 => 
                           REG_27_25_port, B2 => n133, ZN => n920);
   U962 : AOI22_X1 port map( A1 => REG_28_25_port, A2 => n187, B1 => 
                           REG_30_25_port, B2 => n169, ZN => n919);
   U963 : AOI22_X1 port map( A1 => REG_24_25_port, A2 => n223_port, B1 => 
                           REG_26_25_port, B2 => n205_port, ZN => n918);
   U964 : AND4_X1 port map( A1 => n921, A2 => n920, A3 => n919, A4 => n918, ZN 
                           => n933);
   U965 : AOI22_X1 port map( A1 => REG_5_25_port, A2 => n115, B1 => 
                           REG_7_25_port, B2 => n97, ZN => n925);
   U966 : AOI22_X1 port map( A1 => REG_1_25_port, A2 => n151, B1 => 
                           REG_3_25_port, B2 => n133, ZN => n924);
   U967 : AOI22_X1 port map( A1 => REG_4_25_port, A2 => n187, B1 => 
                           REG_6_25_port, B2 => n169, ZN => n923);
   U968 : AOI22_X1 port map( A1 => REG_0_25_port, A2 => n223_port, B1 => 
                           REG_2_25_port, B2 => n205_port, ZN => n922);
   U969 : NAND4_X1 port map( A1 => n925, A2 => n924, A3 => n923, A4 => n922, ZN
                           => n931);
   U970 : AOI22_X1 port map( A1 => REG_13_25_port, A2 => n115, B1 => 
                           REG_15_25_port, B2 => n97, ZN => n929);
   U971 : AOI22_X1 port map( A1 => REG_9_25_port, A2 => n151, B1 => 
                           REG_11_25_port, B2 => n133, ZN => n928);
   U972 : AOI22_X1 port map( A1 => REG_12_25_port, A2 => n187, B1 => 
                           REG_14_25_port, B2 => n169, ZN => n927);
   U973 : AOI22_X1 port map( A1 => REG_8_25_port, A2 => n223_port, B1 => 
                           REG_10_25_port, B2 => n205_port, ZN => n926);
   U974 : NAND4_X1 port map( A1 => n929, A2 => n928, A3 => n927, A4 => n926, ZN
                           => n930);
   U975 : AOI22_X1 port map( A1 => n931, A2 => n85, B1 => n930, B2 => n83, ZN 
                           => n932);
   U976 : OAI221_X1 port map( B1 => n1061, B2 => n934, C1 => n1059, C2 => n933,
                           A => n932, ZN => N258);
   U977 : AOI22_X1 port map( A1 => REG_21_26_port, A2 => n115, B1 => 
                           REG_23_26_port, B2 => n97, ZN => n938);
   U978 : AOI22_X1 port map( A1 => REG_17_26_port, A2 => n151, B1 => 
                           REG_19_26_port, B2 => n133, ZN => n937);
   U979 : AOI22_X1 port map( A1 => REG_20_26_port, A2 => n187, B1 => 
                           REG_22_26_port, B2 => n169, ZN => n936);
   U980 : AOI22_X1 port map( A1 => REG_16_26_port, A2 => n223_port, B1 => 
                           REG_18_26_port, B2 => n205_port, ZN => n935);
   U981 : AND4_X1 port map( A1 => n938, A2 => n937, A3 => n936, A4 => n935, ZN 
                           => n955);
   U982 : AOI22_X1 port map( A1 => REG_29_26_port, A2 => n115, B1 => 
                           REG_31_26_port, B2 => n97, ZN => n942);
   U983 : AOI22_X1 port map( A1 => REG_25_26_port, A2 => n151, B1 => 
                           REG_27_26_port, B2 => n133, ZN => n941);
   U984 : AOI22_X1 port map( A1 => REG_28_26_port, A2 => n187, B1 => 
                           REG_30_26_port, B2 => n169, ZN => n940);
   U985 : AOI22_X1 port map( A1 => REG_24_26_port, A2 => n223_port, B1 => 
                           REG_26_26_port, B2 => n205_port, ZN => n939);
   U986 : AND4_X1 port map( A1 => n942, A2 => n941, A3 => n940, A4 => n939, ZN 
                           => n954);
   U987 : AOI22_X1 port map( A1 => REG_5_26_port, A2 => n115, B1 => 
                           REG_7_26_port, B2 => n97, ZN => n946);
   U988 : AOI22_X1 port map( A1 => REG_1_26_port, A2 => n151, B1 => 
                           REG_3_26_port, B2 => n133, ZN => n945);
   U989 : AOI22_X1 port map( A1 => REG_4_26_port, A2 => n187, B1 => 
                           REG_6_26_port, B2 => n169, ZN => n944);
   U990 : AOI22_X1 port map( A1 => REG_0_26_port, A2 => n223_port, B1 => 
                           REG_2_26_port, B2 => n205_port, ZN => n943);
   U991 : NAND4_X1 port map( A1 => n946, A2 => n945, A3 => n944, A4 => n943, ZN
                           => n952);
   U992 : AOI22_X1 port map( A1 => REG_13_26_port, A2 => n115, B1 => 
                           REG_15_26_port, B2 => n97, ZN => n950);
   U993 : AOI22_X1 port map( A1 => REG_9_26_port, A2 => n151, B1 => 
                           REG_11_26_port, B2 => n133, ZN => n949);
   U994 : AOI22_X1 port map( A1 => REG_12_26_port, A2 => n187, B1 => 
                           REG_14_26_port, B2 => n169, ZN => n948);
   U995 : AOI22_X1 port map( A1 => REG_8_26_port, A2 => n223_port, B1 => 
                           REG_10_26_port, B2 => n205_port, ZN => n947);
   U996 : NAND4_X1 port map( A1 => n950, A2 => n949, A3 => n948, A4 => n947, ZN
                           => n951);
   U997 : AOI22_X1 port map( A1 => n952, A2 => n85, B1 => n951, B2 => n83, ZN 
                           => n953);
   U998 : OAI221_X1 port map( B1 => n1061, B2 => n955, C1 => n1059, C2 => n954,
                           A => n953, ZN => N257);
   U999 : AOI22_X1 port map( A1 => REG_21_27_port, A2 => n115, B1 => 
                           REG_23_27_port, B2 => n97, ZN => n959);
   U1000 : AOI22_X1 port map( A1 => REG_17_27_port, A2 => n151, B1 => 
                           REG_19_27_port, B2 => n133, ZN => n958);
   U1001 : AOI22_X1 port map( A1 => REG_20_27_port, A2 => n187, B1 => 
                           REG_22_27_port, B2 => n169, ZN => n957);
   U1002 : AOI22_X1 port map( A1 => REG_16_27_port, A2 => n223_port, B1 => 
                           REG_18_27_port, B2 => n205_port, ZN => n956);
   U1003 : AND4_X1 port map( A1 => n959, A2 => n958, A3 => n957, A4 => n956, ZN
                           => n976);
   U1004 : AOI22_X1 port map( A1 => REG_29_27_port, A2 => n115, B1 => 
                           REG_31_27_port, B2 => n97, ZN => n963);
   U1005 : AOI22_X1 port map( A1 => REG_25_27_port, A2 => n151, B1 => 
                           REG_27_27_port, B2 => n133, ZN => n962);
   U1006 : AOI22_X1 port map( A1 => REG_28_27_port, A2 => n187, B1 => 
                           REG_30_27_port, B2 => n169, ZN => n961);
   U1007 : AOI22_X1 port map( A1 => REG_24_27_port, A2 => n223_port, B1 => 
                           REG_26_27_port, B2 => n205_port, ZN => n960);
   U1008 : AND4_X1 port map( A1 => n963, A2 => n962, A3 => n961, A4 => n960, ZN
                           => n975);
   U1009 : AOI22_X1 port map( A1 => REG_5_27_port, A2 => n116, B1 => 
                           REG_7_27_port, B2 => n98, ZN => n967);
   U1010 : AOI22_X1 port map( A1 => REG_1_27_port, A2 => n152, B1 => 
                           REG_3_27_port, B2 => n134, ZN => n966);
   U1011 : AOI22_X1 port map( A1 => REG_4_27_port, A2 => n188_port, B1 => 
                           REG_6_27_port, B2 => n170, ZN => n965);
   U1012 : AOI22_X1 port map( A1 => REG_0_27_port, A2 => n224_port, B1 => 
                           REG_2_27_port, B2 => n206_port, ZN => n964);
   U1013 : NAND4_X1 port map( A1 => n967, A2 => n966, A3 => n965, A4 => n964, 
                           ZN => n973);
   U1014 : AOI22_X1 port map( A1 => REG_13_27_port, A2 => n116, B1 => 
                           REG_15_27_port, B2 => n98, ZN => n971);
   U1015 : AOI22_X1 port map( A1 => REG_9_27_port, A2 => n152, B1 => 
                           REG_11_27_port, B2 => n134, ZN => n970);
   U1016 : AOI22_X1 port map( A1 => REG_12_27_port, A2 => n188_port, B1 => 
                           REG_14_27_port, B2 => n170, ZN => n969);
   U1017 : AOI22_X1 port map( A1 => REG_8_27_port, A2 => n224_port, B1 => 
                           REG_10_27_port, B2 => n206_port, ZN => n968);
   U1018 : NAND4_X1 port map( A1 => n971, A2 => n970, A3 => n969, A4 => n968, 
                           ZN => n972);
   U1019 : AOI22_X1 port map( A1 => n973, A2 => n85, B1 => n972, B2 => n83, ZN 
                           => n974);
   U1020 : OAI221_X1 port map( B1 => n1061, B2 => n976, C1 => n1059, C2 => n975
                           , A => n974, ZN => N256);
   U1021 : AOI22_X1 port map( A1 => REG_21_28_port, A2 => n116, B1 => 
                           REG_23_28_port, B2 => n98, ZN => n980);
   U1022 : AOI22_X1 port map( A1 => REG_17_28_port, A2 => n152, B1 => 
                           REG_19_28_port, B2 => n134, ZN => n979);
   U1023 : AOI22_X1 port map( A1 => REG_20_28_port, A2 => n188_port, B1 => 
                           REG_22_28_port, B2 => n170, ZN => n978);
   U1024 : AOI22_X1 port map( A1 => REG_16_28_port, A2 => n224_port, B1 => 
                           REG_18_28_port, B2 => n206_port, ZN => n977);
   U1025 : AND4_X1 port map( A1 => n980, A2 => n979, A3 => n978, A4 => n977, ZN
                           => n997);
   U1026 : AOI22_X1 port map( A1 => REG_29_28_port, A2 => n116, B1 => 
                           REG_31_28_port, B2 => n98, ZN => n984);
   U1027 : AOI22_X1 port map( A1 => REG_25_28_port, A2 => n152, B1 => 
                           REG_27_28_port, B2 => n134, ZN => n983);
   U1028 : AOI22_X1 port map( A1 => REG_28_28_port, A2 => n188_port, B1 => 
                           REG_30_28_port, B2 => n170, ZN => n982);
   U1029 : AOI22_X1 port map( A1 => REG_24_28_port, A2 => n224_port, B1 => 
                           REG_26_28_port, B2 => n206_port, ZN => n981);
   U1030 : AND4_X1 port map( A1 => n984, A2 => n983, A3 => n982, A4 => n981, ZN
                           => n996);
   U1031 : AOI22_X1 port map( A1 => REG_5_28_port, A2 => n116, B1 => 
                           REG_7_28_port, B2 => n98, ZN => n988);
   U1032 : AOI22_X1 port map( A1 => REG_1_28_port, A2 => n152, B1 => 
                           REG_3_28_port, B2 => n134, ZN => n987);
   U1033 : AOI22_X1 port map( A1 => REG_4_28_port, A2 => n188_port, B1 => 
                           REG_6_28_port, B2 => n170, ZN => n986);
   U1034 : AOI22_X1 port map( A1 => REG_0_28_port, A2 => n224_port, B1 => 
                           REG_2_28_port, B2 => n206_port, ZN => n985);
   U1035 : NAND4_X1 port map( A1 => n988, A2 => n987, A3 => n986, A4 => n985, 
                           ZN => n994);
   U1036 : AOI22_X1 port map( A1 => REG_13_28_port, A2 => n116, B1 => 
                           REG_15_28_port, B2 => n98, ZN => n992);
   U1037 : AOI22_X1 port map( A1 => REG_9_28_port, A2 => n152, B1 => 
                           REG_11_28_port, B2 => n134, ZN => n991);
   U1038 : AOI22_X1 port map( A1 => REG_12_28_port, A2 => n188_port, B1 => 
                           REG_14_28_port, B2 => n170, ZN => n990);
   U1039 : AOI22_X1 port map( A1 => REG_8_28_port, A2 => n224_port, B1 => 
                           REG_10_28_port, B2 => n206_port, ZN => n989);
   U1040 : NAND4_X1 port map( A1 => n992, A2 => n991, A3 => n990, A4 => n989, 
                           ZN => n993);
   U1041 : AOI22_X1 port map( A1 => n994, A2 => n85, B1 => n993, B2 => n83, ZN 
                           => n995);
   U1042 : OAI221_X1 port map( B1 => n1061, B2 => n997, C1 => n1059, C2 => n996
                           , A => n995, ZN => N255);
   U1043 : AOI22_X1 port map( A1 => REG_21_29_port, A2 => n116, B1 => 
                           REG_23_29_port, B2 => n98, ZN => n1001);
   U1044 : AOI22_X1 port map( A1 => REG_17_29_port, A2 => n152, B1 => 
                           REG_19_29_port, B2 => n134, ZN => n1000);
   U1045 : AOI22_X1 port map( A1 => REG_20_29_port, A2 => n188_port, B1 => 
                           REG_22_29_port, B2 => n170, ZN => n999);
   U1046 : AOI22_X1 port map( A1 => REG_16_29_port, A2 => n224_port, B1 => 
                           REG_18_29_port, B2 => n206_port, ZN => n998);
   U1047 : AND4_X1 port map( A1 => n1001, A2 => n1000, A3 => n999, A4 => n998, 
                           ZN => n1018);
   U1048 : AOI22_X1 port map( A1 => REG_29_29_port, A2 => n116, B1 => 
                           REG_31_29_port, B2 => n98, ZN => n1005);
   U1049 : AOI22_X1 port map( A1 => REG_25_29_port, A2 => n152, B1 => 
                           REG_27_29_port, B2 => n134, ZN => n1004);
   U1050 : AOI22_X1 port map( A1 => REG_28_29_port, A2 => n188_port, B1 => 
                           REG_30_29_port, B2 => n170, ZN => n1003);
   U1051 : AOI22_X1 port map( A1 => REG_24_29_port, A2 => n224_port, B1 => 
                           REG_26_29_port, B2 => n206_port, ZN => n1002);
   U1052 : AND4_X1 port map( A1 => n1005, A2 => n1004, A3 => n1003, A4 => n1002
                           , ZN => n1017);
   U1053 : AOI22_X1 port map( A1 => REG_5_29_port, A2 => n116, B1 => 
                           REG_7_29_port, B2 => n98, ZN => n1009);
   U1054 : AOI22_X1 port map( A1 => REG_1_29_port, A2 => n152, B1 => 
                           REG_3_29_port, B2 => n134, ZN => n1008);
   U1055 : AOI22_X1 port map( A1 => REG_4_29_port, A2 => n188_port, B1 => 
                           REG_6_29_port, B2 => n170, ZN => n1007);
   U1056 : AOI22_X1 port map( A1 => REG_0_29_port, A2 => n224_port, B1 => 
                           REG_2_29_port, B2 => n206_port, ZN => n1006);
   U1057 : NAND4_X1 port map( A1 => n1009, A2 => n1008, A3 => n1007, A4 => 
                           n1006, ZN => n1015);
   U1058 : AOI22_X1 port map( A1 => REG_13_29_port, A2 => n116, B1 => 
                           REG_15_29_port, B2 => n98, ZN => n1013);
   U1059 : AOI22_X1 port map( A1 => REG_9_29_port, A2 => n152, B1 => 
                           REG_11_29_port, B2 => n134, ZN => n1012);
   U1060 : AOI22_X1 port map( A1 => REG_12_29_port, A2 => n188_port, B1 => 
                           REG_14_29_port, B2 => n170, ZN => n1011);
   U1061 : AOI22_X1 port map( A1 => REG_8_29_port, A2 => n224_port, B1 => 
                           REG_10_29_port, B2 => n206_port, ZN => n1010);
   U1062 : NAND4_X1 port map( A1 => n1013, A2 => n1012, A3 => n1011, A4 => 
                           n1010, ZN => n1014);
   U1063 : AOI22_X1 port map( A1 => n1015, A2 => n85, B1 => n1014, B2 => n83, 
                           ZN => n1016);
   U1064 : OAI221_X1 port map( B1 => n1061, B2 => n1018, C1 => n1059, C2 => 
                           n1017, A => n1016, ZN => N254);
   U1065 : AOI22_X1 port map( A1 => REG_21_30_port, A2 => n116, B1 => 
                           REG_23_30_port, B2 => n98, ZN => n1022);
   U1066 : AOI22_X1 port map( A1 => REG_17_30_port, A2 => n152, B1 => 
                           REG_19_30_port, B2 => n134, ZN => n1021);
   U1067 : AOI22_X1 port map( A1 => REG_20_30_port, A2 => n188_port, B1 => 
                           REG_22_30_port, B2 => n170, ZN => n1020);
   U1068 : AOI22_X1 port map( A1 => REG_16_30_port, A2 => n224_port, B1 => 
                           REG_18_30_port, B2 => n206_port, ZN => n1019);
   U1069 : AND4_X1 port map( A1 => n1022, A2 => n1021, A3 => n1020, A4 => n1019
                           , ZN => n1039);
   U1070 : AOI22_X1 port map( A1 => REG_29_30_port, A2 => n117, B1 => 
                           REG_31_30_port, B2 => n99, ZN => n1026);
   U1071 : AOI22_X1 port map( A1 => REG_25_30_port, A2 => n153, B1 => 
                           REG_27_30_port, B2 => n135, ZN => n1025);
   U1072 : AOI22_X1 port map( A1 => REG_28_30_port, A2 => n189_port, B1 => 
                           REG_30_30_port, B2 => n171, ZN => n1024);
   U1073 : AOI22_X1 port map( A1 => REG_24_30_port, A2 => n225_port, B1 => 
                           REG_26_30_port, B2 => n207_port, ZN => n1023);
   U1074 : AND4_X1 port map( A1 => n1026, A2 => n1025, A3 => n1024, A4 => n1023
                           , ZN => n1038);
   U1075 : AOI22_X1 port map( A1 => REG_5_30_port, A2 => n117, B1 => 
                           REG_7_30_port, B2 => n99, ZN => n1030);
   U1076 : AOI22_X1 port map( A1 => REG_1_30_port, A2 => n153, B1 => 
                           REG_3_30_port, B2 => n135, ZN => n1029);
   U1077 : AOI22_X1 port map( A1 => REG_4_30_port, A2 => n189_port, B1 => 
                           REG_6_30_port, B2 => n171, ZN => n1028);
   U1078 : AOI22_X1 port map( A1 => REG_0_30_port, A2 => n225_port, B1 => 
                           REG_2_30_port, B2 => n207_port, ZN => n1027);
   U1079 : NAND4_X1 port map( A1 => n1030, A2 => n1029, A3 => n1028, A4 => 
                           n1027, ZN => n1036);
   U1080 : AOI22_X1 port map( A1 => REG_13_30_port, A2 => n117, B1 => 
                           REG_15_30_port, B2 => n99, ZN => n1034);
   U1081 : AOI22_X1 port map( A1 => REG_9_30_port, A2 => n153, B1 => 
                           REG_11_30_port, B2 => n135, ZN => n1033);
   U1082 : AOI22_X1 port map( A1 => REG_12_30_port, A2 => n189_port, B1 => 
                           REG_14_30_port, B2 => n171, ZN => n1032);
   U1083 : AOI22_X1 port map( A1 => REG_8_30_port, A2 => n225_port, B1 => 
                           REG_10_30_port, B2 => n207_port, ZN => n1031);
   U1084 : NAND4_X1 port map( A1 => n1034, A2 => n1033, A3 => n1032, A4 => 
                           n1031, ZN => n1035);
   U1085 : AOI22_X1 port map( A1 => n1036, A2 => n85, B1 => n1035, B2 => n83, 
                           ZN => n1037);
   U1086 : OAI221_X1 port map( B1 => n1061, B2 => n1039, C1 => n1059, C2 => 
                           n1038, A => n1037, ZN => N253);
   U1087 : AOI22_X1 port map( A1 => REG_21_31_port, A2 => n117, B1 => 
                           REG_23_31_port, B2 => n99, ZN => n1043);
   U1088 : AOI22_X1 port map( A1 => REG_17_31_port, A2 => n153, B1 => 
                           REG_19_31_port, B2 => n135, ZN => n1042);
   U1089 : AOI22_X1 port map( A1 => REG_20_31_port, A2 => n189_port, B1 => 
                           REG_22_31_port, B2 => n171, ZN => n1041);
   U1090 : AOI22_X1 port map( A1 => REG_16_31_port, A2 => n225_port, B1 => 
                           REG_18_31_port, B2 => n207_port, ZN => n1040);
   U1091 : AND4_X1 port map( A1 => n1043, A2 => n1042, A3 => n1041, A4 => n1040
                           , ZN => n1062);
   U1092 : AOI22_X1 port map( A1 => REG_29_31_port, A2 => n117, B1 => 
                           REG_31_31_port, B2 => n99, ZN => n1047);
   U1093 : AOI22_X1 port map( A1 => REG_25_31_port, A2 => n153, B1 => 
                           REG_27_31_port, B2 => n135, ZN => n1046);
   U1094 : AOI22_X1 port map( A1 => REG_28_31_port, A2 => n189_port, B1 => 
                           REG_30_31_port, B2 => n171, ZN => n1045);
   U1095 : AOI22_X1 port map( A1 => REG_24_31_port, A2 => n225_port, B1 => 
                           REG_26_31_port, B2 => n207_port, ZN => n1044);
   U1096 : AND4_X1 port map( A1 => n1047, A2 => n1046, A3 => n1045, A4 => n1044
                           , ZN => n1060);
   U1097 : AOI22_X1 port map( A1 => REG_5_31_port, A2 => n117, B1 => 
                           REG_7_31_port, B2 => n99, ZN => n1051);
   U1098 : AOI22_X1 port map( A1 => REG_1_31_port, A2 => n153, B1 => 
                           REG_3_31_port, B2 => n135, ZN => n1050);
   U1099 : AOI22_X1 port map( A1 => REG_4_31_port, A2 => n189_port, B1 => 
                           REG_6_31_port, B2 => n171, ZN => n1049);
   U1100 : AOI22_X1 port map( A1 => REG_0_31_port, A2 => n225_port, B1 => 
                           REG_2_31_port, B2 => n207_port, ZN => n1048);
   U1101 : NAND4_X1 port map( A1 => n1051, A2 => n1050, A3 => n1049, A4 => 
                           n1048, ZN => n1057);
   U1102 : AOI22_X1 port map( A1 => REG_13_31_port, A2 => n117, B1 => 
                           REG_15_31_port, B2 => n99, ZN => n1055);
   U1103 : AOI22_X1 port map( A1 => REG_9_31_port, A2 => n153, B1 => 
                           REG_11_31_port, B2 => n135, ZN => n1054);
   U1104 : AOI22_X1 port map( A1 => REG_12_31_port, A2 => n189_port, B1 => 
                           REG_14_31_port, B2 => n171, ZN => n1053);
   U1105 : AOI22_X1 port map( A1 => REG_8_31_port, A2 => n225_port, B1 => 
                           REG_10_31_port, B2 => n207_port, ZN => n1052);
   U1106 : NAND4_X1 port map( A1 => n1055, A2 => n1054, A3 => n1053, A4 => 
                           n1052, ZN => n1056);
   U1107 : AOI22_X1 port map( A1 => n85, A2 => n1057, B1 => n83, B2 => n1056, 
                           ZN => n1058);
   U1108 : OAI221_X1 port map( B1 => n1062, B2 => n1061, C1 => n1060, C2 => 
                           n1059, A => n1058, ZN => N252);
   U1109 : NOR2_X1 port map( A1 => n1746, A2 => ADD_RD2(1), ZN => n1067);
   U1110 : NOR2_X1 port map( A1 => n1746, A2 => n1747, ZN => n1068);
   U1111 : AOI22_X1 port map( A1 => REG_21_0_port, A2 => n250_port, B1 => 
                           REG_23_0_port, B2 => n232_port, ZN => n1074);
   U1112 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1069);
   U1113 : NOR2_X1 port map( A1 => n1747, A2 => ADD_RD2(2), ZN => n1070);
   U1114 : AOI22_X1 port map( A1 => REG_17_0_port, A2 => n286_port, B1 => 
                           REG_19_0_port, B2 => n268_port, ZN => n1073);
   U1115 : AOI22_X1 port map( A1 => REG_20_0_port, A2 => n322, B1 => 
                           REG_22_0_port, B2 => n304_port, ZN => n1072);
   U1116 : AOI22_X1 port map( A1 => REG_16_0_port, A2 => n358, B1 => 
                           REG_18_0_port, B2 => n340, ZN => n1071);
   U1117 : AND4_X1 port map( A1 => n1074, A2 => n1073, A3 => n1072, A4 => n1071
                           , ZN => n1091);
   U1118 : AOI22_X1 port map( A1 => REG_29_0_port, A2 => n250_port, B1 => 
                           REG_31_0_port, B2 => n232_port, ZN => n1078);
   U1119 : AOI22_X1 port map( A1 => REG_25_0_port, A2 => n286_port, B1 => 
                           REG_27_0_port, B2 => n268_port, ZN => n1077);
   U1120 : AOI22_X1 port map( A1 => REG_28_0_port, A2 => n322, B1 => 
                           REG_30_0_port, B2 => n304_port, ZN => n1076);
   U1121 : AOI22_X1 port map( A1 => REG_24_0_port, A2 => n358, B1 => 
                           REG_26_0_port, B2 => n340, ZN => n1075);
   U1122 : AND4_X1 port map( A1 => n1078, A2 => n1077, A3 => n1076, A4 => n1075
                           , ZN => n1090);
   U1123 : AOI22_X1 port map( A1 => REG_5_0_port, A2 => n250_port, B1 => 
                           REG_7_0_port, B2 => n232_port, ZN => n1082);
   U1124 : AOI22_X1 port map( A1 => REG_1_0_port, A2 => n286_port, B1 => 
                           REG_3_0_port, B2 => n268_port, ZN => n1081);
   U1125 : AOI22_X1 port map( A1 => REG_4_0_port, A2 => n322, B1 => 
                           REG_6_0_port, B2 => n304_port, ZN => n1080);
   U1126 : AOI22_X1 port map( A1 => REG_0_0_port, A2 => n358, B1 => 
                           REG_2_0_port, B2 => n340, ZN => n1079);
   U1127 : NAND4_X1 port map( A1 => n1082, A2 => n1081, A3 => n1080, A4 => 
                           n1079, ZN => n1088);
   U1128 : AOI22_X1 port map( A1 => REG_13_0_port, A2 => n250_port, B1 => 
                           REG_15_0_port, B2 => n232_port, ZN => n1086);
   U1129 : AOI22_X1 port map( A1 => REG_9_0_port, A2 => n286_port, B1 => 
                           REG_11_0_port, B2 => n268_port, ZN => n1085);
   U1130 : AOI22_X1 port map( A1 => REG_12_0_port, A2 => n322, B1 => 
                           REG_14_0_port, B2 => n304_port, ZN => n1084);
   U1131 : AOI22_X1 port map( A1 => REG_8_0_port, A2 => n358, B1 => 
                           REG_10_0_port, B2 => n340, ZN => n1083);
   U1132 : NAND4_X1 port map( A1 => n1086, A2 => n1085, A3 => n1084, A4 => 
                           n1083, ZN => n1087);
   U1133 : AOI22_X1 port map( A1 => n1088, A2 => n86, B1 => n1087, B2 => n84, 
                           ZN => n1089);
   U1134 : OAI221_X1 port map( B1 => n1743, B2 => n1091, C1 => n1741, C2 => 
                           n1090, A => n1089, ZN => N315);
   U1135 : AOI22_X1 port map( A1 => REG_21_1_port, A2 => n250_port, B1 => 
                           REG_23_1_port, B2 => n232_port, ZN => n1095);
   U1136 : AOI22_X1 port map( A1 => REG_17_1_port, A2 => n286_port, B1 => 
                           REG_19_1_port, B2 => n268_port, ZN => n1094);
   U1137 : AOI22_X1 port map( A1 => REG_20_1_port, A2 => n322, B1 => 
                           REG_22_1_port, B2 => n304_port, ZN => n1093);
   U1138 : AOI22_X1 port map( A1 => REG_16_1_port, A2 => n358, B1 => 
                           REG_18_1_port, B2 => n340, ZN => n1092);
   U1139 : AND4_X1 port map( A1 => n1095, A2 => n1094, A3 => n1093, A4 => n1092
                           , ZN => n1112);
   U1140 : AOI22_X1 port map( A1 => REG_29_1_port, A2 => n250_port, B1 => 
                           REG_31_1_port, B2 => n232_port, ZN => n1099);
   U1141 : AOI22_X1 port map( A1 => REG_25_1_port, A2 => n286_port, B1 => 
                           REG_27_1_port, B2 => n268_port, ZN => n1098);
   U1142 : AOI22_X1 port map( A1 => REG_28_1_port, A2 => n322, B1 => 
                           REG_30_1_port, B2 => n304_port, ZN => n1097);
   U1143 : AOI22_X1 port map( A1 => REG_24_1_port, A2 => n358, B1 => 
                           REG_26_1_port, B2 => n340, ZN => n1096);
   U1144 : AND4_X1 port map( A1 => n1099, A2 => n1098, A3 => n1097, A4 => n1096
                           , ZN => n1111);
   U1145 : AOI22_X1 port map( A1 => REG_5_1_port, A2 => n250_port, B1 => 
                           REG_7_1_port, B2 => n232_port, ZN => n1103);
   U1146 : AOI22_X1 port map( A1 => REG_1_1_port, A2 => n286_port, B1 => 
                           REG_3_1_port, B2 => n268_port, ZN => n1102);
   U1147 : AOI22_X1 port map( A1 => REG_4_1_port, A2 => n322, B1 => 
                           REG_6_1_port, B2 => n304_port, ZN => n1101);
   U1148 : AOI22_X1 port map( A1 => REG_0_1_port, A2 => n358, B1 => 
                           REG_2_1_port, B2 => n340, ZN => n1100);
   U1149 : NAND4_X1 port map( A1 => n1103, A2 => n1102, A3 => n1101, A4 => 
                           n1100, ZN => n1109);
   U1150 : AOI22_X1 port map( A1 => REG_13_1_port, A2 => n250_port, B1 => 
                           REG_15_1_port, B2 => n232_port, ZN => n1107);
   U1151 : AOI22_X1 port map( A1 => REG_9_1_port, A2 => n286_port, B1 => 
                           REG_11_1_port, B2 => n268_port, ZN => n1106);
   U1152 : AOI22_X1 port map( A1 => REG_12_1_port, A2 => n322, B1 => 
                           REG_14_1_port, B2 => n304_port, ZN => n1105);
   U1153 : AOI22_X1 port map( A1 => REG_8_1_port, A2 => n358, B1 => 
                           REG_10_1_port, B2 => n340, ZN => n1104);
   U1154 : NAND4_X1 port map( A1 => n1107, A2 => n1106, A3 => n1105, A4 => 
                           n1104, ZN => n1108);
   U1155 : AOI22_X1 port map( A1 => n1109, A2 => n86, B1 => n1108, B2 => n84, 
                           ZN => n1110);
   U1156 : OAI221_X1 port map( B1 => n1743, B2 => n1112, C1 => n1741, C2 => 
                           n1111, A => n1110, ZN => N314);
   U1157 : AOI22_X1 port map( A1 => REG_21_2_port, A2 => n250_port, B1 => 
                           REG_23_2_port, B2 => n232_port, ZN => n1116);
   U1158 : AOI22_X1 port map( A1 => REG_17_2_port, A2 => n286_port, B1 => 
                           REG_19_2_port, B2 => n268_port, ZN => n1115);
   U1159 : AOI22_X1 port map( A1 => REG_20_2_port, A2 => n322, B1 => 
                           REG_22_2_port, B2 => n304_port, ZN => n1114);
   U1160 : AOI22_X1 port map( A1 => REG_16_2_port, A2 => n358, B1 => 
                           REG_18_2_port, B2 => n340, ZN => n1113);
   U1161 : AND4_X1 port map( A1 => n1116, A2 => n1115, A3 => n1114, A4 => n1113
                           , ZN => n1133);
   U1162 : AOI22_X1 port map( A1 => REG_29_2_port, A2 => n250_port, B1 => 
                           REG_31_2_port, B2 => n232_port, ZN => n1120);
   U1163 : AOI22_X1 port map( A1 => REG_25_2_port, A2 => n286_port, B1 => 
                           REG_27_2_port, B2 => n268_port, ZN => n1119);
   U1164 : AOI22_X1 port map( A1 => REG_28_2_port, A2 => n322, B1 => 
                           REG_30_2_port, B2 => n304_port, ZN => n1118);
   U1165 : AOI22_X1 port map( A1 => REG_24_2_port, A2 => n358, B1 => 
                           REG_26_2_port, B2 => n340, ZN => n1117);
   U1166 : AND4_X1 port map( A1 => n1120, A2 => n1119, A3 => n1118, A4 => n1117
                           , ZN => n1132);
   U1167 : AOI22_X1 port map( A1 => REG_5_2_port, A2 => n250_port, B1 => 
                           REG_7_2_port, B2 => n232_port, ZN => n1124);
   U1168 : AOI22_X1 port map( A1 => REG_1_2_port, A2 => n286_port, B1 => 
                           REG_3_2_port, B2 => n268_port, ZN => n1123);
   U1169 : AOI22_X1 port map( A1 => REG_4_2_port, A2 => n322, B1 => 
                           REG_6_2_port, B2 => n304_port, ZN => n1122);
   U1170 : AOI22_X1 port map( A1 => REG_0_2_port, A2 => n358, B1 => 
                           REG_2_2_port, B2 => n340, ZN => n1121);
   U1171 : NAND4_X1 port map( A1 => n1124, A2 => n1123, A3 => n1122, A4 => 
                           n1121, ZN => n1130);
   U1172 : AOI22_X1 port map( A1 => REG_13_2_port, A2 => n251, B1 => 
                           REG_15_2_port, B2 => n233_port, ZN => n1128);
   U1173 : AOI22_X1 port map( A1 => REG_9_2_port, A2 => n287_port, B1 => 
                           REG_11_2_port, B2 => n269_port, ZN => n1127);
   U1174 : AOI22_X1 port map( A1 => REG_12_2_port, A2 => n323, B1 => 
                           REG_14_2_port, B2 => n305_port, ZN => n1126);
   U1175 : AOI22_X1 port map( A1 => REG_8_2_port, A2 => n359, B1 => 
                           REG_10_2_port, B2 => n341, ZN => n1125);
   U1176 : NAND4_X1 port map( A1 => n1128, A2 => n1127, A3 => n1126, A4 => 
                           n1125, ZN => n1129);
   U1177 : AOI22_X1 port map( A1 => n1130, A2 => n86, B1 => n1129, B2 => n84, 
                           ZN => n1131);
   U1178 : OAI221_X1 port map( B1 => n1743, B2 => n1133, C1 => n1741, C2 => 
                           n1132, A => n1131, ZN => N313);
   U1179 : AOI22_X1 port map( A1 => REG_21_3_port, A2 => n251, B1 => 
                           REG_23_3_port, B2 => n233_port, ZN => n1137);
   U1180 : AOI22_X1 port map( A1 => REG_17_3_port, A2 => n287_port, B1 => 
                           REG_19_3_port, B2 => n269_port, ZN => n1136);
   U1181 : AOI22_X1 port map( A1 => REG_20_3_port, A2 => n323, B1 => 
                           REG_22_3_port, B2 => n305_port, ZN => n1135);
   U1182 : AOI22_X1 port map( A1 => REG_16_3_port, A2 => n359, B1 => 
                           REG_18_3_port, B2 => n341, ZN => n1134);
   U1183 : AND4_X1 port map( A1 => n1137, A2 => n1136, A3 => n1135, A4 => n1134
                           , ZN => n1154);
   U1184 : AOI22_X1 port map( A1 => REG_29_3_port, A2 => n251, B1 => 
                           REG_31_3_port, B2 => n233_port, ZN => n1141);
   U1185 : AOI22_X1 port map( A1 => REG_25_3_port, A2 => n287_port, B1 => 
                           REG_27_3_port, B2 => n269_port, ZN => n1140);
   U1186 : AOI22_X1 port map( A1 => REG_28_3_port, A2 => n323, B1 => 
                           REG_30_3_port, B2 => n305_port, ZN => n1139);
   U1187 : AOI22_X1 port map( A1 => REG_24_3_port, A2 => n359, B1 => 
                           REG_26_3_port, B2 => n341, ZN => n1138);
   U1188 : AND4_X1 port map( A1 => n1141, A2 => n1140, A3 => n1139, A4 => n1138
                           , ZN => n1153);
   U1189 : AOI22_X1 port map( A1 => REG_5_3_port, A2 => n251, B1 => 
                           REG_7_3_port, B2 => n233_port, ZN => n1145);
   U1190 : AOI22_X1 port map( A1 => REG_1_3_port, A2 => n287_port, B1 => 
                           REG_3_3_port, B2 => n269_port, ZN => n1144);
   U1191 : AOI22_X1 port map( A1 => REG_4_3_port, A2 => n323, B1 => 
                           REG_6_3_port, B2 => n305_port, ZN => n1143);
   U1192 : AOI22_X1 port map( A1 => REG_0_3_port, A2 => n359, B1 => 
                           REG_2_3_port, B2 => n341, ZN => n1142);
   U1193 : NAND4_X1 port map( A1 => n1145, A2 => n1144, A3 => n1143, A4 => 
                           n1142, ZN => n1151);
   U1194 : AOI22_X1 port map( A1 => REG_13_3_port, A2 => n251, B1 => 
                           REG_15_3_port, B2 => n233_port, ZN => n1149);
   U1195 : AOI22_X1 port map( A1 => REG_9_3_port, A2 => n287_port, B1 => 
                           REG_11_3_port, B2 => n269_port, ZN => n1148);
   U1196 : AOI22_X1 port map( A1 => REG_12_3_port, A2 => n323, B1 => 
                           REG_14_3_port, B2 => n305_port, ZN => n1147);
   U1197 : AOI22_X1 port map( A1 => REG_8_3_port, A2 => n359, B1 => 
                           REG_10_3_port, B2 => n341, ZN => n1146);
   U1198 : NAND4_X1 port map( A1 => n1149, A2 => n1148, A3 => n1147, A4 => 
                           n1146, ZN => n1150);
   U1199 : AOI22_X1 port map( A1 => n1151, A2 => n86, B1 => n1150, B2 => n84, 
                           ZN => n1152);
   U1200 : OAI221_X1 port map( B1 => n1743, B2 => n1154, C1 => n1741, C2 => 
                           n1153, A => n1152, ZN => N312);
   U1201 : AOI22_X1 port map( A1 => REG_21_4_port, A2 => n251, B1 => 
                           REG_23_4_port, B2 => n233_port, ZN => n1158);
   U1202 : AOI22_X1 port map( A1 => REG_17_4_port, A2 => n287_port, B1 => 
                           REG_19_4_port, B2 => n269_port, ZN => n1157);
   U1203 : AOI22_X1 port map( A1 => REG_20_4_port, A2 => n323, B1 => 
                           REG_22_4_port, B2 => n305_port, ZN => n1156);
   U1204 : AOI22_X1 port map( A1 => REG_16_4_port, A2 => n359, B1 => 
                           REG_18_4_port, B2 => n341, ZN => n1155);
   U1205 : AND4_X1 port map( A1 => n1158, A2 => n1157, A3 => n1156, A4 => n1155
                           , ZN => n1175);
   U1206 : AOI22_X1 port map( A1 => REG_29_4_port, A2 => n251, B1 => 
                           REG_31_4_port, B2 => n233_port, ZN => n1162);
   U1207 : AOI22_X1 port map( A1 => REG_25_4_port, A2 => n287_port, B1 => 
                           REG_27_4_port, B2 => n269_port, ZN => n1161);
   U1208 : AOI22_X1 port map( A1 => REG_28_4_port, A2 => n323, B1 => 
                           REG_30_4_port, B2 => n305_port, ZN => n1160);
   U1209 : AOI22_X1 port map( A1 => REG_24_4_port, A2 => n359, B1 => 
                           REG_26_4_port, B2 => n341, ZN => n1159);
   U1210 : AND4_X1 port map( A1 => n1162, A2 => n1161, A3 => n1160, A4 => n1159
                           , ZN => n1174);
   U1211 : AOI22_X1 port map( A1 => REG_5_4_port, A2 => n251, B1 => 
                           REG_7_4_port, B2 => n233_port, ZN => n1166);
   U1212 : AOI22_X1 port map( A1 => REG_1_4_port, A2 => n287_port, B1 => 
                           REG_3_4_port, B2 => n269_port, ZN => n1165);
   U1213 : AOI22_X1 port map( A1 => REG_4_4_port, A2 => n323, B1 => 
                           REG_6_4_port, B2 => n305_port, ZN => n1164);
   U1214 : AOI22_X1 port map( A1 => REG_0_4_port, A2 => n359, B1 => 
                           REG_2_4_port, B2 => n341, ZN => n1163);
   U1215 : NAND4_X1 port map( A1 => n1166, A2 => n1165, A3 => n1164, A4 => 
                           n1163, ZN => n1172);
   U1216 : AOI22_X1 port map( A1 => REG_13_4_port, A2 => n251, B1 => 
                           REG_15_4_port, B2 => n233_port, ZN => n1170);
   U1217 : AOI22_X1 port map( A1 => REG_9_4_port, A2 => n287_port, B1 => 
                           REG_11_4_port, B2 => n269_port, ZN => n1169);
   U1218 : AOI22_X1 port map( A1 => REG_12_4_port, A2 => n323, B1 => 
                           REG_14_4_port, B2 => n305_port, ZN => n1168);
   U1219 : AOI22_X1 port map( A1 => REG_8_4_port, A2 => n359, B1 => 
                           REG_10_4_port, B2 => n341, ZN => n1167);
   U1220 : NAND4_X1 port map( A1 => n1170, A2 => n1169, A3 => n1168, A4 => 
                           n1167, ZN => n1171);
   U1221 : AOI22_X1 port map( A1 => n1172, A2 => n86, B1 => n1171, B2 => n84, 
                           ZN => n1173);
   U1222 : OAI221_X1 port map( B1 => n1743, B2 => n1175, C1 => n1741, C2 => 
                           n1174, A => n1173, ZN => N311);
   U1223 : AOI22_X1 port map( A1 => REG_21_5_port, A2 => n251, B1 => 
                           REG_23_5_port, B2 => n233_port, ZN => n1179);
   U1224 : AOI22_X1 port map( A1 => REG_17_5_port, A2 => n287_port, B1 => 
                           REG_19_5_port, B2 => n269_port, ZN => n1178);
   U1225 : AOI22_X1 port map( A1 => REG_20_5_port, A2 => n323, B1 => 
                           REG_22_5_port, B2 => n305_port, ZN => n1177);
   U1226 : AOI22_X1 port map( A1 => REG_16_5_port, A2 => n359, B1 => 
                           REG_18_5_port, B2 => n341, ZN => n1176);
   U1227 : AND4_X1 port map( A1 => n1179, A2 => n1178, A3 => n1177, A4 => n1176
                           , ZN => n1196);
   U1228 : AOI22_X1 port map( A1 => REG_29_5_port, A2 => n251, B1 => 
                           REG_31_5_port, B2 => n233_port, ZN => n1183);
   U1229 : AOI22_X1 port map( A1 => REG_25_5_port, A2 => n287_port, B1 => 
                           REG_27_5_port, B2 => n269_port, ZN => n1182);
   U1230 : AOI22_X1 port map( A1 => REG_28_5_port, A2 => n323, B1 => 
                           REG_30_5_port, B2 => n305_port, ZN => n1181);
   U1231 : AOI22_X1 port map( A1 => REG_24_5_port, A2 => n359, B1 => 
                           REG_26_5_port, B2 => n341, ZN => n1180);
   U1232 : AND4_X1 port map( A1 => n1183, A2 => n1182, A3 => n1181, A4 => n1180
                           , ZN => n1195);
   U1233 : AOI22_X1 port map( A1 => REG_5_5_port, A2 => n252_port, B1 => 
                           REG_7_5_port, B2 => n234_port, ZN => n1187);
   U1234 : AOI22_X1 port map( A1 => REG_1_5_port, A2 => n288_port, B1 => 
                           REG_3_5_port, B2 => n270_port, ZN => n1186);
   U1235 : AOI22_X1 port map( A1 => REG_4_5_port, A2 => n324, B1 => 
                           REG_6_5_port, B2 => n306_port, ZN => n1185);
   U1236 : AOI22_X1 port map( A1 => REG_0_5_port, A2 => n360, B1 => 
                           REG_2_5_port, B2 => n342, ZN => n1184);
   U1237 : NAND4_X1 port map( A1 => n1187, A2 => n1186, A3 => n1185, A4 => 
                           n1184, ZN => n1193);
   U1238 : AOI22_X1 port map( A1 => REG_13_5_port, A2 => n252_port, B1 => 
                           REG_15_5_port, B2 => n234_port, ZN => n1191);
   U1239 : AOI22_X1 port map( A1 => REG_9_5_port, A2 => n288_port, B1 => 
                           REG_11_5_port, B2 => n270_port, ZN => n1190);
   U1240 : AOI22_X1 port map( A1 => REG_12_5_port, A2 => n324, B1 => 
                           REG_14_5_port, B2 => n306_port, ZN => n1189);
   U1241 : AOI22_X1 port map( A1 => REG_8_5_port, A2 => n360, B1 => 
                           REG_10_5_port, B2 => n342, ZN => n1188);
   U1242 : NAND4_X1 port map( A1 => n1191, A2 => n1190, A3 => n1189, A4 => 
                           n1188, ZN => n1192);
   U1243 : AOI22_X1 port map( A1 => n1193, A2 => n86, B1 => n1192, B2 => n84, 
                           ZN => n1194);
   U1244 : OAI221_X1 port map( B1 => n1743, B2 => n1196, C1 => n1741, C2 => 
                           n1195, A => n1194, ZN => N310);
   U1245 : AOI22_X1 port map( A1 => REG_21_6_port, A2 => n252_port, B1 => 
                           REG_23_6_port, B2 => n234_port, ZN => n1200);
   U1246 : AOI22_X1 port map( A1 => REG_17_6_port, A2 => n288_port, B1 => 
                           REG_19_6_port, B2 => n270_port, ZN => n1199);
   U1247 : AOI22_X1 port map( A1 => REG_20_6_port, A2 => n324, B1 => 
                           REG_22_6_port, B2 => n306_port, ZN => n1198);
   U1248 : AOI22_X1 port map( A1 => REG_16_6_port, A2 => n360, B1 => 
                           REG_18_6_port, B2 => n342, ZN => n1197);
   U1249 : AND4_X1 port map( A1 => n1200, A2 => n1199, A3 => n1198, A4 => n1197
                           , ZN => n1217);
   U1250 : AOI22_X1 port map( A1 => REG_29_6_port, A2 => n252_port, B1 => 
                           REG_31_6_port, B2 => n234_port, ZN => n1204);
   U1251 : AOI22_X1 port map( A1 => REG_25_6_port, A2 => n288_port, B1 => 
                           REG_27_6_port, B2 => n270_port, ZN => n1203);
   U1252 : AOI22_X1 port map( A1 => REG_28_6_port, A2 => n324, B1 => 
                           REG_30_6_port, B2 => n306_port, ZN => n1202);
   U1253 : AOI22_X1 port map( A1 => REG_24_6_port, A2 => n360, B1 => 
                           REG_26_6_port, B2 => n342, ZN => n1201);
   U1254 : AND4_X1 port map( A1 => n1204, A2 => n1203, A3 => n1202, A4 => n1201
                           , ZN => n1216);
   U1255 : AOI22_X1 port map( A1 => REG_5_6_port, A2 => n252_port, B1 => 
                           REG_7_6_port, B2 => n234_port, ZN => n1208);
   U1256 : AOI22_X1 port map( A1 => REG_1_6_port, A2 => n288_port, B1 => 
                           REG_3_6_port, B2 => n270_port, ZN => n1207);
   U1257 : AOI22_X1 port map( A1 => REG_4_6_port, A2 => n324, B1 => 
                           REG_6_6_port, B2 => n306_port, ZN => n1206);
   U1258 : AOI22_X1 port map( A1 => REG_0_6_port, A2 => n360, B1 => 
                           REG_2_6_port, B2 => n342, ZN => n1205);
   U1259 : NAND4_X1 port map( A1 => n1208, A2 => n1207, A3 => n1206, A4 => 
                           n1205, ZN => n1214);
   U1260 : AOI22_X1 port map( A1 => REG_13_6_port, A2 => n252_port, B1 => 
                           REG_15_6_port, B2 => n234_port, ZN => n1212);
   U1261 : AOI22_X1 port map( A1 => REG_9_6_port, A2 => n288_port, B1 => 
                           REG_11_6_port, B2 => n270_port, ZN => n1211);
   U1262 : AOI22_X1 port map( A1 => REG_12_6_port, A2 => n324, B1 => 
                           REG_14_6_port, B2 => n306_port, ZN => n1210);
   U1263 : AOI22_X1 port map( A1 => REG_8_6_port, A2 => n360, B1 => 
                           REG_10_6_port, B2 => n342, ZN => n1209);
   U1264 : NAND4_X1 port map( A1 => n1212, A2 => n1211, A3 => n1210, A4 => 
                           n1209, ZN => n1213);
   U1265 : AOI22_X1 port map( A1 => n1214, A2 => n86, B1 => n1213, B2 => n84, 
                           ZN => n1215);
   U1266 : OAI221_X1 port map( B1 => n1743, B2 => n1217, C1 => n1741, C2 => 
                           n1216, A => n1215, ZN => N309);
   U1267 : AOI22_X1 port map( A1 => REG_21_7_port, A2 => n252_port, B1 => 
                           REG_23_7_port, B2 => n234_port, ZN => n1221);
   U1268 : AOI22_X1 port map( A1 => REG_17_7_port, A2 => n288_port, B1 => 
                           REG_19_7_port, B2 => n270_port, ZN => n1220);
   U1269 : AOI22_X1 port map( A1 => REG_20_7_port, A2 => n324, B1 => 
                           REG_22_7_port, B2 => n306_port, ZN => n1219);
   U1270 : AOI22_X1 port map( A1 => REG_16_7_port, A2 => n360, B1 => 
                           REG_18_7_port, B2 => n342, ZN => n1218);
   U1271 : AND4_X1 port map( A1 => n1221, A2 => n1220, A3 => n1219, A4 => n1218
                           , ZN => n1238);
   U1272 : AOI22_X1 port map( A1 => REG_29_7_port, A2 => n252_port, B1 => 
                           REG_31_7_port, B2 => n234_port, ZN => n1225);
   U1273 : AOI22_X1 port map( A1 => REG_25_7_port, A2 => n288_port, B1 => 
                           REG_27_7_port, B2 => n270_port, ZN => n1224);
   U1274 : AOI22_X1 port map( A1 => REG_28_7_port, A2 => n324, B1 => 
                           REG_30_7_port, B2 => n306_port, ZN => n1223);
   U1275 : AOI22_X1 port map( A1 => REG_24_7_port, A2 => n360, B1 => 
                           REG_26_7_port, B2 => n342, ZN => n1222);
   U1276 : AND4_X1 port map( A1 => n1225, A2 => n1224, A3 => n1223, A4 => n1222
                           , ZN => n1237);
   U1277 : AOI22_X1 port map( A1 => REG_5_7_port, A2 => n252_port, B1 => 
                           REG_7_7_port, B2 => n234_port, ZN => n1229);
   U1278 : AOI22_X1 port map( A1 => REG_1_7_port, A2 => n288_port, B1 => 
                           REG_3_7_port, B2 => n270_port, ZN => n1228);
   U1279 : AOI22_X1 port map( A1 => REG_4_7_port, A2 => n324, B1 => 
                           REG_6_7_port, B2 => n306_port, ZN => n1227);
   U1280 : AOI22_X1 port map( A1 => REG_0_7_port, A2 => n360, B1 => 
                           REG_2_7_port, B2 => n342, ZN => n1226);
   U1281 : NAND4_X1 port map( A1 => n1229, A2 => n1228, A3 => n1227, A4 => 
                           n1226, ZN => n1235);
   U1282 : AOI22_X1 port map( A1 => REG_13_7_port, A2 => n252_port, B1 => 
                           REG_15_7_port, B2 => n234_port, ZN => n1233);
   U1283 : AOI22_X1 port map( A1 => REG_9_7_port, A2 => n288_port, B1 => 
                           REG_11_7_port, B2 => n270_port, ZN => n1232);
   U1284 : AOI22_X1 port map( A1 => REG_12_7_port, A2 => n324, B1 => 
                           REG_14_7_port, B2 => n306_port, ZN => n1231);
   U1285 : AOI22_X1 port map( A1 => REG_8_7_port, A2 => n360, B1 => 
                           REG_10_7_port, B2 => n342, ZN => n1230);
   U1286 : NAND4_X1 port map( A1 => n1233, A2 => n1232, A3 => n1231, A4 => 
                           n1230, ZN => n1234);
   U1287 : AOI22_X1 port map( A1 => n1235, A2 => n86, B1 => n1234, B2 => n84, 
                           ZN => n1236);
   U1288 : OAI221_X1 port map( B1 => n1743, B2 => n1238, C1 => n1741, C2 => 
                           n1237, A => n1236, ZN => N308);
   U1289 : AOI22_X1 port map( A1 => REG_21_8_port, A2 => n252_port, B1 => 
                           REG_23_8_port, B2 => n234_port, ZN => n1242);
   U1290 : AOI22_X1 port map( A1 => REG_17_8_port, A2 => n288_port, B1 => 
                           REG_19_8_port, B2 => n270_port, ZN => n1241);
   U1291 : AOI22_X1 port map( A1 => REG_20_8_port, A2 => n324, B1 => 
                           REG_22_8_port, B2 => n306_port, ZN => n1240);
   U1292 : AOI22_X1 port map( A1 => REG_16_8_port, A2 => n360, B1 => 
                           REG_18_8_port, B2 => n342, ZN => n1239);
   U1293 : AND4_X1 port map( A1 => n1242, A2 => n1241, A3 => n1240, A4 => n1239
                           , ZN => n1259);
   U1294 : AOI22_X1 port map( A1 => REG_29_8_port, A2 => n253_port, B1 => 
                           REG_31_8_port, B2 => n235_port, ZN => n1246);
   U1295 : AOI22_X1 port map( A1 => REG_25_8_port, A2 => n289_port, B1 => 
                           REG_27_8_port, B2 => n271_port, ZN => n1245);
   U1296 : AOI22_X1 port map( A1 => REG_28_8_port, A2 => n325, B1 => 
                           REG_30_8_port, B2 => n307_port, ZN => n1244);
   U1297 : AOI22_X1 port map( A1 => REG_24_8_port, A2 => n361, B1 => 
                           REG_26_8_port, B2 => n343, ZN => n1243);
   U1298 : AND4_X1 port map( A1 => n1246, A2 => n1245, A3 => n1244, A4 => n1243
                           , ZN => n1258);
   U1299 : AOI22_X1 port map( A1 => REG_5_8_port, A2 => n253_port, B1 => 
                           REG_7_8_port, B2 => n235_port, ZN => n1250);
   U1300 : AOI22_X1 port map( A1 => REG_1_8_port, A2 => n289_port, B1 => 
                           REG_3_8_port, B2 => n271_port, ZN => n1249);
   U1301 : AOI22_X1 port map( A1 => REG_4_8_port, A2 => n325, B1 => 
                           REG_6_8_port, B2 => n307_port, ZN => n1248);
   U1302 : AOI22_X1 port map( A1 => REG_0_8_port, A2 => n361, B1 => 
                           REG_2_8_port, B2 => n343, ZN => n1247);
   U1303 : NAND4_X1 port map( A1 => n1250, A2 => n1249, A3 => n1248, A4 => 
                           n1247, ZN => n1256);
   U1304 : AOI22_X1 port map( A1 => REG_13_8_port, A2 => n253_port, B1 => 
                           REG_15_8_port, B2 => n235_port, ZN => n1254);
   U1305 : AOI22_X1 port map( A1 => REG_9_8_port, A2 => n289_port, B1 => 
                           REG_11_8_port, B2 => n271_port, ZN => n1253);
   U1306 : AOI22_X1 port map( A1 => REG_12_8_port, A2 => n325, B1 => 
                           REG_14_8_port, B2 => n307_port, ZN => n1252);
   U1307 : AOI22_X1 port map( A1 => REG_8_8_port, A2 => n361, B1 => 
                           REG_10_8_port, B2 => n343, ZN => n1251);
   U1308 : NAND4_X1 port map( A1 => n1254, A2 => n1253, A3 => n1252, A4 => 
                           n1251, ZN => n1255);
   U1309 : AOI22_X1 port map( A1 => n1256, A2 => n86, B1 => n1255, B2 => n84, 
                           ZN => n1257);
   U1310 : OAI221_X1 port map( B1 => n1743, B2 => n1259, C1 => n1741, C2 => 
                           n1258, A => n1257, ZN => N307);
   U1311 : AOI22_X1 port map( A1 => REG_21_9_port, A2 => n253_port, B1 => 
                           REG_23_9_port, B2 => n235_port, ZN => n1263);
   U1312 : AOI22_X1 port map( A1 => REG_17_9_port, A2 => n289_port, B1 => 
                           REG_19_9_port, B2 => n271_port, ZN => n1262);
   U1313 : AOI22_X1 port map( A1 => REG_20_9_port, A2 => n325, B1 => 
                           REG_22_9_port, B2 => n307_port, ZN => n1261);
   U1314 : AOI22_X1 port map( A1 => REG_16_9_port, A2 => n361, B1 => 
                           REG_18_9_port, B2 => n343, ZN => n1260);
   U1315 : AND4_X1 port map( A1 => n1263, A2 => n1262, A3 => n1261, A4 => n1260
                           , ZN => n1280);
   U1316 : AOI22_X1 port map( A1 => REG_29_9_port, A2 => n253_port, B1 => 
                           REG_31_9_port, B2 => n235_port, ZN => n1267);
   U1317 : AOI22_X1 port map( A1 => REG_25_9_port, A2 => n289_port, B1 => 
                           REG_27_9_port, B2 => n271_port, ZN => n1266);
   U1318 : AOI22_X1 port map( A1 => REG_28_9_port, A2 => n325, B1 => 
                           REG_30_9_port, B2 => n307_port, ZN => n1265);
   U1319 : AOI22_X1 port map( A1 => REG_24_9_port, A2 => n361, B1 => 
                           REG_26_9_port, B2 => n343, ZN => n1264);
   U1320 : AND4_X1 port map( A1 => n1267, A2 => n1266, A3 => n1265, A4 => n1264
                           , ZN => n1279);
   U1321 : AOI22_X1 port map( A1 => REG_5_9_port, A2 => n253_port, B1 => 
                           REG_7_9_port, B2 => n235_port, ZN => n1271);
   U1322 : AOI22_X1 port map( A1 => REG_1_9_port, A2 => n289_port, B1 => 
                           REG_3_9_port, B2 => n271_port, ZN => n1270);
   U1323 : AOI22_X1 port map( A1 => REG_4_9_port, A2 => n325, B1 => 
                           REG_6_9_port, B2 => n307_port, ZN => n1269);
   U1324 : AOI22_X1 port map( A1 => REG_0_9_port, A2 => n361, B1 => 
                           REG_2_9_port, B2 => n343, ZN => n1268);
   U1325 : NAND4_X1 port map( A1 => n1271, A2 => n1270, A3 => n1269, A4 => 
                           n1268, ZN => n1277);
   U1326 : AOI22_X1 port map( A1 => REG_13_9_port, A2 => n253_port, B1 => 
                           REG_15_9_port, B2 => n235_port, ZN => n1275);
   U1327 : AOI22_X1 port map( A1 => REG_9_9_port, A2 => n289_port, B1 => 
                           REG_11_9_port, B2 => n271_port, ZN => n1274);
   U1328 : AOI22_X1 port map( A1 => REG_12_9_port, A2 => n325, B1 => 
                           REG_14_9_port, B2 => n307_port, ZN => n1273);
   U1329 : AOI22_X1 port map( A1 => REG_8_9_port, A2 => n361, B1 => 
                           REG_10_9_port, B2 => n343, ZN => n1272);
   U1330 : NAND4_X1 port map( A1 => n1275, A2 => n1274, A3 => n1273, A4 => 
                           n1272, ZN => n1276);
   U1331 : AOI22_X1 port map( A1 => n1277, A2 => n86, B1 => n1276, B2 => n84, 
                           ZN => n1278);
   U1332 : OAI221_X1 port map( B1 => n1743, B2 => n1280, C1 => n1741, C2 => 
                           n1279, A => n1278, ZN => N306);
   U1333 : AOI22_X1 port map( A1 => REG_21_10_port, A2 => n253_port, B1 => 
                           REG_23_10_port, B2 => n235_port, ZN => n1284);
   U1334 : AOI22_X1 port map( A1 => REG_17_10_port, A2 => n289_port, B1 => 
                           REG_19_10_port, B2 => n271_port, ZN => n1283);
   U1335 : AOI22_X1 port map( A1 => REG_20_10_port, A2 => n325, B1 => 
                           REG_22_10_port, B2 => n307_port, ZN => n1282);
   U1336 : AOI22_X1 port map( A1 => REG_16_10_port, A2 => n361, B1 => 
                           REG_18_10_port, B2 => n343, ZN => n1281);
   U1337 : AND4_X1 port map( A1 => n1284, A2 => n1283, A3 => n1282, A4 => n1281
                           , ZN => n1301);
   U1338 : AOI22_X1 port map( A1 => REG_29_10_port, A2 => n253_port, B1 => 
                           REG_31_10_port, B2 => n235_port, ZN => n1288);
   U1339 : AOI22_X1 port map( A1 => REG_25_10_port, A2 => n289_port, B1 => 
                           REG_27_10_port, B2 => n271_port, ZN => n1287);
   U1340 : AOI22_X1 port map( A1 => REG_28_10_port, A2 => n325, B1 => 
                           REG_30_10_port, B2 => n307_port, ZN => n1286);
   U1341 : AOI22_X1 port map( A1 => REG_24_10_port, A2 => n361, B1 => 
                           REG_26_10_port, B2 => n343, ZN => n1285);
   U1342 : AND4_X1 port map( A1 => n1288, A2 => n1287, A3 => n1286, A4 => n1285
                           , ZN => n1300);
   U1343 : AOI22_X1 port map( A1 => REG_5_10_port, A2 => n253_port, B1 => 
                           REG_7_10_port, B2 => n235_port, ZN => n1292);
   U1344 : AOI22_X1 port map( A1 => REG_1_10_port, A2 => n289_port, B1 => 
                           REG_3_10_port, B2 => n271_port, ZN => n1291);
   U1345 : AOI22_X1 port map( A1 => REG_4_10_port, A2 => n325, B1 => 
                           REG_6_10_port, B2 => n307_port, ZN => n1290);
   U1346 : AOI22_X1 port map( A1 => REG_0_10_port, A2 => n361, B1 => 
                           REG_2_10_port, B2 => n343, ZN => n1289);
   U1347 : NAND4_X1 port map( A1 => n1292, A2 => n1291, A3 => n1290, A4 => 
                           n1289, ZN => n1298);
   U1348 : AOI22_X1 port map( A1 => REG_13_10_port, A2 => n253_port, B1 => 
                           REG_15_10_port, B2 => n235_port, ZN => n1296);
   U1349 : AOI22_X1 port map( A1 => REG_9_10_port, A2 => n289_port, B1 => 
                           REG_11_10_port, B2 => n271_port, ZN => n1295);
   U1350 : AOI22_X1 port map( A1 => REG_12_10_port, A2 => n325, B1 => 
                           REG_14_10_port, B2 => n307_port, ZN => n1294);
   U1351 : AOI22_X1 port map( A1 => REG_8_10_port, A2 => n361, B1 => 
                           REG_10_10_port, B2 => n343, ZN => n1293);
   U1352 : NAND4_X1 port map( A1 => n1296, A2 => n1295, A3 => n1294, A4 => 
                           n1293, ZN => n1297);
   U1353 : AOI22_X1 port map( A1 => n1298, A2 => n86, B1 => n1297, B2 => n84, 
                           ZN => n1299);
   U1354 : OAI221_X1 port map( B1 => n1743, B2 => n1301, C1 => n1741, C2 => 
                           n1300, A => n1299, ZN => N305);
   U1355 : AOI22_X1 port map( A1 => REG_21_11_port, A2 => n254_port, B1 => 
                           REG_23_11_port, B2 => n236_port, ZN => n1305);
   U1356 : AOI22_X1 port map( A1 => REG_17_11_port, A2 => n290_port, B1 => 
                           REG_19_11_port, B2 => n272_port, ZN => n1304);
   U1357 : AOI22_X1 port map( A1 => REG_20_11_port, A2 => n326, B1 => 
                           REG_22_11_port, B2 => n308_port, ZN => n1303);
   U1358 : AOI22_X1 port map( A1 => REG_16_11_port, A2 => n362, B1 => 
                           REG_18_11_port, B2 => n344, ZN => n1302);
   U1359 : AND4_X1 port map( A1 => n1305, A2 => n1304, A3 => n1303, A4 => n1302
                           , ZN => n1322);
   U1360 : AOI22_X1 port map( A1 => REG_29_11_port, A2 => n254_port, B1 => 
                           REG_31_11_port, B2 => n236_port, ZN => n1309);
   U1361 : AOI22_X1 port map( A1 => REG_25_11_port, A2 => n290_port, B1 => 
                           REG_27_11_port, B2 => n272_port, ZN => n1308);
   U1362 : AOI22_X1 port map( A1 => REG_28_11_port, A2 => n326, B1 => 
                           REG_30_11_port, B2 => n308_port, ZN => n1307);
   U1363 : AOI22_X1 port map( A1 => REG_24_11_port, A2 => n362, B1 => 
                           REG_26_11_port, B2 => n344, ZN => n1306);
   U1364 : AND4_X1 port map( A1 => n1309, A2 => n1308, A3 => n1307, A4 => n1306
                           , ZN => n1321);
   U1365 : AOI22_X1 port map( A1 => REG_5_11_port, A2 => n254_port, B1 => 
                           REG_7_11_port, B2 => n236_port, ZN => n1313);
   U1366 : AOI22_X1 port map( A1 => REG_1_11_port, A2 => n290_port, B1 => 
                           REG_3_11_port, B2 => n272_port, ZN => n1312);
   U1367 : AOI22_X1 port map( A1 => REG_4_11_port, A2 => n326, B1 => 
                           REG_6_11_port, B2 => n308_port, ZN => n1311);
   U1368 : AOI22_X1 port map( A1 => REG_0_11_port, A2 => n362, B1 => 
                           REG_2_11_port, B2 => n344, ZN => n1310);
   U1369 : NAND4_X1 port map( A1 => n1313, A2 => n1312, A3 => n1311, A4 => 
                           n1310, ZN => n1319);
   U1370 : AOI22_X1 port map( A1 => REG_13_11_port, A2 => n254_port, B1 => 
                           REG_15_11_port, B2 => n236_port, ZN => n1317);
   U1371 : AOI22_X1 port map( A1 => REG_9_11_port, A2 => n290_port, B1 => 
                           REG_11_11_port, B2 => n272_port, ZN => n1316);
   U1372 : AOI22_X1 port map( A1 => REG_12_11_port, A2 => n326, B1 => 
                           REG_14_11_port, B2 => n308_port, ZN => n1315);
   U1373 : AOI22_X1 port map( A1 => REG_8_11_port, A2 => n362, B1 => 
                           REG_10_11_port, B2 => n344, ZN => n1314);
   U1374 : NAND4_X1 port map( A1 => n1317, A2 => n1316, A3 => n1315, A4 => 
                           n1314, ZN => n1318);
   U1375 : AOI22_X1 port map( A1 => n1319, A2 => n86, B1 => n1318, B2 => n84, 
                           ZN => n1320);
   U1376 : OAI221_X1 port map( B1 => n1743, B2 => n1322, C1 => n1741, C2 => 
                           n1321, A => n1320, ZN => N304);
   U1377 : AOI22_X1 port map( A1 => REG_21_12_port, A2 => n254_port, B1 => 
                           REG_23_12_port, B2 => n236_port, ZN => n1326);
   U1378 : AOI22_X1 port map( A1 => REG_17_12_port, A2 => n290_port, B1 => 
                           REG_19_12_port, B2 => n272_port, ZN => n1325);
   U1379 : AOI22_X1 port map( A1 => REG_20_12_port, A2 => n326, B1 => 
                           REG_22_12_port, B2 => n308_port, ZN => n1324);
   U1380 : AOI22_X1 port map( A1 => REG_16_12_port, A2 => n362, B1 => 
                           REG_18_12_port, B2 => n344, ZN => n1323);
   U1381 : AND4_X1 port map( A1 => n1326, A2 => n1325, A3 => n1324, A4 => n1323
                           , ZN => n1343);
   U1382 : AOI22_X1 port map( A1 => REG_29_12_port, A2 => n254_port, B1 => 
                           REG_31_12_port, B2 => n236_port, ZN => n1330);
   U1383 : AOI22_X1 port map( A1 => REG_25_12_port, A2 => n290_port, B1 => 
                           REG_27_12_port, B2 => n272_port, ZN => n1329);
   U1384 : AOI22_X1 port map( A1 => REG_28_12_port, A2 => n326, B1 => 
                           REG_30_12_port, B2 => n308_port, ZN => n1328);
   U1385 : AOI22_X1 port map( A1 => REG_24_12_port, A2 => n362, B1 => 
                           REG_26_12_port, B2 => n344, ZN => n1327);
   U1386 : AND4_X1 port map( A1 => n1330, A2 => n1329, A3 => n1328, A4 => n1327
                           , ZN => n1342);
   U1387 : AOI22_X1 port map( A1 => REG_5_12_port, A2 => n254_port, B1 => 
                           REG_7_12_port, B2 => n236_port, ZN => n1334);
   U1388 : AOI22_X1 port map( A1 => REG_1_12_port, A2 => n290_port, B1 => 
                           REG_3_12_port, B2 => n272_port, ZN => n1333);
   U1389 : AOI22_X1 port map( A1 => REG_4_12_port, A2 => n326, B1 => 
                           REG_6_12_port, B2 => n308_port, ZN => n1332);
   U1390 : AOI22_X1 port map( A1 => REG_0_12_port, A2 => n362, B1 => 
                           REG_2_12_port, B2 => n344, ZN => n1331);
   U1391 : NAND4_X1 port map( A1 => n1334, A2 => n1333, A3 => n1332, A4 => 
                           n1331, ZN => n1340);
   U1392 : AOI22_X1 port map( A1 => REG_13_12_port, A2 => n254_port, B1 => 
                           REG_15_12_port, B2 => n236_port, ZN => n1338);
   U1393 : AOI22_X1 port map( A1 => REG_9_12_port, A2 => n290_port, B1 => 
                           REG_11_12_port, B2 => n272_port, ZN => n1337);
   U1394 : AOI22_X1 port map( A1 => REG_12_12_port, A2 => n326, B1 => 
                           REG_14_12_port, B2 => n308_port, ZN => n1336);
   U1395 : AOI22_X1 port map( A1 => REG_8_12_port, A2 => n362, B1 => 
                           REG_10_12_port, B2 => n344, ZN => n1335);
   U1396 : NAND4_X1 port map( A1 => n1338, A2 => n1337, A3 => n1336, A4 => 
                           n1335, ZN => n1339);
   U1397 : AOI22_X1 port map( A1 => n1340, A2 => n86, B1 => n1339, B2 => n84, 
                           ZN => n1341);
   U1398 : OAI221_X1 port map( B1 => n1743, B2 => n1343, C1 => n1741, C2 => 
                           n1342, A => n1341, ZN => N303);
   U1399 : AOI22_X1 port map( A1 => REG_21_13_port, A2 => n254_port, B1 => 
                           REG_23_13_port, B2 => n236_port, ZN => n1347);
   U1400 : AOI22_X1 port map( A1 => REG_17_13_port, A2 => n290_port, B1 => 
                           REG_19_13_port, B2 => n272_port, ZN => n1346);
   U1401 : AOI22_X1 port map( A1 => REG_20_13_port, A2 => n326, B1 => 
                           REG_22_13_port, B2 => n308_port, ZN => n1345);
   U1402 : AOI22_X1 port map( A1 => REG_16_13_port, A2 => n362, B1 => 
                           REG_18_13_port, B2 => n344, ZN => n1344);
   U1403 : AND4_X1 port map( A1 => n1347, A2 => n1346, A3 => n1345, A4 => n1344
                           , ZN => n1364);
   U1404 : AOI22_X1 port map( A1 => REG_29_13_port, A2 => n254_port, B1 => 
                           REG_31_13_port, B2 => n236_port, ZN => n1351);
   U1405 : AOI22_X1 port map( A1 => REG_25_13_port, A2 => n290_port, B1 => 
                           REG_27_13_port, B2 => n272_port, ZN => n1350);
   U1406 : AOI22_X1 port map( A1 => REG_28_13_port, A2 => n326, B1 => 
                           REG_30_13_port, B2 => n308_port, ZN => n1349);
   U1407 : AOI22_X1 port map( A1 => REG_24_13_port, A2 => n362, B1 => 
                           REG_26_13_port, B2 => n344, ZN => n1348);
   U1408 : AND4_X1 port map( A1 => n1351, A2 => n1350, A3 => n1349, A4 => n1348
                           , ZN => n1363);
   U1409 : AOI22_X1 port map( A1 => REG_5_13_port, A2 => n254_port, B1 => 
                           REG_7_13_port, B2 => n236_port, ZN => n1355);
   U1410 : AOI22_X1 port map( A1 => REG_1_13_port, A2 => n290_port, B1 => 
                           REG_3_13_port, B2 => n272_port, ZN => n1354);
   U1411 : AOI22_X1 port map( A1 => REG_4_13_port, A2 => n326, B1 => 
                           REG_6_13_port, B2 => n308_port, ZN => n1353);
   U1412 : AOI22_X1 port map( A1 => REG_0_13_port, A2 => n362, B1 => 
                           REG_2_13_port, B2 => n344, ZN => n1352);
   U1413 : NAND4_X1 port map( A1 => n1355, A2 => n1354, A3 => n1353, A4 => 
                           n1352, ZN => n1361);
   U1414 : AOI22_X1 port map( A1 => REG_13_13_port, A2 => n255_port, B1 => 
                           REG_15_13_port, B2 => n237_port, ZN => n1359);
   U1415 : AOI22_X1 port map( A1 => REG_9_13_port, A2 => n291_port, B1 => 
                           REG_11_13_port, B2 => n273_port, ZN => n1358);
   U1416 : AOI22_X1 port map( A1 => REG_12_13_port, A2 => n327, B1 => 
                           REG_14_13_port, B2 => n309_port, ZN => n1357);
   U1417 : AOI22_X1 port map( A1 => REG_8_13_port, A2 => n363, B1 => 
                           REG_10_13_port, B2 => n345, ZN => n1356);
   U1418 : NAND4_X1 port map( A1 => n1359, A2 => n1358, A3 => n1357, A4 => 
                           n1356, ZN => n1360);
   U1419 : AOI22_X1 port map( A1 => n1361, A2 => n86, B1 => n1360, B2 => n84, 
                           ZN => n1362);
   U1420 : OAI221_X1 port map( B1 => n1743, B2 => n1364, C1 => n1741, C2 => 
                           n1363, A => n1362, ZN => N302);
   U1421 : AOI22_X1 port map( A1 => REG_21_14_port, A2 => n255_port, B1 => 
                           REG_23_14_port, B2 => n237_port, ZN => n1368);
   U1422 : AOI22_X1 port map( A1 => REG_17_14_port, A2 => n291_port, B1 => 
                           REG_19_14_port, B2 => n273_port, ZN => n1367);
   U1423 : AOI22_X1 port map( A1 => REG_20_14_port, A2 => n327, B1 => 
                           REG_22_14_port, B2 => n309_port, ZN => n1366);
   U1424 : AOI22_X1 port map( A1 => REG_16_14_port, A2 => n363, B1 => 
                           REG_18_14_port, B2 => n345, ZN => n1365);
   U1425 : AND4_X1 port map( A1 => n1368, A2 => n1367, A3 => n1366, A4 => n1365
                           , ZN => n1385);
   U1426 : AOI22_X1 port map( A1 => REG_29_14_port, A2 => n255_port, B1 => 
                           REG_31_14_port, B2 => n237_port, ZN => n1372);
   U1427 : AOI22_X1 port map( A1 => REG_25_14_port, A2 => n291_port, B1 => 
                           REG_27_14_port, B2 => n273_port, ZN => n1371);
   U1428 : AOI22_X1 port map( A1 => REG_28_14_port, A2 => n327, B1 => 
                           REG_30_14_port, B2 => n309_port, ZN => n1370);
   U1429 : AOI22_X1 port map( A1 => REG_24_14_port, A2 => n363, B1 => 
                           REG_26_14_port, B2 => n345, ZN => n1369);
   U1430 : AND4_X1 port map( A1 => n1372, A2 => n1371, A3 => n1370, A4 => n1369
                           , ZN => n1384);
   U1431 : AOI22_X1 port map( A1 => REG_5_14_port, A2 => n255_port, B1 => 
                           REG_7_14_port, B2 => n237_port, ZN => n1376);
   U1432 : AOI22_X1 port map( A1 => REG_1_14_port, A2 => n291_port, B1 => 
                           REG_3_14_port, B2 => n273_port, ZN => n1375);
   U1433 : AOI22_X1 port map( A1 => REG_4_14_port, A2 => n327, B1 => 
                           REG_6_14_port, B2 => n309_port, ZN => n1374);
   U1434 : AOI22_X1 port map( A1 => REG_0_14_port, A2 => n363, B1 => 
                           REG_2_14_port, B2 => n345, ZN => n1373);
   U1435 : NAND4_X1 port map( A1 => n1376, A2 => n1375, A3 => n1374, A4 => 
                           n1373, ZN => n1382);
   U1436 : AOI22_X1 port map( A1 => REG_13_14_port, A2 => n255_port, B1 => 
                           REG_15_14_port, B2 => n237_port, ZN => n1380);
   U1437 : AOI22_X1 port map( A1 => REG_9_14_port, A2 => n291_port, B1 => 
                           REG_11_14_port, B2 => n273_port, ZN => n1379);
   U1438 : AOI22_X1 port map( A1 => REG_12_14_port, A2 => n327, B1 => 
                           REG_14_14_port, B2 => n309_port, ZN => n1378);
   U1439 : AOI22_X1 port map( A1 => REG_8_14_port, A2 => n363, B1 => 
                           REG_10_14_port, B2 => n345, ZN => n1377);
   U1440 : NAND4_X1 port map( A1 => n1380, A2 => n1379, A3 => n1378, A4 => 
                           n1377, ZN => n1381);
   U1441 : AOI22_X1 port map( A1 => n1382, A2 => n86, B1 => n1381, B2 => n84, 
                           ZN => n1383);
   U1442 : OAI221_X1 port map( B1 => n1743, B2 => n1385, C1 => n1741, C2 => 
                           n1384, A => n1383, ZN => N301);
   U1443 : AOI22_X1 port map( A1 => REG_21_15_port, A2 => n255_port, B1 => 
                           REG_23_15_port, B2 => n237_port, ZN => n1389);
   U1444 : AOI22_X1 port map( A1 => REG_17_15_port, A2 => n291_port, B1 => 
                           REG_19_15_port, B2 => n273_port, ZN => n1388);
   U1445 : AOI22_X1 port map( A1 => REG_20_15_port, A2 => n327, B1 => 
                           REG_22_15_port, B2 => n309_port, ZN => n1387);
   U1446 : AOI22_X1 port map( A1 => REG_16_15_port, A2 => n363, B1 => 
                           REG_18_15_port, B2 => n345, ZN => n1386);
   U1447 : AND4_X1 port map( A1 => n1389, A2 => n1388, A3 => n1387, A4 => n1386
                           , ZN => n1406);
   U1448 : AOI22_X1 port map( A1 => REG_29_15_port, A2 => n255_port, B1 => 
                           REG_31_15_port, B2 => n237_port, ZN => n1393);
   U1449 : AOI22_X1 port map( A1 => REG_25_15_port, A2 => n291_port, B1 => 
                           REG_27_15_port, B2 => n273_port, ZN => n1392);
   U1450 : AOI22_X1 port map( A1 => REG_28_15_port, A2 => n327, B1 => 
                           REG_30_15_port, B2 => n309_port, ZN => n1391);
   U1451 : AOI22_X1 port map( A1 => REG_24_15_port, A2 => n363, B1 => 
                           REG_26_15_port, B2 => n345, ZN => n1390);
   U1452 : AND4_X1 port map( A1 => n1393, A2 => n1392, A3 => n1391, A4 => n1390
                           , ZN => n1405);
   U1453 : AOI22_X1 port map( A1 => REG_5_15_port, A2 => n255_port, B1 => 
                           REG_7_15_port, B2 => n237_port, ZN => n1397);
   U1454 : AOI22_X1 port map( A1 => REG_1_15_port, A2 => n291_port, B1 => 
                           REG_3_15_port, B2 => n273_port, ZN => n1396);
   U1455 : AOI22_X1 port map( A1 => REG_4_15_port, A2 => n327, B1 => 
                           REG_6_15_port, B2 => n309_port, ZN => n1395);
   U1456 : AOI22_X1 port map( A1 => REG_0_15_port, A2 => n363, B1 => 
                           REG_2_15_port, B2 => n345, ZN => n1394);
   U1457 : NAND4_X1 port map( A1 => n1397, A2 => n1396, A3 => n1395, A4 => 
                           n1394, ZN => n1403);
   U1458 : AOI22_X1 port map( A1 => REG_13_15_port, A2 => n255_port, B1 => 
                           REG_15_15_port, B2 => n237_port, ZN => n1401);
   U1459 : AOI22_X1 port map( A1 => REG_9_15_port, A2 => n291_port, B1 => 
                           REG_11_15_port, B2 => n273_port, ZN => n1400);
   U1460 : AOI22_X1 port map( A1 => REG_12_15_port, A2 => n327, B1 => 
                           REG_14_15_port, B2 => n309_port, ZN => n1399);
   U1461 : AOI22_X1 port map( A1 => REG_8_15_port, A2 => n363, B1 => 
                           REG_10_15_port, B2 => n345, ZN => n1398);
   U1462 : NAND4_X1 port map( A1 => n1401, A2 => n1400, A3 => n1399, A4 => 
                           n1398, ZN => n1402);
   U1463 : AOI22_X1 port map( A1 => n1403, A2 => n86, B1 => n1402, B2 => n84, 
                           ZN => n1404);
   U1464 : OAI221_X1 port map( B1 => n1743, B2 => n1406, C1 => n1741, C2 => 
                           n1405, A => n1404, ZN => N300);
   U1465 : AOI22_X1 port map( A1 => REG_21_16_port, A2 => n255_port, B1 => 
                           REG_23_16_port, B2 => n237_port, ZN => n1410);
   U1466 : AOI22_X1 port map( A1 => REG_17_16_port, A2 => n291_port, B1 => 
                           REG_19_16_port, B2 => n273_port, ZN => n1409);
   U1467 : AOI22_X1 port map( A1 => REG_20_16_port, A2 => n327, B1 => 
                           REG_22_16_port, B2 => n309_port, ZN => n1408);
   U1468 : AOI22_X1 port map( A1 => REG_16_16_port, A2 => n363, B1 => 
                           REG_18_16_port, B2 => n345, ZN => n1407);
   U1469 : AND4_X1 port map( A1 => n1410, A2 => n1409, A3 => n1408, A4 => n1407
                           , ZN => n1427);
   U1470 : AOI22_X1 port map( A1 => REG_29_16_port, A2 => n255_port, B1 => 
                           REG_31_16_port, B2 => n237_port, ZN => n1414);
   U1471 : AOI22_X1 port map( A1 => REG_25_16_port, A2 => n291_port, B1 => 
                           REG_27_16_port, B2 => n273_port, ZN => n1413);
   U1472 : AOI22_X1 port map( A1 => REG_28_16_port, A2 => n327, B1 => 
                           REG_30_16_port, B2 => n309_port, ZN => n1412);
   U1473 : AOI22_X1 port map( A1 => REG_24_16_port, A2 => n363, B1 => 
                           REG_26_16_port, B2 => n345, ZN => n1411);
   U1474 : AND4_X1 port map( A1 => n1414, A2 => n1413, A3 => n1412, A4 => n1411
                           , ZN => n1426);
   U1475 : AOI22_X1 port map( A1 => REG_5_16_port, A2 => n256_port, B1 => 
                           REG_7_16_port, B2 => n238_port, ZN => n1418);
   U1476 : AOI22_X1 port map( A1 => REG_1_16_port, A2 => n292_port, B1 => 
                           REG_3_16_port, B2 => n274_port, ZN => n1417);
   U1477 : AOI22_X1 port map( A1 => REG_4_16_port, A2 => n328, B1 => 
                           REG_6_16_port, B2 => n310_port, ZN => n1416);
   U1478 : AOI22_X1 port map( A1 => REG_0_16_port, A2 => n364, B1 => 
                           REG_2_16_port, B2 => n346, ZN => n1415);
   U1479 : NAND4_X1 port map( A1 => n1418, A2 => n1417, A3 => n1416, A4 => 
                           n1415, ZN => n1424);
   U1480 : AOI22_X1 port map( A1 => REG_13_16_port, A2 => n256_port, B1 => 
                           REG_15_16_port, B2 => n238_port, ZN => n1422);
   U1481 : AOI22_X1 port map( A1 => REG_9_16_port, A2 => n292_port, B1 => 
                           REG_11_16_port, B2 => n274_port, ZN => n1421);
   U1482 : AOI22_X1 port map( A1 => REG_12_16_port, A2 => n328, B1 => 
                           REG_14_16_port, B2 => n310_port, ZN => n1420);
   U1483 : AOI22_X1 port map( A1 => REG_8_16_port, A2 => n364, B1 => 
                           REG_10_16_port, B2 => n346, ZN => n1419);
   U1484 : NAND4_X1 port map( A1 => n1422, A2 => n1421, A3 => n1420, A4 => 
                           n1419, ZN => n1423);
   U1485 : AOI22_X1 port map( A1 => n1424, A2 => n86, B1 => n1423, B2 => n84, 
                           ZN => n1425);
   U1486 : OAI221_X1 port map( B1 => n1743, B2 => n1427, C1 => n1741, C2 => 
                           n1426, A => n1425, ZN => N299);
   U1487 : AOI22_X1 port map( A1 => REG_21_17_port, A2 => n256_port, B1 => 
                           REG_23_17_port, B2 => n238_port, ZN => n1431);
   U1488 : AOI22_X1 port map( A1 => REG_17_17_port, A2 => n292_port, B1 => 
                           REG_19_17_port, B2 => n274_port, ZN => n1430);
   U1489 : AOI22_X1 port map( A1 => REG_20_17_port, A2 => n328, B1 => 
                           REG_22_17_port, B2 => n310_port, ZN => n1429);
   U1490 : AOI22_X1 port map( A1 => REG_16_17_port, A2 => n364, B1 => 
                           REG_18_17_port, B2 => n346, ZN => n1428);
   U1491 : AND4_X1 port map( A1 => n1431, A2 => n1430, A3 => n1429, A4 => n1428
                           , ZN => n1448);
   U1492 : AOI22_X1 port map( A1 => REG_29_17_port, A2 => n256_port, B1 => 
                           REG_31_17_port, B2 => n238_port, ZN => n1435);
   U1493 : AOI22_X1 port map( A1 => REG_25_17_port, A2 => n292_port, B1 => 
                           REG_27_17_port, B2 => n274_port, ZN => n1434);
   U1494 : AOI22_X1 port map( A1 => REG_28_17_port, A2 => n328, B1 => 
                           REG_30_17_port, B2 => n310_port, ZN => n1433);
   U1495 : AOI22_X1 port map( A1 => REG_24_17_port, A2 => n364, B1 => 
                           REG_26_17_port, B2 => n346, ZN => n1432);
   U1496 : AND4_X1 port map( A1 => n1435, A2 => n1434, A3 => n1433, A4 => n1432
                           , ZN => n1447);
   U1497 : AOI22_X1 port map( A1 => REG_5_17_port, A2 => n256_port, B1 => 
                           REG_7_17_port, B2 => n238_port, ZN => n1439);
   U1498 : AOI22_X1 port map( A1 => REG_1_17_port, A2 => n292_port, B1 => 
                           REG_3_17_port, B2 => n274_port, ZN => n1438);
   U1499 : AOI22_X1 port map( A1 => REG_4_17_port, A2 => n328, B1 => 
                           REG_6_17_port, B2 => n310_port, ZN => n1437);
   U1500 : AOI22_X1 port map( A1 => REG_0_17_port, A2 => n364, B1 => 
                           REG_2_17_port, B2 => n346, ZN => n1436);
   U1501 : NAND4_X1 port map( A1 => n1439, A2 => n1438, A3 => n1437, A4 => 
                           n1436, ZN => n1445);
   U1502 : AOI22_X1 port map( A1 => REG_13_17_port, A2 => n256_port, B1 => 
                           REG_15_17_port, B2 => n238_port, ZN => n1443);
   U1503 : AOI22_X1 port map( A1 => REG_9_17_port, A2 => n292_port, B1 => 
                           REG_11_17_port, B2 => n274_port, ZN => n1442);
   U1504 : AOI22_X1 port map( A1 => REG_12_17_port, A2 => n328, B1 => 
                           REG_14_17_port, B2 => n310_port, ZN => n1441);
   U1505 : AOI22_X1 port map( A1 => REG_8_17_port, A2 => n364, B1 => 
                           REG_10_17_port, B2 => n346, ZN => n1440);
   U1506 : NAND4_X1 port map( A1 => n1443, A2 => n1442, A3 => n1441, A4 => 
                           n1440, ZN => n1444);
   U1507 : AOI22_X1 port map( A1 => n1445, A2 => n86, B1 => n1444, B2 => n84, 
                           ZN => n1446);
   U1508 : OAI221_X1 port map( B1 => n1743, B2 => n1448, C1 => n1741, C2 => 
                           n1447, A => n1446, ZN => N298);
   U1509 : AOI22_X1 port map( A1 => REG_21_18_port, A2 => n256_port, B1 => 
                           REG_23_18_port, B2 => n238_port, ZN => n1452);
   U1510 : AOI22_X1 port map( A1 => REG_17_18_port, A2 => n292_port, B1 => 
                           REG_19_18_port, B2 => n274_port, ZN => n1451);
   U1511 : AOI22_X1 port map( A1 => REG_20_18_port, A2 => n328, B1 => 
                           REG_22_18_port, B2 => n310_port, ZN => n1450);
   U1512 : AOI22_X1 port map( A1 => REG_16_18_port, A2 => n364, B1 => 
                           REG_18_18_port, B2 => n346, ZN => n1449);
   U1513 : AND4_X1 port map( A1 => n1452, A2 => n1451, A3 => n1450, A4 => n1449
                           , ZN => n1469);
   U1514 : AOI22_X1 port map( A1 => REG_29_18_port, A2 => n256_port, B1 => 
                           REG_31_18_port, B2 => n238_port, ZN => n1456);
   U1515 : AOI22_X1 port map( A1 => REG_25_18_port, A2 => n292_port, B1 => 
                           REG_27_18_port, B2 => n274_port, ZN => n1455);
   U1516 : AOI22_X1 port map( A1 => REG_28_18_port, A2 => n328, B1 => 
                           REG_30_18_port, B2 => n310_port, ZN => n1454);
   U1517 : AOI22_X1 port map( A1 => REG_24_18_port, A2 => n364, B1 => 
                           REG_26_18_port, B2 => n346, ZN => n1453);
   U1518 : AND4_X1 port map( A1 => n1456, A2 => n1455, A3 => n1454, A4 => n1453
                           , ZN => n1468);
   U1519 : AOI22_X1 port map( A1 => REG_5_18_port, A2 => n256_port, B1 => 
                           REG_7_18_port, B2 => n238_port, ZN => n1460);
   U1520 : AOI22_X1 port map( A1 => REG_1_18_port, A2 => n292_port, B1 => 
                           REG_3_18_port, B2 => n274_port, ZN => n1459);
   U1521 : AOI22_X1 port map( A1 => REG_4_18_port, A2 => n328, B1 => 
                           REG_6_18_port, B2 => n310_port, ZN => n1458);
   U1522 : AOI22_X1 port map( A1 => REG_0_18_port, A2 => n364, B1 => 
                           REG_2_18_port, B2 => n346, ZN => n1457);
   U1523 : NAND4_X1 port map( A1 => n1460, A2 => n1459, A3 => n1458, A4 => 
                           n1457, ZN => n1466);
   U1524 : AOI22_X1 port map( A1 => REG_13_18_port, A2 => n256_port, B1 => 
                           REG_15_18_port, B2 => n238_port, ZN => n1464);
   U1525 : AOI22_X1 port map( A1 => REG_9_18_port, A2 => n292_port, B1 => 
                           REG_11_18_port, B2 => n274_port, ZN => n1463);
   U1526 : AOI22_X1 port map( A1 => REG_12_18_port, A2 => n328, B1 => 
                           REG_14_18_port, B2 => n310_port, ZN => n1462);
   U1527 : AOI22_X1 port map( A1 => REG_8_18_port, A2 => n364, B1 => 
                           REG_10_18_port, B2 => n346, ZN => n1461);
   U1528 : NAND4_X1 port map( A1 => n1464, A2 => n1463, A3 => n1462, A4 => 
                           n1461, ZN => n1465);
   U1529 : AOI22_X1 port map( A1 => n1466, A2 => n86, B1 => n1465, B2 => n84, 
                           ZN => n1467);
   U1530 : OAI221_X1 port map( B1 => n1743, B2 => n1469, C1 => n1741, C2 => 
                           n1468, A => n1467, ZN => N297);
   U1531 : AOI22_X1 port map( A1 => REG_21_19_port, A2 => n256_port, B1 => 
                           REG_23_19_port, B2 => n238_port, ZN => n1473);
   U1532 : AOI22_X1 port map( A1 => REG_17_19_port, A2 => n292_port, B1 => 
                           REG_19_19_port, B2 => n274_port, ZN => n1472);
   U1533 : AOI22_X1 port map( A1 => REG_20_19_port, A2 => n328, B1 => 
                           REG_22_19_port, B2 => n310_port, ZN => n1471);
   U1534 : AOI22_X1 port map( A1 => REG_16_19_port, A2 => n364, B1 => 
                           REG_18_19_port, B2 => n346, ZN => n1470);
   U1535 : AND4_X1 port map( A1 => n1473, A2 => n1472, A3 => n1471, A4 => n1470
                           , ZN => n1490);
   U1536 : AOI22_X1 port map( A1 => REG_29_19_port, A2 => n257_port, B1 => 
                           REG_31_19_port, B2 => n239_port, ZN => n1477);
   U1537 : AOI22_X1 port map( A1 => REG_25_19_port, A2 => n293_port, B1 => 
                           REG_27_19_port, B2 => n275_port, ZN => n1476);
   U1538 : AOI22_X1 port map( A1 => REG_28_19_port, A2 => n329, B1 => 
                           REG_30_19_port, B2 => n311_port, ZN => n1475);
   U1539 : AOI22_X1 port map( A1 => REG_24_19_port, A2 => n365, B1 => 
                           REG_26_19_port, B2 => n347, ZN => n1474);
   U1540 : AND4_X1 port map( A1 => n1477, A2 => n1476, A3 => n1475, A4 => n1474
                           , ZN => n1489);
   U1541 : AOI22_X1 port map( A1 => REG_5_19_port, A2 => n257_port, B1 => 
                           REG_7_19_port, B2 => n239_port, ZN => n1481);
   U1542 : AOI22_X1 port map( A1 => REG_1_19_port, A2 => n293_port, B1 => 
                           REG_3_19_port, B2 => n275_port, ZN => n1480);
   U1543 : AOI22_X1 port map( A1 => REG_4_19_port, A2 => n329, B1 => 
                           REG_6_19_port, B2 => n311_port, ZN => n1479);
   U1544 : AOI22_X1 port map( A1 => REG_0_19_port, A2 => n365, B1 => 
                           REG_2_19_port, B2 => n347, ZN => n1478);
   U1545 : NAND4_X1 port map( A1 => n1481, A2 => n1480, A3 => n1479, A4 => 
                           n1478, ZN => n1487);
   U1546 : AOI22_X1 port map( A1 => REG_13_19_port, A2 => n257_port, B1 => 
                           REG_15_19_port, B2 => n239_port, ZN => n1485);
   U1547 : AOI22_X1 port map( A1 => REG_9_19_port, A2 => n293_port, B1 => 
                           REG_11_19_port, B2 => n275_port, ZN => n1484);
   U1548 : AOI22_X1 port map( A1 => REG_12_19_port, A2 => n329, B1 => 
                           REG_14_19_port, B2 => n311_port, ZN => n1483);
   U1549 : AOI22_X1 port map( A1 => REG_8_19_port, A2 => n365, B1 => 
                           REG_10_19_port, B2 => n347, ZN => n1482);
   U1550 : NAND4_X1 port map( A1 => n1485, A2 => n1484, A3 => n1483, A4 => 
                           n1482, ZN => n1486);
   U1551 : AOI22_X1 port map( A1 => n1487, A2 => n86, B1 => n1486, B2 => n84, 
                           ZN => n1488);
   U1552 : OAI221_X1 port map( B1 => n1743, B2 => n1490, C1 => n1741, C2 => 
                           n1489, A => n1488, ZN => N296);
   U1553 : AOI22_X1 port map( A1 => REG_21_20_port, A2 => n257_port, B1 => 
                           REG_23_20_port, B2 => n239_port, ZN => n1494);
   U1554 : AOI22_X1 port map( A1 => REG_17_20_port, A2 => n293_port, B1 => 
                           REG_19_20_port, B2 => n275_port, ZN => n1493);
   U1555 : AOI22_X1 port map( A1 => REG_20_20_port, A2 => n329, B1 => 
                           REG_22_20_port, B2 => n311_port, ZN => n1492);
   U1556 : AOI22_X1 port map( A1 => REG_16_20_port, A2 => n365, B1 => 
                           REG_18_20_port, B2 => n347, ZN => n1491);
   U1557 : AND4_X1 port map( A1 => n1494, A2 => n1493, A3 => n1492, A4 => n1491
                           , ZN => n1511);
   U1558 : AOI22_X1 port map( A1 => REG_29_20_port, A2 => n257_port, B1 => 
                           REG_31_20_port, B2 => n239_port, ZN => n1498);
   U1559 : AOI22_X1 port map( A1 => REG_25_20_port, A2 => n293_port, B1 => 
                           REG_27_20_port, B2 => n275_port, ZN => n1497);
   U1560 : AOI22_X1 port map( A1 => REG_28_20_port, A2 => n329, B1 => 
                           REG_30_20_port, B2 => n311_port, ZN => n1496);
   U1561 : AOI22_X1 port map( A1 => REG_24_20_port, A2 => n365, B1 => 
                           REG_26_20_port, B2 => n347, ZN => n1495);
   U1562 : AND4_X1 port map( A1 => n1498, A2 => n1497, A3 => n1496, A4 => n1495
                           , ZN => n1510);
   U1563 : AOI22_X1 port map( A1 => REG_5_20_port, A2 => n257_port, B1 => 
                           REG_7_20_port, B2 => n239_port, ZN => n1502);
   U1564 : AOI22_X1 port map( A1 => REG_1_20_port, A2 => n293_port, B1 => 
                           REG_3_20_port, B2 => n275_port, ZN => n1501);
   U1565 : AOI22_X1 port map( A1 => REG_4_20_port, A2 => n329, B1 => 
                           REG_6_20_port, B2 => n311_port, ZN => n1500);
   U1566 : AOI22_X1 port map( A1 => REG_0_20_port, A2 => n365, B1 => 
                           REG_2_20_port, B2 => n347, ZN => n1499);
   U1567 : NAND4_X1 port map( A1 => n1502, A2 => n1501, A3 => n1500, A4 => 
                           n1499, ZN => n1508);
   U1568 : AOI22_X1 port map( A1 => REG_13_20_port, A2 => n257_port, B1 => 
                           REG_15_20_port, B2 => n239_port, ZN => n1506);
   U1569 : AOI22_X1 port map( A1 => REG_9_20_port, A2 => n293_port, B1 => 
                           REG_11_20_port, B2 => n275_port, ZN => n1505);
   U1570 : AOI22_X1 port map( A1 => REG_12_20_port, A2 => n329, B1 => 
                           REG_14_20_port, B2 => n311_port, ZN => n1504);
   U1571 : AOI22_X1 port map( A1 => REG_8_20_port, A2 => n365, B1 => 
                           REG_10_20_port, B2 => n347, ZN => n1503);
   U1572 : NAND4_X1 port map( A1 => n1506, A2 => n1505, A3 => n1504, A4 => 
                           n1503, ZN => n1507);
   U1573 : AOI22_X1 port map( A1 => n1508, A2 => n86, B1 => n1507, B2 => n84, 
                           ZN => n1509);
   U1574 : OAI221_X1 port map( B1 => n1743, B2 => n1511, C1 => n1741, C2 => 
                           n1510, A => n1509, ZN => N295);
   U1575 : AOI22_X1 port map( A1 => REG_21_21_port, A2 => n257_port, B1 => 
                           REG_23_21_port, B2 => n239_port, ZN => n1515);
   U1576 : AOI22_X1 port map( A1 => REG_17_21_port, A2 => n293_port, B1 => 
                           REG_19_21_port, B2 => n275_port, ZN => n1514);
   U1577 : AOI22_X1 port map( A1 => REG_20_21_port, A2 => n329, B1 => 
                           REG_22_21_port, B2 => n311_port, ZN => n1513);
   U1578 : AOI22_X1 port map( A1 => REG_16_21_port, A2 => n365, B1 => 
                           REG_18_21_port, B2 => n347, ZN => n1512);
   U1579 : AND4_X1 port map( A1 => n1515, A2 => n1514, A3 => n1513, A4 => n1512
                           , ZN => n1532);
   U1580 : AOI22_X1 port map( A1 => REG_29_21_port, A2 => n257_port, B1 => 
                           REG_31_21_port, B2 => n239_port, ZN => n1519);
   U1581 : AOI22_X1 port map( A1 => REG_25_21_port, A2 => n293_port, B1 => 
                           REG_27_21_port, B2 => n275_port, ZN => n1518);
   U1582 : AOI22_X1 port map( A1 => REG_28_21_port, A2 => n329, B1 => 
                           REG_30_21_port, B2 => n311_port, ZN => n1517);
   U1583 : AOI22_X1 port map( A1 => REG_24_21_port, A2 => n365, B1 => 
                           REG_26_21_port, B2 => n347, ZN => n1516);
   U1584 : AND4_X1 port map( A1 => n1519, A2 => n1518, A3 => n1517, A4 => n1516
                           , ZN => n1531);
   U1585 : AOI22_X1 port map( A1 => REG_5_21_port, A2 => n257_port, B1 => 
                           REG_7_21_port, B2 => n239_port, ZN => n1523);
   U1586 : AOI22_X1 port map( A1 => REG_1_21_port, A2 => n293_port, B1 => 
                           REG_3_21_port, B2 => n275_port, ZN => n1522);
   U1587 : AOI22_X1 port map( A1 => REG_4_21_port, A2 => n329, B1 => 
                           REG_6_21_port, B2 => n311_port, ZN => n1521);
   U1588 : AOI22_X1 port map( A1 => REG_0_21_port, A2 => n365, B1 => 
                           REG_2_21_port, B2 => n347, ZN => n1520);
   U1589 : NAND4_X1 port map( A1 => n1523, A2 => n1522, A3 => n1521, A4 => 
                           n1520, ZN => n1529);
   U1590 : AOI22_X1 port map( A1 => REG_13_21_port, A2 => n257_port, B1 => 
                           REG_15_21_port, B2 => n239_port, ZN => n1527);
   U1591 : AOI22_X1 port map( A1 => REG_9_21_port, A2 => n293_port, B1 => 
                           REG_11_21_port, B2 => n275_port, ZN => n1526);
   U1592 : AOI22_X1 port map( A1 => REG_12_21_port, A2 => n329, B1 => 
                           REG_14_21_port, B2 => n311_port, ZN => n1525);
   U1593 : AOI22_X1 port map( A1 => REG_8_21_port, A2 => n365, B1 => 
                           REG_10_21_port, B2 => n347, ZN => n1524);
   U1594 : NAND4_X1 port map( A1 => n1527, A2 => n1526, A3 => n1525, A4 => 
                           n1524, ZN => n1528);
   U1595 : AOI22_X1 port map( A1 => n1529, A2 => n86, B1 => n1528, B2 => n84, 
                           ZN => n1530);
   U1596 : OAI221_X1 port map( B1 => n1743, B2 => n1532, C1 => n1741, C2 => 
                           n1531, A => n1530, ZN => N294);
   U1597 : AOI22_X1 port map( A1 => REG_21_22_port, A2 => n258_port, B1 => 
                           REG_23_22_port, B2 => n240_port, ZN => n1536);
   U1598 : AOI22_X1 port map( A1 => REG_17_22_port, A2 => n294_port, B1 => 
                           REG_19_22_port, B2 => n276_port, ZN => n1535);
   U1599 : AOI22_X1 port map( A1 => REG_20_22_port, A2 => n330, B1 => 
                           REG_22_22_port, B2 => n312_port, ZN => n1534);
   U1600 : AOI22_X1 port map( A1 => REG_16_22_port, A2 => n366, B1 => 
                           REG_18_22_port, B2 => n348, ZN => n1533);
   U1601 : AND4_X1 port map( A1 => n1536, A2 => n1535, A3 => n1534, A4 => n1533
                           , ZN => n1553);
   U1602 : AOI22_X1 port map( A1 => REG_29_22_port, A2 => n258_port, B1 => 
                           REG_31_22_port, B2 => n240_port, ZN => n1540);
   U1603 : AOI22_X1 port map( A1 => REG_25_22_port, A2 => n294_port, B1 => 
                           REG_27_22_port, B2 => n276_port, ZN => n1539);
   U1604 : AOI22_X1 port map( A1 => REG_28_22_port, A2 => n330, B1 => 
                           REG_30_22_port, B2 => n312_port, ZN => n1538);
   U1605 : AOI22_X1 port map( A1 => REG_24_22_port, A2 => n366, B1 => 
                           REG_26_22_port, B2 => n348, ZN => n1537);
   U1606 : AND4_X1 port map( A1 => n1540, A2 => n1539, A3 => n1538, A4 => n1537
                           , ZN => n1552);
   U1607 : AOI22_X1 port map( A1 => REG_5_22_port, A2 => n258_port, B1 => 
                           REG_7_22_port, B2 => n240_port, ZN => n1544);
   U1608 : AOI22_X1 port map( A1 => REG_1_22_port, A2 => n294_port, B1 => 
                           REG_3_22_port, B2 => n276_port, ZN => n1543);
   U1609 : AOI22_X1 port map( A1 => REG_4_22_port, A2 => n330, B1 => 
                           REG_6_22_port, B2 => n312_port, ZN => n1542);
   U1610 : AOI22_X1 port map( A1 => REG_0_22_port, A2 => n366, B1 => 
                           REG_2_22_port, B2 => n348, ZN => n1541);
   U1611 : NAND4_X1 port map( A1 => n1544, A2 => n1543, A3 => n1542, A4 => 
                           n1541, ZN => n1550);
   U1612 : AOI22_X1 port map( A1 => REG_13_22_port, A2 => n258_port, B1 => 
                           REG_15_22_port, B2 => n240_port, ZN => n1548);
   U1613 : AOI22_X1 port map( A1 => REG_9_22_port, A2 => n294_port, B1 => 
                           REG_11_22_port, B2 => n276_port, ZN => n1547);
   U1614 : AOI22_X1 port map( A1 => REG_12_22_port, A2 => n330, B1 => 
                           REG_14_22_port, B2 => n312_port, ZN => n1546);
   U1615 : AOI22_X1 port map( A1 => REG_8_22_port, A2 => n366, B1 => 
                           REG_10_22_port, B2 => n348, ZN => n1545);
   U1616 : NAND4_X1 port map( A1 => n1548, A2 => n1547, A3 => n1546, A4 => 
                           n1545, ZN => n1549);
   U1617 : AOI22_X1 port map( A1 => n1550, A2 => n86, B1 => n1549, B2 => n84, 
                           ZN => n1551);
   U1618 : OAI221_X1 port map( B1 => n1743, B2 => n1553, C1 => n1741, C2 => 
                           n1552, A => n1551, ZN => N293);
   U1619 : AOI22_X1 port map( A1 => REG_21_23_port, A2 => n258_port, B1 => 
                           REG_23_23_port, B2 => n240_port, ZN => n1557);
   U1620 : AOI22_X1 port map( A1 => REG_17_23_port, A2 => n294_port, B1 => 
                           REG_19_23_port, B2 => n276_port, ZN => n1556);
   U1621 : AOI22_X1 port map( A1 => REG_20_23_port, A2 => n330, B1 => 
                           REG_22_23_port, B2 => n312_port, ZN => n1555);
   U1622 : AOI22_X1 port map( A1 => REG_16_23_port, A2 => n366, B1 => 
                           REG_18_23_port, B2 => n348, ZN => n1554);
   U1623 : AND4_X1 port map( A1 => n1557, A2 => n1556, A3 => n1555, A4 => n1554
                           , ZN => n1574);
   U1624 : AOI22_X1 port map( A1 => REG_29_23_port, A2 => n258_port, B1 => 
                           REG_31_23_port, B2 => n240_port, ZN => n1561);
   U1625 : AOI22_X1 port map( A1 => REG_25_23_port, A2 => n294_port, B1 => 
                           REG_27_23_port, B2 => n276_port, ZN => n1560);
   U1626 : AOI22_X1 port map( A1 => REG_28_23_port, A2 => n330, B1 => 
                           REG_30_23_port, B2 => n312_port, ZN => n1559);
   U1627 : AOI22_X1 port map( A1 => REG_24_23_port, A2 => n366, B1 => 
                           REG_26_23_port, B2 => n348, ZN => n1558);
   U1628 : AND4_X1 port map( A1 => n1561, A2 => n1560, A3 => n1559, A4 => n1558
                           , ZN => n1573);
   U1629 : AOI22_X1 port map( A1 => REG_5_23_port, A2 => n258_port, B1 => 
                           REG_7_23_port, B2 => n240_port, ZN => n1565);
   U1630 : AOI22_X1 port map( A1 => REG_1_23_port, A2 => n294_port, B1 => 
                           REG_3_23_port, B2 => n276_port, ZN => n1564);
   U1631 : AOI22_X1 port map( A1 => REG_4_23_port, A2 => n330, B1 => 
                           REG_6_23_port, B2 => n312_port, ZN => n1563);
   U1632 : AOI22_X1 port map( A1 => REG_0_23_port, A2 => n366, B1 => 
                           REG_2_23_port, B2 => n348, ZN => n1562);
   U1633 : NAND4_X1 port map( A1 => n1565, A2 => n1564, A3 => n1563, A4 => 
                           n1562, ZN => n1571);
   U1634 : AOI22_X1 port map( A1 => REG_13_23_port, A2 => n258_port, B1 => 
                           REG_15_23_port, B2 => n240_port, ZN => n1569);
   U1635 : AOI22_X1 port map( A1 => REG_9_23_port, A2 => n294_port, B1 => 
                           REG_11_23_port, B2 => n276_port, ZN => n1568);
   U1636 : AOI22_X1 port map( A1 => REG_12_23_port, A2 => n330, B1 => 
                           REG_14_23_port, B2 => n312_port, ZN => n1567);
   U1637 : AOI22_X1 port map( A1 => REG_8_23_port, A2 => n366, B1 => 
                           REG_10_23_port, B2 => n348, ZN => n1566);
   U1638 : NAND4_X1 port map( A1 => n1569, A2 => n1568, A3 => n1567, A4 => 
                           n1566, ZN => n1570);
   U1639 : AOI22_X1 port map( A1 => n1571, A2 => n86, B1 => n1570, B2 => n84, 
                           ZN => n1572);
   U1640 : OAI221_X1 port map( B1 => n1743, B2 => n1574, C1 => n1741, C2 => 
                           n1573, A => n1572, ZN => N292);
   U1641 : AOI22_X1 port map( A1 => REG_21_24_port, A2 => n258_port, B1 => 
                           REG_23_24_port, B2 => n240_port, ZN => n1578);
   U1642 : AOI22_X1 port map( A1 => REG_17_24_port, A2 => n294_port, B1 => 
                           REG_19_24_port, B2 => n276_port, ZN => n1577);
   U1643 : AOI22_X1 port map( A1 => REG_20_24_port, A2 => n330, B1 => 
                           REG_22_24_port, B2 => n312_port, ZN => n1576);
   U1644 : AOI22_X1 port map( A1 => REG_16_24_port, A2 => n366, B1 => 
                           REG_18_24_port, B2 => n348, ZN => n1575);
   U1645 : AND4_X1 port map( A1 => n1578, A2 => n1577, A3 => n1576, A4 => n1575
                           , ZN => n1595);
   U1646 : AOI22_X1 port map( A1 => REG_29_24_port, A2 => n258_port, B1 => 
                           REG_31_24_port, B2 => n240_port, ZN => n1582);
   U1647 : AOI22_X1 port map( A1 => REG_25_24_port, A2 => n294_port, B1 => 
                           REG_27_24_port, B2 => n276_port, ZN => n1581);
   U1648 : AOI22_X1 port map( A1 => REG_28_24_port, A2 => n330, B1 => 
                           REG_30_24_port, B2 => n312_port, ZN => n1580);
   U1649 : AOI22_X1 port map( A1 => REG_24_24_port, A2 => n366, B1 => 
                           REG_26_24_port, B2 => n348, ZN => n1579);
   U1650 : AND4_X1 port map( A1 => n1582, A2 => n1581, A3 => n1580, A4 => n1579
                           , ZN => n1594);
   U1651 : AOI22_X1 port map( A1 => REG_5_24_port, A2 => n258_port, B1 => 
                           REG_7_24_port, B2 => n240_port, ZN => n1586);
   U1652 : AOI22_X1 port map( A1 => REG_1_24_port, A2 => n294_port, B1 => 
                           REG_3_24_port, B2 => n276_port, ZN => n1585);
   U1653 : AOI22_X1 port map( A1 => REG_4_24_port, A2 => n330, B1 => 
                           REG_6_24_port, B2 => n312_port, ZN => n1584);
   U1654 : AOI22_X1 port map( A1 => REG_0_24_port, A2 => n366, B1 => 
                           REG_2_24_port, B2 => n348, ZN => n1583);
   U1655 : NAND4_X1 port map( A1 => n1586, A2 => n1585, A3 => n1584, A4 => 
                           n1583, ZN => n1592);
   U1656 : AOI22_X1 port map( A1 => REG_13_24_port, A2 => n259_port, B1 => 
                           REG_15_24_port, B2 => n241_port, ZN => n1590);
   U1657 : AOI22_X1 port map( A1 => REG_9_24_port, A2 => n295_port, B1 => 
                           REG_11_24_port, B2 => n277_port, ZN => n1589);
   U1658 : AOI22_X1 port map( A1 => REG_12_24_port, A2 => n331, B1 => 
                           REG_14_24_port, B2 => n313_port, ZN => n1588);
   U1659 : AOI22_X1 port map( A1 => REG_8_24_port, A2 => n367, B1 => 
                           REG_10_24_port, B2 => n349, ZN => n1587);
   U1660 : NAND4_X1 port map( A1 => n1590, A2 => n1589, A3 => n1588, A4 => 
                           n1587, ZN => n1591);
   U1661 : AOI22_X1 port map( A1 => n1592, A2 => n86, B1 => n1591, B2 => n84, 
                           ZN => n1593);
   U1662 : OAI221_X1 port map( B1 => n1743, B2 => n1595, C1 => n1741, C2 => 
                           n1594, A => n1593, ZN => N291);
   U1663 : AOI22_X1 port map( A1 => REG_21_25_port, A2 => n259_port, B1 => 
                           REG_23_25_port, B2 => n241_port, ZN => n1599);
   U1664 : AOI22_X1 port map( A1 => REG_17_25_port, A2 => n295_port, B1 => 
                           REG_19_25_port, B2 => n277_port, ZN => n1598);
   U1665 : AOI22_X1 port map( A1 => REG_20_25_port, A2 => n331, B1 => 
                           REG_22_25_port, B2 => n313_port, ZN => n1597);
   U1666 : AOI22_X1 port map( A1 => REG_16_25_port, A2 => n367, B1 => 
                           REG_18_25_port, B2 => n349, ZN => n1596);
   U1667 : AND4_X1 port map( A1 => n1599, A2 => n1598, A3 => n1597, A4 => n1596
                           , ZN => n1616);
   U1668 : AOI22_X1 port map( A1 => REG_29_25_port, A2 => n259_port, B1 => 
                           REG_31_25_port, B2 => n241_port, ZN => n1603);
   U1669 : AOI22_X1 port map( A1 => REG_25_25_port, A2 => n295_port, B1 => 
                           REG_27_25_port, B2 => n277_port, ZN => n1602);
   U1670 : AOI22_X1 port map( A1 => REG_28_25_port, A2 => n331, B1 => 
                           REG_30_25_port, B2 => n313_port, ZN => n1601);
   U1671 : AOI22_X1 port map( A1 => REG_24_25_port, A2 => n367, B1 => 
                           REG_26_25_port, B2 => n349, ZN => n1600);
   U1672 : AND4_X1 port map( A1 => n1603, A2 => n1602, A3 => n1601, A4 => n1600
                           , ZN => n1615);
   U1673 : AOI22_X1 port map( A1 => REG_5_25_port, A2 => n259_port, B1 => 
                           REG_7_25_port, B2 => n241_port, ZN => n1607);
   U1674 : AOI22_X1 port map( A1 => REG_1_25_port, A2 => n295_port, B1 => 
                           REG_3_25_port, B2 => n277_port, ZN => n1606);
   U1675 : AOI22_X1 port map( A1 => REG_4_25_port, A2 => n331, B1 => 
                           REG_6_25_port, B2 => n313_port, ZN => n1605);
   U1676 : AOI22_X1 port map( A1 => REG_0_25_port, A2 => n367, B1 => 
                           REG_2_25_port, B2 => n349, ZN => n1604);
   U1677 : NAND4_X1 port map( A1 => n1607, A2 => n1606, A3 => n1605, A4 => 
                           n1604, ZN => n1613);
   U1678 : AOI22_X1 port map( A1 => REG_13_25_port, A2 => n259_port, B1 => 
                           REG_15_25_port, B2 => n241_port, ZN => n1611);
   U1679 : AOI22_X1 port map( A1 => REG_9_25_port, A2 => n295_port, B1 => 
                           REG_11_25_port, B2 => n277_port, ZN => n1610);
   U1680 : AOI22_X1 port map( A1 => REG_12_25_port, A2 => n331, B1 => 
                           REG_14_25_port, B2 => n313_port, ZN => n1609);
   U1681 : AOI22_X1 port map( A1 => REG_8_25_port, A2 => n367, B1 => 
                           REG_10_25_port, B2 => n349, ZN => n1608);
   U1682 : NAND4_X1 port map( A1 => n1611, A2 => n1610, A3 => n1609, A4 => 
                           n1608, ZN => n1612);
   U1683 : AOI22_X1 port map( A1 => n1613, A2 => n86, B1 => n1612, B2 => n84, 
                           ZN => n1614);
   U1684 : OAI221_X1 port map( B1 => n1743, B2 => n1616, C1 => n1741, C2 => 
                           n1615, A => n1614, ZN => N290);
   U1685 : AOI22_X1 port map( A1 => REG_21_26_port, A2 => n259_port, B1 => 
                           REG_23_26_port, B2 => n241_port, ZN => n1620);
   U1686 : AOI22_X1 port map( A1 => REG_17_26_port, A2 => n295_port, B1 => 
                           REG_19_26_port, B2 => n277_port, ZN => n1619);
   U1687 : AOI22_X1 port map( A1 => REG_20_26_port, A2 => n331, B1 => 
                           REG_22_26_port, B2 => n313_port, ZN => n1618);
   U1688 : AOI22_X1 port map( A1 => REG_16_26_port, A2 => n367, B1 => 
                           REG_18_26_port, B2 => n349, ZN => n1617);
   U1689 : AND4_X1 port map( A1 => n1620, A2 => n1619, A3 => n1618, A4 => n1617
                           , ZN => n1637);
   U1690 : AOI22_X1 port map( A1 => REG_29_26_port, A2 => n259_port, B1 => 
                           REG_31_26_port, B2 => n241_port, ZN => n1624);
   U1691 : AOI22_X1 port map( A1 => REG_25_26_port, A2 => n295_port, B1 => 
                           REG_27_26_port, B2 => n277_port, ZN => n1623);
   U1692 : AOI22_X1 port map( A1 => REG_28_26_port, A2 => n331, B1 => 
                           REG_30_26_port, B2 => n313_port, ZN => n1622);
   U1693 : AOI22_X1 port map( A1 => REG_24_26_port, A2 => n367, B1 => 
                           REG_26_26_port, B2 => n349, ZN => n1621);
   U1694 : AND4_X1 port map( A1 => n1624, A2 => n1623, A3 => n1622, A4 => n1621
                           , ZN => n1636);
   U1695 : AOI22_X1 port map( A1 => REG_5_26_port, A2 => n259_port, B1 => 
                           REG_7_26_port, B2 => n241_port, ZN => n1628);
   U1696 : AOI22_X1 port map( A1 => REG_1_26_port, A2 => n295_port, B1 => 
                           REG_3_26_port, B2 => n277_port, ZN => n1627);
   U1697 : AOI22_X1 port map( A1 => REG_4_26_port, A2 => n331, B1 => 
                           REG_6_26_port, B2 => n313_port, ZN => n1626);
   U1698 : AOI22_X1 port map( A1 => REG_0_26_port, A2 => n367, B1 => 
                           REG_2_26_port, B2 => n349, ZN => n1625);
   U1699 : NAND4_X1 port map( A1 => n1628, A2 => n1627, A3 => n1626, A4 => 
                           n1625, ZN => n1634);
   U1700 : AOI22_X1 port map( A1 => REG_13_26_port, A2 => n259_port, B1 => 
                           REG_15_26_port, B2 => n241_port, ZN => n1632);
   U1701 : AOI22_X1 port map( A1 => REG_9_26_port, A2 => n295_port, B1 => 
                           REG_11_26_port, B2 => n277_port, ZN => n1631);
   U1702 : AOI22_X1 port map( A1 => REG_12_26_port, A2 => n331, B1 => 
                           REG_14_26_port, B2 => n313_port, ZN => n1630);
   U1703 : AOI22_X1 port map( A1 => REG_8_26_port, A2 => n367, B1 => 
                           REG_10_26_port, B2 => n349, ZN => n1629);
   U1704 : NAND4_X1 port map( A1 => n1632, A2 => n1631, A3 => n1630, A4 => 
                           n1629, ZN => n1633);
   U1705 : AOI22_X1 port map( A1 => n1634, A2 => n86, B1 => n1633, B2 => n84, 
                           ZN => n1635);
   U1706 : OAI221_X1 port map( B1 => n1743, B2 => n1637, C1 => n1741, C2 => 
                           n1636, A => n1635, ZN => N289);
   U1707 : AOI22_X1 port map( A1 => REG_21_27_port, A2 => n259_port, B1 => 
                           REG_23_27_port, B2 => n241_port, ZN => n1641);
   U1708 : AOI22_X1 port map( A1 => REG_17_27_port, A2 => n295_port, B1 => 
                           REG_19_27_port, B2 => n277_port, ZN => n1640);
   U1709 : AOI22_X1 port map( A1 => REG_20_27_port, A2 => n331, B1 => 
                           REG_22_27_port, B2 => n313_port, ZN => n1639);
   U1710 : AOI22_X1 port map( A1 => REG_16_27_port, A2 => n367, B1 => 
                           REG_18_27_port, B2 => n349, ZN => n1638);
   U1711 : AND4_X1 port map( A1 => n1641, A2 => n1640, A3 => n1639, A4 => n1638
                           , ZN => n1658);
   U1712 : AOI22_X1 port map( A1 => REG_29_27_port, A2 => n259_port, B1 => 
                           REG_31_27_port, B2 => n241_port, ZN => n1645);
   U1713 : AOI22_X1 port map( A1 => REG_25_27_port, A2 => n295_port, B1 => 
                           REG_27_27_port, B2 => n277_port, ZN => n1644);
   U1714 : AOI22_X1 port map( A1 => REG_28_27_port, A2 => n331, B1 => 
                           REG_30_27_port, B2 => n313_port, ZN => n1643);
   U1715 : AOI22_X1 port map( A1 => REG_24_27_port, A2 => n367, B1 => 
                           REG_26_27_port, B2 => n349, ZN => n1642);
   U1716 : AND4_X1 port map( A1 => n1645, A2 => n1644, A3 => n1643, A4 => n1642
                           , ZN => n1657);
   U1717 : AOI22_X1 port map( A1 => REG_5_27_port, A2 => n260_port, B1 => 
                           REG_7_27_port, B2 => n242_port, ZN => n1649);
   U1718 : AOI22_X1 port map( A1 => REG_1_27_port, A2 => n296_port, B1 => 
                           REG_3_27_port, B2 => n278_port, ZN => n1648);
   U1719 : AOI22_X1 port map( A1 => REG_4_27_port, A2 => n332, B1 => 
                           REG_6_27_port, B2 => n314_port, ZN => n1647);
   U1720 : AOI22_X1 port map( A1 => REG_0_27_port, A2 => n368, B1 => 
                           REG_2_27_port, B2 => n350, ZN => n1646);
   U1721 : NAND4_X1 port map( A1 => n1649, A2 => n1648, A3 => n1647, A4 => 
                           n1646, ZN => n1655);
   U1722 : AOI22_X1 port map( A1 => REG_13_27_port, A2 => n260_port, B1 => 
                           REG_15_27_port, B2 => n242_port, ZN => n1653);
   U1723 : AOI22_X1 port map( A1 => REG_9_27_port, A2 => n296_port, B1 => 
                           REG_11_27_port, B2 => n278_port, ZN => n1652);
   U1724 : AOI22_X1 port map( A1 => REG_12_27_port, A2 => n332, B1 => 
                           REG_14_27_port, B2 => n314_port, ZN => n1651);
   U1725 : AOI22_X1 port map( A1 => REG_8_27_port, A2 => n368, B1 => 
                           REG_10_27_port, B2 => n350, ZN => n1650);
   U1726 : NAND4_X1 port map( A1 => n1653, A2 => n1652, A3 => n1651, A4 => 
                           n1650, ZN => n1654);
   U1727 : AOI22_X1 port map( A1 => n1655, A2 => n86, B1 => n1654, B2 => n84, 
                           ZN => n1656);
   U1728 : OAI221_X1 port map( B1 => n1743, B2 => n1658, C1 => n1741, C2 => 
                           n1657, A => n1656, ZN => N288);
   U1729 : AOI22_X1 port map( A1 => REG_21_28_port, A2 => n260_port, B1 => 
                           REG_23_28_port, B2 => n242_port, ZN => n1662);
   U1730 : AOI22_X1 port map( A1 => REG_17_28_port, A2 => n296_port, B1 => 
                           REG_19_28_port, B2 => n278_port, ZN => n1661);
   U1731 : AOI22_X1 port map( A1 => REG_20_28_port, A2 => n332, B1 => 
                           REG_22_28_port, B2 => n314_port, ZN => n1660);
   U1732 : AOI22_X1 port map( A1 => REG_16_28_port, A2 => n368, B1 => 
                           REG_18_28_port, B2 => n350, ZN => n1659);
   U1733 : AND4_X1 port map( A1 => n1662, A2 => n1661, A3 => n1660, A4 => n1659
                           , ZN => n1679);
   U1734 : AOI22_X1 port map( A1 => REG_29_28_port, A2 => n260_port, B1 => 
                           REG_31_28_port, B2 => n242_port, ZN => n1666);
   U1735 : AOI22_X1 port map( A1 => REG_25_28_port, A2 => n296_port, B1 => 
                           REG_27_28_port, B2 => n278_port, ZN => n1665);
   U1736 : AOI22_X1 port map( A1 => REG_28_28_port, A2 => n332, B1 => 
                           REG_30_28_port, B2 => n314_port, ZN => n1664);
   U1737 : AOI22_X1 port map( A1 => REG_24_28_port, A2 => n368, B1 => 
                           REG_26_28_port, B2 => n350, ZN => n1663);
   U1738 : AND4_X1 port map( A1 => n1666, A2 => n1665, A3 => n1664, A4 => n1663
                           , ZN => n1678);
   U1739 : AOI22_X1 port map( A1 => REG_5_28_port, A2 => n260_port, B1 => 
                           REG_7_28_port, B2 => n242_port, ZN => n1670);
   U1740 : AOI22_X1 port map( A1 => REG_1_28_port, A2 => n296_port, B1 => 
                           REG_3_28_port, B2 => n278_port, ZN => n1669);
   U1741 : AOI22_X1 port map( A1 => REG_4_28_port, A2 => n332, B1 => 
                           REG_6_28_port, B2 => n314_port, ZN => n1668);
   U1742 : AOI22_X1 port map( A1 => REG_0_28_port, A2 => n368, B1 => 
                           REG_2_28_port, B2 => n350, ZN => n1667);
   U1743 : NAND4_X1 port map( A1 => n1670, A2 => n1669, A3 => n1668, A4 => 
                           n1667, ZN => n1676);
   U1744 : AOI22_X1 port map( A1 => REG_13_28_port, A2 => n260_port, B1 => 
                           REG_15_28_port, B2 => n242_port, ZN => n1674);
   U1745 : AOI22_X1 port map( A1 => REG_9_28_port, A2 => n296_port, B1 => 
                           REG_11_28_port, B2 => n278_port, ZN => n1673);
   U1746 : AOI22_X1 port map( A1 => REG_12_28_port, A2 => n332, B1 => 
                           REG_14_28_port, B2 => n314_port, ZN => n1672);
   U1747 : AOI22_X1 port map( A1 => REG_8_28_port, A2 => n368, B1 => 
                           REG_10_28_port, B2 => n350, ZN => n1671);
   U1748 : NAND4_X1 port map( A1 => n1674, A2 => n1673, A3 => n1672, A4 => 
                           n1671, ZN => n1675);
   U1749 : AOI22_X1 port map( A1 => n1676, A2 => n86, B1 => n1675, B2 => n84, 
                           ZN => n1677);
   U1750 : OAI221_X1 port map( B1 => n1743, B2 => n1679, C1 => n1741, C2 => 
                           n1678, A => n1677, ZN => N287);
   U1751 : AOI22_X1 port map( A1 => REG_21_29_port, A2 => n260_port, B1 => 
                           REG_23_29_port, B2 => n242_port, ZN => n1683);
   U1752 : AOI22_X1 port map( A1 => REG_17_29_port, A2 => n296_port, B1 => 
                           REG_19_29_port, B2 => n278_port, ZN => n1682);
   U1753 : AOI22_X1 port map( A1 => REG_20_29_port, A2 => n332, B1 => 
                           REG_22_29_port, B2 => n314_port, ZN => n1681);
   U1754 : AOI22_X1 port map( A1 => REG_16_29_port, A2 => n368, B1 => 
                           REG_18_29_port, B2 => n350, ZN => n1680);
   U1755 : AND4_X1 port map( A1 => n1683, A2 => n1682, A3 => n1681, A4 => n1680
                           , ZN => n1700);
   U1756 : AOI22_X1 port map( A1 => REG_29_29_port, A2 => n260_port, B1 => 
                           REG_31_29_port, B2 => n242_port, ZN => n1687);
   U1757 : AOI22_X1 port map( A1 => REG_25_29_port, A2 => n296_port, B1 => 
                           REG_27_29_port, B2 => n278_port, ZN => n1686);
   U1758 : AOI22_X1 port map( A1 => REG_28_29_port, A2 => n332, B1 => 
                           REG_30_29_port, B2 => n314_port, ZN => n1685);
   U1759 : AOI22_X1 port map( A1 => REG_24_29_port, A2 => n368, B1 => 
                           REG_26_29_port, B2 => n350, ZN => n1684);
   U1760 : AND4_X1 port map( A1 => n1687, A2 => n1686, A3 => n1685, A4 => n1684
                           , ZN => n1699);
   U1761 : AOI22_X1 port map( A1 => REG_5_29_port, A2 => n260_port, B1 => 
                           REG_7_29_port, B2 => n242_port, ZN => n1691);
   U1762 : AOI22_X1 port map( A1 => REG_1_29_port, A2 => n296_port, B1 => 
                           REG_3_29_port, B2 => n278_port, ZN => n1690);
   U1763 : AOI22_X1 port map( A1 => REG_4_29_port, A2 => n332, B1 => 
                           REG_6_29_port, B2 => n314_port, ZN => n1689);
   U1764 : AOI22_X1 port map( A1 => REG_0_29_port, A2 => n368, B1 => 
                           REG_2_29_port, B2 => n350, ZN => n1688);
   U1765 : NAND4_X1 port map( A1 => n1691, A2 => n1690, A3 => n1689, A4 => 
                           n1688, ZN => n1697);
   U1766 : AOI22_X1 port map( A1 => REG_13_29_port, A2 => n260_port, B1 => 
                           REG_15_29_port, B2 => n242_port, ZN => n1695);
   U1767 : AOI22_X1 port map( A1 => REG_9_29_port, A2 => n296_port, B1 => 
                           REG_11_29_port, B2 => n278_port, ZN => n1694);
   U1768 : AOI22_X1 port map( A1 => REG_12_29_port, A2 => n332, B1 => 
                           REG_14_29_port, B2 => n314_port, ZN => n1693);
   U1769 : AOI22_X1 port map( A1 => REG_8_29_port, A2 => n368, B1 => 
                           REG_10_29_port, B2 => n350, ZN => n1692);
   U1770 : NAND4_X1 port map( A1 => n1695, A2 => n1694, A3 => n1693, A4 => 
                           n1692, ZN => n1696);
   U1771 : AOI22_X1 port map( A1 => n1697, A2 => n86, B1 => n1696, B2 => n84, 
                           ZN => n1698);
   U1772 : OAI221_X1 port map( B1 => n1743, B2 => n1700, C1 => n1741, C2 => 
                           n1699, A => n1698, ZN => N286);
   U1773 : AOI22_X1 port map( A1 => REG_21_30_port, A2 => n260_port, B1 => 
                           REG_23_30_port, B2 => n242_port, ZN => n1704);
   U1774 : AOI22_X1 port map( A1 => REG_17_30_port, A2 => n296_port, B1 => 
                           REG_19_30_port, B2 => n278_port, ZN => n1703);
   U1775 : AOI22_X1 port map( A1 => REG_20_30_port, A2 => n332, B1 => 
                           REG_22_30_port, B2 => n314_port, ZN => n1702);
   U1776 : AOI22_X1 port map( A1 => REG_16_30_port, A2 => n368, B1 => 
                           REG_18_30_port, B2 => n350, ZN => n1701);
   U1777 : AND4_X1 port map( A1 => n1704, A2 => n1703, A3 => n1702, A4 => n1701
                           , ZN => n1721);
   U1778 : AOI22_X1 port map( A1 => REG_29_30_port, A2 => n261_port, B1 => 
                           REG_31_30_port, B2 => n243_port, ZN => n1708);
   U1779 : AOI22_X1 port map( A1 => REG_25_30_port, A2 => n297_port, B1 => 
                           REG_27_30_port, B2 => n279_port, ZN => n1707);
   U1780 : AOI22_X1 port map( A1 => REG_28_30_port, A2 => n333, B1 => 
                           REG_30_30_port, B2 => n315_port, ZN => n1706);
   U1781 : AOI22_X1 port map( A1 => REG_24_30_port, A2 => n369, B1 => 
                           REG_26_30_port, B2 => n351, ZN => n1705);
   U1782 : AND4_X1 port map( A1 => n1708, A2 => n1707, A3 => n1706, A4 => n1705
                           , ZN => n1720);
   U1783 : AOI22_X1 port map( A1 => REG_5_30_port, A2 => n261_port, B1 => 
                           REG_7_30_port, B2 => n243_port, ZN => n1712);
   U1784 : AOI22_X1 port map( A1 => REG_1_30_port, A2 => n297_port, B1 => 
                           REG_3_30_port, B2 => n279_port, ZN => n1711);
   U1785 : AOI22_X1 port map( A1 => REG_4_30_port, A2 => n333, B1 => 
                           REG_6_30_port, B2 => n315_port, ZN => n1710);
   U1786 : AOI22_X1 port map( A1 => REG_0_30_port, A2 => n369, B1 => 
                           REG_2_30_port, B2 => n351, ZN => n1709);
   U1787 : NAND4_X1 port map( A1 => n1712, A2 => n1711, A3 => n1710, A4 => 
                           n1709, ZN => n1718);
   U1788 : AOI22_X1 port map( A1 => REG_13_30_port, A2 => n261_port, B1 => 
                           REG_15_30_port, B2 => n243_port, ZN => n1716);
   U1789 : AOI22_X1 port map( A1 => REG_9_30_port, A2 => n297_port, B1 => 
                           REG_11_30_port, B2 => n279_port, ZN => n1715);
   U1790 : AOI22_X1 port map( A1 => REG_12_30_port, A2 => n333, B1 => 
                           REG_14_30_port, B2 => n315_port, ZN => n1714);
   U1791 : AOI22_X1 port map( A1 => REG_8_30_port, A2 => n369, B1 => 
                           REG_10_30_port, B2 => n351, ZN => n1713);
   U1792 : NAND4_X1 port map( A1 => n1716, A2 => n1715, A3 => n1714, A4 => 
                           n1713, ZN => n1717);
   U1793 : AOI22_X1 port map( A1 => n1718, A2 => n86, B1 => n1717, B2 => n84, 
                           ZN => n1719);
   U1794 : OAI221_X1 port map( B1 => n1743, B2 => n1721, C1 => n1741, C2 => 
                           n1720, A => n1719, ZN => N285);
   U1795 : AOI22_X1 port map( A1 => REG_21_31_port, A2 => n261_port, B1 => 
                           REG_23_31_port, B2 => n243_port, ZN => n1725);
   U1796 : AOI22_X1 port map( A1 => REG_17_31_port, A2 => n297_port, B1 => 
                           REG_19_31_port, B2 => n279_port, ZN => n1724);
   U1797 : AOI22_X1 port map( A1 => REG_20_31_port, A2 => n333, B1 => 
                           REG_22_31_port, B2 => n315_port, ZN => n1723);
   U1798 : AOI22_X1 port map( A1 => REG_16_31_port, A2 => n369, B1 => 
                           REG_18_31_port, B2 => n351, ZN => n1722);
   U1799 : AND4_X1 port map( A1 => n1725, A2 => n1724, A3 => n1723, A4 => n1722
                           , ZN => n1744);
   U1800 : AOI22_X1 port map( A1 => REG_29_31_port, A2 => n261_port, B1 => 
                           REG_31_31_port, B2 => n243_port, ZN => n1729);
   U1801 : AOI22_X1 port map( A1 => REG_25_31_port, A2 => n297_port, B1 => 
                           REG_27_31_port, B2 => n279_port, ZN => n1728);
   U1802 : AOI22_X1 port map( A1 => REG_28_31_port, A2 => n333, B1 => 
                           REG_30_31_port, B2 => n315_port, ZN => n1727);
   U1803 : AOI22_X1 port map( A1 => REG_24_31_port, A2 => n369, B1 => 
                           REG_26_31_port, B2 => n351, ZN => n1726);
   U1804 : AND4_X1 port map( A1 => n1729, A2 => n1728, A3 => n1727, A4 => n1726
                           , ZN => n1742);
   U1805 : AOI22_X1 port map( A1 => REG_5_31_port, A2 => n261_port, B1 => 
                           REG_7_31_port, B2 => n243_port, ZN => n1733);
   U1806 : AOI22_X1 port map( A1 => REG_1_31_port, A2 => n297_port, B1 => 
                           REG_3_31_port, B2 => n279_port, ZN => n1732);
   U1807 : AOI22_X1 port map( A1 => REG_4_31_port, A2 => n333, B1 => 
                           REG_6_31_port, B2 => n315_port, ZN => n1731);
   U1808 : AOI22_X1 port map( A1 => REG_0_31_port, A2 => n369, B1 => 
                           REG_2_31_port, B2 => n351, ZN => n1730);
   U1809 : NAND4_X1 port map( A1 => n1733, A2 => n1732, A3 => n1731, A4 => 
                           n1730, ZN => n1739);
   U1810 : AOI22_X1 port map( A1 => REG_13_31_port, A2 => n261_port, B1 => 
                           REG_15_31_port, B2 => n243_port, ZN => n1737);
   U1811 : AOI22_X1 port map( A1 => REG_9_31_port, A2 => n297_port, B1 => 
                           REG_11_31_port, B2 => n279_port, ZN => n1736);
   U1812 : AOI22_X1 port map( A1 => REG_12_31_port, A2 => n333, B1 => 
                           REG_14_31_port, B2 => n315_port, ZN => n1735);
   U1813 : AOI22_X1 port map( A1 => REG_8_31_port, A2 => n369, B1 => 
                           REG_10_31_port, B2 => n351, ZN => n1734);
   U1814 : NAND4_X1 port map( A1 => n1737, A2 => n1736, A3 => n1735, A4 => 
                           n1734, ZN => n1738);
   U1815 : AOI22_X1 port map( A1 => n86, A2 => n1739, B1 => n84, B2 => n1738, 
                           ZN => n1740);
   U1816 : OAI221_X1 port map( B1 => n1744, B2 => n1743, C1 => n1742, C2 => 
                           n1741, A => n1740, ZN => N284);
   U1817 : INV_X1 port map( A => n1749, ZN => n1801);
   U1818 : INV_X1 port map( A => n1750, ZN => n1802);
   U1819 : INV_X1 port map( A => n1751, ZN => n1803);
   U1820 : INV_X1 port map( A => n1752, ZN => n1804);
   U1821 : INV_X1 port map( A => n1753, ZN => n1805);
   U1822 : INV_X1 port map( A => n1754, ZN => n1806);
   U1823 : INV_X1 port map( A => n1755, ZN => n1807);
   U1824 : INV_X1 port map( A => n1756, ZN => n1808);
   U1825 : INV_X1 port map( A => n1757, ZN => n1809);
   U1826 : INV_X1 port map( A => n1758, ZN => n1810);
   U1827 : INV_X1 port map( A => n1759, ZN => n1811);
   U1828 : INV_X1 port map( A => n1760, ZN => n1812);
   U1829 : INV_X1 port map( A => n1761, ZN => n1813);
   U1830 : INV_X1 port map( A => n1762, ZN => n1814);
   U1831 : INV_X1 port map( A => n1763, ZN => n1815);
   U1832 : INV_X1 port map( A => n1764, ZN => n1816);
   U1833 : INV_X1 port map( A => n1765, ZN => n1817);
   U1834 : INV_X1 port map( A => n1766, ZN => n1818);
   U1835 : INV_X1 port map( A => n1767, ZN => n1819);
   U1836 : INV_X1 port map( A => n1768, ZN => n1820);
   U1837 : INV_X1 port map( A => n1769, ZN => n1821);
   U1838 : INV_X1 port map( A => n1770, ZN => n1822);
   U1839 : INV_X1 port map( A => n1771, ZN => n1823);
   U1840 : INV_X1 port map( A => n1772, ZN => n1824);
   U1841 : INV_X1 port map( A => n1773, ZN => n1825);
   U1842 : INV_X1 port map( A => n1774, ZN => n1826);
   U1843 : INV_X1 port map( A => n1775, ZN => n1827);
   U1844 : INV_X1 port map( A => n1776, ZN => n1828);
   U1845 : INV_X1 port map( A => n1777, ZN => n1829);
   U1846 : INV_X1 port map( A => n1778, ZN => n1830);
   U1847 : INV_X1 port map( A => n1779, ZN => n1831);
   U1848 : INV_X1 port map( A => n1780, ZN => n1832);
   U1849 : AND2_X1 port map( A1 => EN_RD2, A2 => EN, ZN => N317);
   U1850 : AND2_X1 port map( A1 => EN_RD1, A2 => EN, ZN => N316);
   U1851 : NOR2_X1 port map( A1 => n87, A2 => n1749, ZN => N250);
   U1852 : NAND2_X1 port map( A1 => n382, A2 => DATAIN(31), ZN => n1749);
   U1853 : NOR2_X1 port map( A1 => n87, A2 => n1750, ZN => N249);
   U1854 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n382, ZN => n1750);
   U1855 : NOR2_X1 port map( A1 => n87, A2 => n1751, ZN => N248);
   U1856 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n382, ZN => n1751);
   U1857 : NOR2_X1 port map( A1 => n87, A2 => n1752, ZN => N247);
   U1858 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n382, ZN => n1752);
   U1859 : NOR2_X1 port map( A1 => n87, A2 => n1753, ZN => N246);
   U1860 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n382, ZN => n1753);
   U1861 : NOR2_X1 port map( A1 => n87, A2 => n1754, ZN => N245);
   U1862 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n382, ZN => n1754);
   U1863 : NOR2_X1 port map( A1 => n87, A2 => n1755, ZN => N244);
   U1864 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n382, ZN => n1755);
   U1865 : NOR2_X1 port map( A1 => n87, A2 => n1756, ZN => N243);
   U1866 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n382, ZN => n1756);
   U1867 : NOR2_X1 port map( A1 => n87, A2 => n1757, ZN => N242);
   U1868 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n382, ZN => n1757);
   U1869 : NOR2_X1 port map( A1 => n87, A2 => n1758, ZN => N241);
   U1870 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n381, ZN => n1758);
   U1871 : NOR2_X1 port map( A1 => n87, A2 => n1759, ZN => N240);
   U1872 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n381, ZN => n1759);
   U1873 : NOR2_X1 port map( A1 => n87, A2 => n1760, ZN => N239);
   U1874 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n381, ZN => n1760);
   U1875 : NOR2_X1 port map( A1 => n87, A2 => n1761, ZN => N238);
   U1876 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n381, ZN => n1761);
   U1877 : NOR2_X1 port map( A1 => n87, A2 => n1762, ZN => N237);
   U1878 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n381, ZN => n1762);
   U1879 : NOR2_X1 port map( A1 => n87, A2 => n1763, ZN => N236);
   U1880 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n381, ZN => n1763);
   U1881 : NOR2_X1 port map( A1 => n87, A2 => n1764, ZN => N235);
   U1882 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n381, ZN => n1764);
   U1883 : NOR2_X1 port map( A1 => n87, A2 => n1765, ZN => N234);
   U1884 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n381, ZN => n1765);
   U1885 : NOR2_X1 port map( A1 => n87, A2 => n1766, ZN => N233);
   U1886 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n381, ZN => n1766);
   U1887 : NOR2_X1 port map( A1 => n87, A2 => n1767, ZN => N232);
   U1888 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n381, ZN => n1767);
   U1889 : NOR2_X1 port map( A1 => n87, A2 => n1768, ZN => N231);
   U1890 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n381, ZN => n1768);
   U1891 : NOR2_X1 port map( A1 => n87, A2 => n1769, ZN => N230);
   U1892 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n380, ZN => n1769);
   U1893 : NOR2_X1 port map( A1 => n87, A2 => n1770, ZN => N229);
   U1894 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n380, ZN => n1770);
   U1895 : NOR2_X1 port map( A1 => n87, A2 => n1771, ZN => N228);
   U1896 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n380, ZN => n1771);
   U1897 : NOR2_X1 port map( A1 => n87, A2 => n1772, ZN => N227);
   U1898 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n380, ZN => n1772);
   U1899 : NOR2_X1 port map( A1 => n87, A2 => n1773, ZN => N226);
   U1900 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n380, ZN => n1773);
   U1901 : NOR2_X1 port map( A1 => n87, A2 => n1774, ZN => N225);
   U1902 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n380, ZN => n1774);
   U1903 : NOR2_X1 port map( A1 => n87, A2 => n1775, ZN => N224);
   U1904 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n380, ZN => n1775);
   U1905 : NOR2_X1 port map( A1 => n87, A2 => n1776, ZN => N223);
   U1906 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n380, ZN => n1776);
   U1907 : NOR2_X1 port map( A1 => n87, A2 => n1777, ZN => N222);
   U1908 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n380, ZN => n1777);
   U1909 : NOR2_X1 port map( A1 => n87, A2 => n1778, ZN => N221);
   U1910 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n380, ZN => n1778);
   U1911 : NOR2_X1 port map( A1 => n87, A2 => n1779, ZN => N220);
   U1912 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n380, ZN => n1779);
   U1913 : NOR2_X1 port map( A1 => n87, A2 => n1780, ZN => N219);
   U1914 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n379, ZN => n1780);
   U1915 : OAI21_X1 port map( B1 => n1784, B2 => n1785, A => n379, ZN => N217);
   U1916 : OAI21_X1 port map( B1 => n1784, B2 => n1786, A => n379, ZN => N216);
   U1917 : OAI21_X1 port map( B1 => n1784, B2 => n1787, A => n379, ZN => N215);
   U1918 : OAI21_X1 port map( B1 => n1784, B2 => n1788, A => n379, ZN => N214);
   U1919 : OAI21_X1 port map( B1 => n1784, B2 => n1789, A => n379, ZN => N213);
   U1920 : OAI21_X1 port map( B1 => n1784, B2 => n1790, A => n379, ZN => N212);
   U1921 : OAI21_X1 port map( B1 => n1784, B2 => n1791, A => n379, ZN => N211);
   U1922 : NAND3_X1 port map( A1 => n1792, A2 => n1793, A3 => n1794, ZN => 
                           n1784);
   U1923 : OAI21_X1 port map( B1 => n1783, B2 => n1795, A => n379, ZN => N210);
   U1924 : OAI21_X1 port map( B1 => n1785, B2 => n1795, A => n379, ZN => N209);
   U1925 : OAI21_X1 port map( B1 => n1786, B2 => n1795, A => n378, ZN => N208);
   U1926 : OAI21_X1 port map( B1 => n1787, B2 => n1795, A => n378, ZN => N207);
   U1927 : OAI21_X1 port map( B1 => n1788, B2 => n1795, A => n378, ZN => N206);
   U1928 : OAI21_X1 port map( B1 => n1789, B2 => n1795, A => n378, ZN => N205);
   U1929 : OAI21_X1 port map( B1 => n1790, B2 => n1795, A => n378, ZN => N204);
   U1930 : OAI21_X1 port map( B1 => n1791, B2 => n1795, A => n378, ZN => N203);
   U1931 : NAND3_X1 port map( A1 => n1794, A2 => n1793, A3 => ADD_WR(3), ZN => 
                           n1795);
   U1932 : INV_X1 port map( A => ADD_WR(4), ZN => n1793);
   U1933 : OAI21_X1 port map( B1 => n1783, B2 => n1796, A => n378, ZN => N202);
   U1934 : OAI21_X1 port map( B1 => n1785, B2 => n1796, A => n378, ZN => N201);
   U1935 : OAI21_X1 port map( B1 => n1786, B2 => n1796, A => n378, ZN => N200);
   U1936 : OAI21_X1 port map( B1 => n1787, B2 => n1796, A => n378, ZN => N199);
   U1937 : OAI21_X1 port map( B1 => n1788, B2 => n1796, A => n378, ZN => N198);
   U1938 : OAI21_X1 port map( B1 => n1789, B2 => n1796, A => n377, ZN => N197);
   U1939 : OAI21_X1 port map( B1 => n1790, B2 => n1796, A => n377, ZN => N196);
   U1940 : OAI21_X1 port map( B1 => n1791, B2 => n1796, A => n377, ZN => N195);
   U1941 : NAND3_X1 port map( A1 => n1794, A2 => n1792, A3 => ADD_WR(4), ZN => 
                           n1796);
   U1942 : INV_X1 port map( A => ADD_WR(3), ZN => n1792);
   U1943 : OAI21_X1 port map( B1 => n1783, B2 => n1797, A => n377, ZN => N194);
   U1944 : NAND3_X1 port map( A1 => n1798, A2 => n1799, A3 => n1800, ZN => 
                           n1783);
   U1945 : OAI21_X1 port map( B1 => n1785, B2 => n1797, A => n377, ZN => N193);
   U1946 : NAND3_X1 port map( A1 => n1798, A2 => n1799, A3 => ADD_WR(0), ZN => 
                           n1785);
   U1947 : OAI21_X1 port map( B1 => n1786, B2 => n1797, A => n377, ZN => N192);
   U1948 : NAND3_X1 port map( A1 => n1800, A2 => n1799, A3 => ADD_WR(1), ZN => 
                           n1786);
   U1949 : OAI21_X1 port map( B1 => n1787, B2 => n1797, A => n377, ZN => N191);
   U1950 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1799, A3 => ADD_WR(1), ZN
                           => n1787);
   U1951 : INV_X1 port map( A => ADD_WR(2), ZN => n1799);
   U1952 : OAI21_X1 port map( B1 => n1788, B2 => n1797, A => n377, ZN => N190);
   U1953 : NAND3_X1 port map( A1 => n1800, A2 => n1798, A3 => ADD_WR(2), ZN => 
                           n1788);
   U1954 : OAI21_X1 port map( B1 => n1789, B2 => n1797, A => n377, ZN => N189);
   U1955 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1798, A3 => ADD_WR(2), ZN
                           => n1789);
   U1956 : INV_X1 port map( A => ADD_WR(1), ZN => n1798);
   U1957 : OAI21_X1 port map( B1 => n1790, B2 => n1797, A => n377, ZN => N188);
   U1958 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n1800, A3 => ADD_WR(2), ZN
                           => n1790);
   U1959 : INV_X1 port map( A => ADD_WR(0), ZN => n1800);
   U1960 : OAI21_X1 port map( B1 => n1791, B2 => n1797, A => n377, ZN => N155);
   U1961 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n1794, A3 => ADD_WR(4), ZN
                           => n1797);
   U1962 : INV_X1 port map( A => n1782, ZN => n1794);
   U1963 : NAND2_X1 port map( A1 => EN_WR, A2 => EN, ZN => n1782);
   U1964 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n1791);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity LDR_N32_6 is

   port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);  
         REGOUT : out std_logic_vector (31 downto 0));

end LDR_N32_6;

architecture SYN_STRUCTURAL of LDR_N32_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component LD_192
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_193
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_194
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_195
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_196
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_197
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_198
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_199
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_200
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_201
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_202
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_203
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_204
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_205
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_206
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_207
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_208
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_209
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_210
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_211
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_212
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_213
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_214
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_215
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_216
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_217
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_218
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_219
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_220
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_221
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_222
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LD_223
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   LDI_31 : LD_223 port map( RST => n1, EN => EN, D => REGIN(31), Q => 
                           REGOUT(31));
   LDI_30 : LD_222 port map( RST => n1, EN => EN, D => REGIN(30), Q => 
                           REGOUT(30));
   LDI_29 : LD_221 port map( RST => n1, EN => EN, D => REGIN(29), Q => 
                           REGOUT(29));
   LDI_28 : LD_220 port map( RST => n1, EN => EN, D => REGIN(28), Q => 
                           REGOUT(28));
   LDI_27 : LD_219 port map( RST => n1, EN => EN, D => REGIN(27), Q => 
                           REGOUT(27));
   LDI_26 : LD_218 port map( RST => n1, EN => EN, D => REGIN(26), Q => 
                           REGOUT(26));
   LDI_25 : LD_217 port map( RST => n1, EN => EN, D => REGIN(25), Q => 
                           REGOUT(25));
   LDI_24 : LD_216 port map( RST => n1, EN => EN, D => REGIN(24), Q => 
                           REGOUT(24));
   LDI_23 : LD_215 port map( RST => n1, EN => EN, D => REGIN(23), Q => 
                           REGOUT(23));
   LDI_22 : LD_214 port map( RST => n1, EN => EN, D => REGIN(22), Q => 
                           REGOUT(22));
   LDI_21 : LD_213 port map( RST => n1, EN => EN, D => REGIN(21), Q => 
                           REGOUT(21));
   LDI_20 : LD_212 port map( RST => n1, EN => EN, D => REGIN(20), Q => 
                           REGOUT(20));
   LDI_19 : LD_211 port map( RST => n2, EN => EN, D => REGIN(19), Q => 
                           REGOUT(19));
   LDI_18 : LD_210 port map( RST => n2, EN => EN, D => REGIN(18), Q => 
                           REGOUT(18));
   LDI_17 : LD_209 port map( RST => n2, EN => EN, D => REGIN(17), Q => 
                           REGOUT(17));
   LDI_16 : LD_208 port map( RST => n2, EN => EN, D => REGIN(16), Q => 
                           REGOUT(16));
   LDI_15 : LD_207 port map( RST => n2, EN => EN, D => REGIN(15), Q => 
                           REGOUT(15));
   LDI_14 : LD_206 port map( RST => n2, EN => EN, D => REGIN(14), Q => 
                           REGOUT(14));
   LDI_13 : LD_205 port map( RST => n2, EN => EN, D => REGIN(13), Q => 
                           REGOUT(13));
   LDI_12 : LD_204 port map( RST => n2, EN => EN, D => REGIN(12), Q => 
                           REGOUT(12));
   LDI_11 : LD_203 port map( RST => n2, EN => EN, D => REGIN(11), Q => 
                           REGOUT(11));
   LDI_10 : LD_202 port map( RST => n2, EN => EN, D => REGIN(10), Q => 
                           REGOUT(10));
   LDI_9 : LD_201 port map( RST => n2, EN => EN, D => REGIN(9), Q => REGOUT(9))
                           ;
   LDI_8 : LD_200 port map( RST => n2, EN => EN, D => REGIN(8), Q => REGOUT(8))
                           ;
   LDI_7 : LD_199 port map( RST => n3, EN => EN, D => REGIN(7), Q => REGOUT(7))
                           ;
   LDI_6 : LD_198 port map( RST => n3, EN => EN, D => REGIN(6), Q => REGOUT(6))
                           ;
   LDI_5 : LD_197 port map( RST => n3, EN => EN, D => REGIN(5), Q => REGOUT(5))
                           ;
   LDI_4 : LD_196 port map( RST => n3, EN => EN, D => REGIN(4), Q => REGOUT(4))
                           ;
   LDI_3 : LD_195 port map( RST => n3, EN => EN, D => REGIN(3), Q => REGOUT(3))
                           ;
   LDI_2 : LD_194 port map( RST => n3, EN => EN, D => REGIN(2), Q => REGOUT(2))
                           ;
   LDI_1 : LD_193 port map( RST => n3, EN => EN, D => REGIN(1), Q => REGOUT(1))
                           ;
   LDI_0 : LD_192 port map( RST => n3, EN => EN, D => REGIN(0), Q => REGOUT(0))
                           ;
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => n4, Z => n1);
   U3 : BUF_X1 port map( A => n4, Z => n2);
   U4 : BUF_X1 port map( A => n4, Z => n3);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MUX21_N32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX21_N32_4;

architecture SYN_BEHAVIORAL of MUX21_N32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(31), B => B(31), S => S, Z => Y(31));
   U2 : MUX2_X1 port map( A => A(30), B => B(30), S => S, Z => Y(30));
   U3 : MUX2_X1 port map( A => A(29), B => B(29), S => S, Z => Y(29));
   U4 : MUX2_X1 port map( A => A(28), B => B(28), S => S, Z => Y(28));
   U5 : MUX2_X1 port map( A => A(27), B => B(27), S => S, Z => Y(27));
   U6 : MUX2_X1 port map( A => A(26), B => B(26), S => S, Z => Y(26));
   U7 : MUX2_X1 port map( A => A(25), B => B(25), S => S, Z => Y(25));
   U8 : MUX2_X1 port map( A => A(24), B => B(24), S => S, Z => Y(24));
   U9 : MUX2_X1 port map( A => A(23), B => B(23), S => S, Z => Y(23));
   U10 : MUX2_X1 port map( A => A(22), B => B(22), S => S, Z => Y(22));
   U11 : MUX2_X1 port map( A => A(21), B => B(21), S => S, Z => Y(21));
   U12 : MUX2_X1 port map( A => A(20), B => B(20), S => S, Z => Y(20));
   U13 : MUX2_X1 port map( A => A(19), B => B(19), S => S, Z => Y(19));
   U14 : MUX2_X1 port map( A => A(18), B => B(18), S => S, Z => Y(18));
   U15 : MUX2_X1 port map( A => A(17), B => B(17), S => S, Z => Y(17));
   U16 : MUX2_X1 port map( A => A(16), B => B(16), S => S, Z => Y(16));
   U17 : MUX2_X1 port map( A => A(15), B => B(15), S => S, Z => Y(15));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => S, Z => Y(14));
   U19 : MUX2_X1 port map( A => A(13), B => B(13), S => S, Z => Y(13));
   U20 : MUX2_X1 port map( A => A(12), B => B(12), S => S, Z => Y(12));
   U21 : MUX2_X1 port map( A => A(11), B => B(11), S => S, Z => Y(11));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => S, Z => Y(10));
   U23 : MUX2_X1 port map( A => A(9), B => B(9), S => S, Z => Y(9));
   U24 : MUX2_X1 port map( A => A(8), B => B(8), S => S, Z => Y(8));
   U25 : MUX2_X1 port map( A => A(7), B => B(7), S => S, Z => Y(7));
   U26 : MUX2_X1 port map( A => A(6), B => B(6), S => S, Z => Y(6));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => S, Z => Y(5));
   U28 : MUX2_X1 port map( A => A(4), B => B(4), S => S, Z => Y(4));
   U29 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U30 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U31 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FFDR_N32 is

   port( CLK, RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 
         0);  REGOUT : out std_logic_vector (31 downto 0));

end FFDR_N32;

architecture SYN_STRUCTURAL of FFDR_N32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FFD_0
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_1
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_2
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_3
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_4
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_5
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_6
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_7
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_8
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_9
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_10
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_11
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_12
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_13
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_14
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_15
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_16
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_17
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_18
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_19
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_20
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_21
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_22
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_23
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_24
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_25
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_26
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_27
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_28
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_29
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_30
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FFD_31
      port( CLK, RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   FFI_31 : FFD_31 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(31), Q 
                           => REGOUT(31));
   FFI_30 : FFD_30 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(30), Q 
                           => REGOUT(30));
   FFI_29 : FFD_29 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(29), Q 
                           => REGOUT(29));
   FFI_28 : FFD_28 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(28), Q 
                           => REGOUT(28));
   FFI_27 : FFD_27 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(27), Q 
                           => REGOUT(27));
   FFI_26 : FFD_26 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(26), Q 
                           => REGOUT(26));
   FFI_25 : FFD_25 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(25), Q 
                           => REGOUT(25));
   FFI_24 : FFD_24 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(24), Q 
                           => REGOUT(24));
   FFI_23 : FFD_23 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(23), Q 
                           => REGOUT(23));
   FFI_22 : FFD_22 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(22), Q 
                           => REGOUT(22));
   FFI_21 : FFD_21 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(21), Q 
                           => REGOUT(21));
   FFI_20 : FFD_20 port map( CLK => n5, RST => n1, EN => EN, D => REGIN(20), Q 
                           => REGOUT(20));
   FFI_19 : FFD_19 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(19), Q 
                           => REGOUT(19));
   FFI_18 : FFD_18 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(18), Q 
                           => REGOUT(18));
   FFI_17 : FFD_17 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(17), Q 
                           => REGOUT(17));
   FFI_16 : FFD_16 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(16), Q 
                           => REGOUT(16));
   FFI_15 : FFD_15 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(15), Q 
                           => REGOUT(15));
   FFI_14 : FFD_14 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(14), Q 
                           => REGOUT(14));
   FFI_13 : FFD_13 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(13), Q 
                           => REGOUT(13));
   FFI_12 : FFD_12 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(12), Q 
                           => REGOUT(12));
   FFI_11 : FFD_11 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(11), Q 
                           => REGOUT(11));
   FFI_10 : FFD_10 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(10), Q 
                           => REGOUT(10));
   FFI_9 : FFD_9 port map( CLK => n6, RST => n2, EN => EN, D => REGIN(9), Q => 
                           REGOUT(9));
   FFI_8 : FFD_8 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(8), Q => 
                           REGOUT(8));
   FFI_7 : FFD_7 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(7), Q => 
                           REGOUT(7));
   FFI_6 : FFD_6 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(6), Q => 
                           REGOUT(6));
   FFI_5 : FFD_5 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(5), Q => 
                           REGOUT(5));
   FFI_4 : FFD_4 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(4), Q => 
                           REGOUT(4));
   FFI_3 : FFD_3 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(3), Q => 
                           REGOUT(3));
   FFI_2 : FFD_2 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(2), Q => 
                           REGOUT(2));
   FFI_1 : FFD_1 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(1), Q => 
                           REGOUT(1));
   FFI_0 : FFD_0 port map( CLK => n7, RST => n3, EN => EN, D => REGIN(0), Q => 
                           REGOUT(0));
   U1 : BUF_X1 port map( A => RST, Z => n4);
   U2 : BUF_X1 port map( A => CLK, Z => n8);
   U3 : BUF_X1 port map( A => n4, Z => n1);
   U4 : BUF_X1 port map( A => n4, Z => n2);
   U5 : BUF_X1 port map( A => n4, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n5);
   U7 : BUF_X1 port map( A => n8, Z => n6);
   U8 : BUF_X1 port map( A => n8, Z => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32 is

   port( CLK, RST : in std_logic;  IR_IN, DRAM_OUT : in std_logic_vector (31 
         downto 0);  IR_LATCH_EN, PC_LATCH_EN, NPC_LATCH_EN, RF_WE, 
         RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, 
         ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
         std_logic_vector (0 to 6);  LMD_LATCH_EN, JUMP_EN, JUMP_COND, 
         WB_MUX_SEL, JAL_MUX_SEL : in std_logic;  IR_OUT, PC_OUT, ALU_OUT, 
         DRAM_IN : out std_logic_vector (31 downto 0));

end DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32;

architecture SYN_DLX_DATAPATH_ARCH of 
   DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component 
      DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component MUX21_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component LDR_N32_0
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component LD_224
      port( RST, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component LDR_N32_1
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component FU_N5
      port( RS1, RS2, RD_MEM, RD_WB : in std_logic_vector (4 downto 0);  
            RF_WE_MEM, RF_WE_WB : in std_logic;  FORWARD_A, FORWARD_B : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component ZERO_DETECTOR_N32_1
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic);
   end component;
   
   component MUX21_L_320
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component ALU_N32_NB8
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  OPC : in 
            std_logic_vector (0 to 6);  Y : out std_logic_vector (31 downto 0);
            Z : out std_logic);
   end component;
   
   component MUX21_N32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_N32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX41_N32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX41_N32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component LDR_N32_2
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component LDR_N32_3
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component LDR_N32_4
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component REGADDR_N32_OPC6_REG5
      port( INSTR : in std_logic_vector (31 downto 0);  RS1, RS2, RD : out 
            std_logic_vector (4 downto 0));
   end component;
   
   component SIGNEX_N32_OPC6_REG5
      port( INSTR : in std_logic_vector (31 downto 0);  IMM : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component RF_N32_NA5
      port( RST, EN, EN_RD1, EN_RD2, EN_WR : in std_logic;  ADD_RD1, ADD_RD2, 
            ADD_WR : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component LDR_N32_5
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component LDR_N32_6
      port( RST, EN : in std_logic;  REGIN : in std_logic_vector (31 downto 0);
            REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_N32_4
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component FFDR_N32
      port( CLK, RST, EN : in std_logic;  REGIN : in std_logic_vector (31 
            downto 0);  REGOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, IR_OUT_31_port, IR_OUT_30_port, 
      IR_OUT_29_port, IR_OUT_28_port, IR_OUT_27_port, IR_OUT_26_port, 
      IR_OUT_25_port, IR_OUT_24_port, IR_OUT_23_port, IR_OUT_22_port, 
      IR_OUT_21_port, IR_OUT_20_port, IR_OUT_19_port, IR_OUT_18_port, 
      IR_OUT_17_port, IR_OUT_16_port, IR_OUT_15_port, IR_OUT_14_port, 
      IR_OUT_13_port, IR_OUT_12_port, IR_OUT_11_port, IR_OUT_10_port, 
      IR_OUT_9_port, IR_OUT_8_port, IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port
      , IR_OUT_4_port, IR_OUT_3_port, IR_OUT_2_port, IR_OUT_1_port, 
      IR_OUT_0_port, PC_OUT_31_port, PC_OUT_30_port, PC_OUT_29_port, 
      PC_OUT_28_port, PC_OUT_27_port, PC_OUT_26_port, PC_OUT_25_port, 
      PC_OUT_24_port, PC_OUT_23_port, PC_OUT_22_port, PC_OUT_21_port, 
      PC_OUT_20_port, PC_OUT_19_port, PC_OUT_18_port, PC_OUT_17_port, 
      PC_OUT_16_port, PC_OUT_15_port, PC_OUT_14_port, PC_OUT_13_port, 
      PC_OUT_12_port, PC_OUT_11_port, PC_OUT_10_port, PC_OUT_9_port, 
      PC_OUT_8_port, PC_OUT_7_port, PC_OUT_6_port, PC_OUT_5_port, PC_OUT_4_port
      , PC_OUT_3_port, PC_OUT_2_port, PC_OUT_1_port, PC_OUT_0_port, 
      ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, ALU_OUT_28_port, 
      ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, ALU_OUT_24_port, 
      ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, ALU_OUT_20_port, 
      ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, ALU_OUT_16_port, 
      ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, ALU_OUT_12_port, 
      ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, ALU_OUT_8_port, 
      ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, ALU_OUT_4_port, 
      ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, ALU_OUT_0_port, 
      IF_ID_IR_31_port, IF_ID_IR_30_port, IF_ID_IR_29_port, IF_ID_IR_28_port, 
      IF_ID_IR_27_port, IF_ID_IR_26_port, IF_ID_IR_25_port, IF_ID_IR_24_port, 
      IF_ID_IR_23_port, IF_ID_IR_22_port, IF_ID_IR_21_port, IF_ID_IR_20_port, 
      IF_ID_IR_19_port, IF_ID_IR_18_port, IF_ID_IR_17_port, IF_ID_IR_16_port, 
      IF_ID_IR_15_port, IF_ID_IR_14_port, IF_ID_IR_13_port, IF_ID_IR_12_port, 
      IF_ID_IR_11_port, IF_ID_IR_10_port, IF_ID_IR_9_port, IF_ID_IR_8_port, 
      IF_ID_IR_7_port, IF_ID_IR_6_port, IF_ID_IR_5_port, IF_ID_IR_4_port, 
      IF_ID_IR_3_port, IF_ID_IR_2_port, IF_ID_IR_1_port, IF_ID_IR_0_port, 
      ID_EX_NPC_31_port, ID_EX_NPC_30_port, ID_EX_NPC_29_port, 
      ID_EX_NPC_28_port, ID_EX_NPC_27_port, ID_EX_NPC_26_port, 
      ID_EX_NPC_25_port, ID_EX_NPC_24_port, ID_EX_NPC_23_port, 
      ID_EX_NPC_22_port, ID_EX_NPC_21_port, ID_EX_NPC_20_port, 
      ID_EX_NPC_19_port, ID_EX_NPC_18_port, ID_EX_NPC_17_port, 
      ID_EX_NPC_16_port, ID_EX_NPC_15_port, ID_EX_NPC_14_port, 
      ID_EX_NPC_13_port, ID_EX_NPC_12_port, ID_EX_NPC_11_port, 
      ID_EX_NPC_10_port, ID_EX_NPC_9_port, ID_EX_NPC_8_port, ID_EX_NPC_7_port, 
      ID_EX_NPC_6_port, ID_EX_NPC_5_port, ID_EX_NPC_4_port, ID_EX_NPC_3_port, 
      ID_EX_NPC_2_port, ID_EX_NPC_1_port, ID_EX_NPC_0_port, ID_EX_RS1_4_port, 
      ID_EX_RS1_3_port, ID_EX_RS1_2_port, ID_EX_RS1_1_port, ID_EX_RS1_0_port, 
      ID_EX_RS2_4_port, ID_EX_RS2_3_port, ID_EX_RS2_2_port, ID_EX_RS2_1_port, 
      ID_EX_RS2_0_port, ID_EX_RF_OUT1_31_port, ID_EX_RF_OUT1_30_port, 
      ID_EX_RF_OUT1_29_port, ID_EX_RF_OUT1_28_port, ID_EX_RF_OUT1_27_port, 
      ID_EX_RF_OUT1_26_port, ID_EX_RF_OUT1_25_port, ID_EX_RF_OUT1_24_port, 
      ID_EX_RF_OUT1_23_port, ID_EX_RF_OUT1_22_port, ID_EX_RF_OUT1_21_port, 
      ID_EX_RF_OUT1_20_port, ID_EX_RF_OUT1_19_port, ID_EX_RF_OUT1_18_port, 
      ID_EX_RF_OUT1_17_port, ID_EX_RF_OUT1_16_port, ID_EX_RF_OUT1_15_port, 
      ID_EX_RF_OUT1_14_port, ID_EX_RF_OUT1_13_port, ID_EX_RF_OUT1_12_port, 
      ID_EX_RF_OUT1_11_port, ID_EX_RF_OUT1_10_port, ID_EX_RF_OUT1_9_port, 
      ID_EX_RF_OUT1_8_port, ID_EX_RF_OUT1_7_port, ID_EX_RF_OUT1_6_port, 
      ID_EX_RF_OUT1_5_port, ID_EX_RF_OUT1_4_port, ID_EX_RF_OUT1_3_port, 
      ID_EX_RF_OUT1_2_port, ID_EX_RF_OUT1_1_port, ID_EX_RF_OUT1_0_port, 
      ID_EX_RF_OUT2_31_port, ID_EX_RF_OUT2_30_port, ID_EX_RF_OUT2_29_port, 
      ID_EX_RF_OUT2_28_port, ID_EX_RF_OUT2_27_port, ID_EX_RF_OUT2_26_port, 
      ID_EX_RF_OUT2_25_port, ID_EX_RF_OUT2_24_port, ID_EX_RF_OUT2_23_port, 
      ID_EX_RF_OUT2_22_port, ID_EX_RF_OUT2_21_port, ID_EX_RF_OUT2_20_port, 
      ID_EX_RF_OUT2_19_port, ID_EX_RF_OUT2_18_port, ID_EX_RF_OUT2_17_port, 
      ID_EX_RF_OUT2_16_port, ID_EX_RF_OUT2_15_port, ID_EX_RF_OUT2_14_port, 
      ID_EX_RF_OUT2_13_port, ID_EX_RF_OUT2_12_port, ID_EX_RF_OUT2_11_port, 
      ID_EX_RF_OUT2_10_port, ID_EX_RF_OUT2_9_port, ID_EX_RF_OUT2_8_port, 
      ID_EX_RF_OUT2_7_port, ID_EX_RF_OUT2_6_port, ID_EX_RF_OUT2_5_port, 
      ID_EX_RF_OUT2_4_port, ID_EX_RF_OUT2_3_port, ID_EX_RF_OUT2_2_port, 
      ID_EX_RF_OUT2_1_port, ID_EX_RF_OUT2_0_port, ID_EX_IMM_31_port, 
      ID_EX_IMM_30_port, ID_EX_IMM_29_port, ID_EX_IMM_28_port, 
      ID_EX_IMM_27_port, ID_EX_IMM_26_port, ID_EX_IMM_25_port, 
      ID_EX_IMM_24_port, ID_EX_IMM_23_port, ID_EX_IMM_22_port, 
      ID_EX_IMM_21_port, ID_EX_IMM_20_port, ID_EX_IMM_19_port, 
      ID_EX_IMM_18_port, ID_EX_IMM_17_port, ID_EX_IMM_16_port, 
      ID_EX_IMM_15_port, ID_EX_IMM_14_port, ID_EX_IMM_13_port, 
      ID_EX_IMM_12_port, ID_EX_IMM_11_port, ID_EX_IMM_10_port, ID_EX_IMM_9_port
      , ID_EX_IMM_8_port, ID_EX_IMM_7_port, ID_EX_IMM_6_port, ID_EX_IMM_5_port,
      ID_EX_IMM_4_port, ID_EX_IMM_3_port, ID_EX_IMM_2_port, ID_EX_IMM_1_port, 
      ID_EX_IMM_0_port, EX_MEM_RF_WE, EX_MEM_BRANCH_DETECT, EX_MEM_RD_4_port, 
      EX_MEM_RD_3_port, EX_MEM_RD_2_port, EX_MEM_RD_1_port, EX_MEM_RD_0_port, 
      MEM_WB_NPC_31_port, MEM_WB_NPC_30_port, MEM_WB_NPC_29_port, 
      MEM_WB_NPC_28_port, MEM_WB_NPC_27_port, MEM_WB_NPC_26_port, 
      MEM_WB_NPC_25_port, MEM_WB_NPC_24_port, MEM_WB_NPC_23_port, 
      MEM_WB_NPC_22_port, MEM_WB_NPC_21_port, MEM_WB_NPC_20_port, 
      MEM_WB_NPC_19_port, MEM_WB_NPC_18_port, MEM_WB_NPC_17_port, 
      MEM_WB_NPC_16_port, MEM_WB_NPC_15_port, MEM_WB_NPC_14_port, 
      MEM_WB_NPC_13_port, MEM_WB_NPC_12_port, MEM_WB_NPC_11_port, 
      MEM_WB_NPC_10_port, MEM_WB_NPC_9_port, MEM_WB_NPC_8_port, 
      MEM_WB_NPC_7_port, MEM_WB_NPC_6_port, MEM_WB_NPC_5_port, 
      MEM_WB_NPC_4_port, MEM_WB_NPC_3_port, MEM_WB_NPC_2_port, 
      MEM_WB_NPC_1_port, MEM_WB_NPC_0_port, MEM_WB_RF_WE, 
      MEM_WB_ALU_OUTPUT_31_port, MEM_WB_ALU_OUTPUT_30_port, 
      MEM_WB_ALU_OUTPUT_29_port, MEM_WB_ALU_OUTPUT_28_port, 
      MEM_WB_ALU_OUTPUT_27_port, MEM_WB_ALU_OUTPUT_26_port, 
      MEM_WB_ALU_OUTPUT_25_port, MEM_WB_ALU_OUTPUT_24_port, 
      MEM_WB_ALU_OUTPUT_23_port, MEM_WB_ALU_OUTPUT_22_port, 
      MEM_WB_ALU_OUTPUT_21_port, MEM_WB_ALU_OUTPUT_20_port, 
      MEM_WB_ALU_OUTPUT_19_port, MEM_WB_ALU_OUTPUT_18_port, 
      MEM_WB_ALU_OUTPUT_17_port, MEM_WB_ALU_OUTPUT_16_port, 
      MEM_WB_ALU_OUTPUT_15_port, MEM_WB_ALU_OUTPUT_14_port, 
      MEM_WB_ALU_OUTPUT_13_port, MEM_WB_ALU_OUTPUT_12_port, 
      MEM_WB_ALU_OUTPUT_11_port, MEM_WB_ALU_OUTPUT_10_port, 
      MEM_WB_ALU_OUTPUT_9_port, MEM_WB_ALU_OUTPUT_8_port, 
      MEM_WB_ALU_OUTPUT_7_port, MEM_WB_ALU_OUTPUT_6_port, 
      MEM_WB_ALU_OUTPUT_5_port, MEM_WB_ALU_OUTPUT_4_port, 
      MEM_WB_ALU_OUTPUT_3_port, MEM_WB_ALU_OUTPUT_2_port, 
      MEM_WB_ALU_OUTPUT_1_port, MEM_WB_ALU_OUTPUT_0_port, 
      MEM_WB_DRAM_OUTPUT_31_port, MEM_WB_DRAM_OUTPUT_30_port, 
      MEM_WB_DRAM_OUTPUT_29_port, MEM_WB_DRAM_OUTPUT_28_port, 
      MEM_WB_DRAM_OUTPUT_27_port, MEM_WB_DRAM_OUTPUT_26_port, 
      MEM_WB_DRAM_OUTPUT_25_port, MEM_WB_DRAM_OUTPUT_24_port, 
      MEM_WB_DRAM_OUTPUT_23_port, MEM_WB_DRAM_OUTPUT_22_port, 
      MEM_WB_DRAM_OUTPUT_21_port, MEM_WB_DRAM_OUTPUT_20_port, 
      MEM_WB_DRAM_OUTPUT_19_port, MEM_WB_DRAM_OUTPUT_18_port, 
      MEM_WB_DRAM_OUTPUT_17_port, MEM_WB_DRAM_OUTPUT_16_port, 
      MEM_WB_DRAM_OUTPUT_15_port, MEM_WB_DRAM_OUTPUT_14_port, 
      MEM_WB_DRAM_OUTPUT_13_port, MEM_WB_DRAM_OUTPUT_12_port, 
      MEM_WB_DRAM_OUTPUT_11_port, MEM_WB_DRAM_OUTPUT_10_port, 
      MEM_WB_DRAM_OUTPUT_9_port, MEM_WB_DRAM_OUTPUT_8_port, 
      MEM_WB_DRAM_OUTPUT_7_port, MEM_WB_DRAM_OUTPUT_6_port, 
      MEM_WB_DRAM_OUTPUT_5_port, MEM_WB_DRAM_OUTPUT_4_port, 
      MEM_WB_DRAM_OUTPUT_3_port, MEM_WB_DRAM_OUTPUT_2_port, 
      MEM_WB_DRAM_OUTPUT_1_port, MEM_WB_DRAM_OUTPUT_0_port, MEM_WB_RD_4_port, 
      MEM_WB_RD_3_port, MEM_WB_RD_2_port, MEM_WB_RD_1_port, MEM_WB_RD_0_port, 
      IF_ID_NPC_NEXT_31_port, IF_ID_NPC_NEXT_30_port, IF_ID_NPC_NEXT_29_port, 
      IF_ID_NPC_NEXT_28_port, IF_ID_NPC_NEXT_27_port, IF_ID_NPC_NEXT_26_port, 
      IF_ID_NPC_NEXT_25_port, IF_ID_NPC_NEXT_24_port, IF_ID_NPC_NEXT_23_port, 
      IF_ID_NPC_NEXT_22_port, IF_ID_NPC_NEXT_21_port, IF_ID_NPC_NEXT_20_port, 
      IF_ID_NPC_NEXT_19_port, IF_ID_NPC_NEXT_18_port, IF_ID_NPC_NEXT_17_port, 
      IF_ID_NPC_NEXT_16_port, IF_ID_NPC_NEXT_15_port, IF_ID_NPC_NEXT_14_port, 
      IF_ID_NPC_NEXT_13_port, IF_ID_NPC_NEXT_12_port, IF_ID_NPC_NEXT_11_port, 
      IF_ID_NPC_NEXT_10_port, IF_ID_NPC_NEXT_9_port, IF_ID_NPC_NEXT_8_port, 
      IF_ID_NPC_NEXT_7_port, IF_ID_NPC_NEXT_6_port, IF_ID_NPC_NEXT_5_port, 
      IF_ID_NPC_NEXT_4_port, IF_ID_NPC_NEXT_3_port, IF_ID_NPC_NEXT_2_port, 
      IF_ID_NPC_NEXT_1_port, IF_ID_NPC_NEXT_0_port, ID_EX_RS1_NEXT_4_port, 
      ID_EX_RS1_NEXT_3_port, ID_EX_RS1_NEXT_2_port, ID_EX_RS1_NEXT_1_port, 
      ID_EX_RS1_NEXT_0_port, ID_EX_RS2_NEXT_4_port, ID_EX_RS2_NEXT_3_port, 
      ID_EX_RS2_NEXT_2_port, ID_EX_RS2_NEXT_1_port, ID_EX_RS2_NEXT_0_port, 
      ID_EX_RD_NEXT_4_port, ID_EX_RD_NEXT_3_port, ID_EX_RD_NEXT_2_port, 
      ID_EX_RD_NEXT_1_port, ID_EX_RD_NEXT_0_port, ID_EX_RF_OUT1_NEXT_31_port, 
      ID_EX_RF_OUT1_NEXT_30_port, ID_EX_RF_OUT1_NEXT_29_port, 
      ID_EX_RF_OUT1_NEXT_28_port, ID_EX_RF_OUT1_NEXT_27_port, 
      ID_EX_RF_OUT1_NEXT_26_port, ID_EX_RF_OUT1_NEXT_25_port, 
      ID_EX_RF_OUT1_NEXT_24_port, ID_EX_RF_OUT1_NEXT_23_port, 
      ID_EX_RF_OUT1_NEXT_22_port, ID_EX_RF_OUT1_NEXT_21_port, 
      ID_EX_RF_OUT1_NEXT_20_port, ID_EX_RF_OUT1_NEXT_19_port, 
      ID_EX_RF_OUT1_NEXT_18_port, ID_EX_RF_OUT1_NEXT_17_port, 
      ID_EX_RF_OUT1_NEXT_16_port, ID_EX_RF_OUT1_NEXT_15_port, 
      ID_EX_RF_OUT1_NEXT_14_port, ID_EX_RF_OUT1_NEXT_13_port, 
      ID_EX_RF_OUT1_NEXT_12_port, ID_EX_RF_OUT1_NEXT_11_port, 
      ID_EX_RF_OUT1_NEXT_10_port, ID_EX_RF_OUT1_NEXT_9_port, 
      ID_EX_RF_OUT1_NEXT_8_port, ID_EX_RF_OUT1_NEXT_7_port, 
      ID_EX_RF_OUT1_NEXT_6_port, ID_EX_RF_OUT1_NEXT_5_port, 
      ID_EX_RF_OUT1_NEXT_4_port, ID_EX_RF_OUT1_NEXT_3_port, 
      ID_EX_RF_OUT1_NEXT_2_port, ID_EX_RF_OUT1_NEXT_1_port, 
      ID_EX_RF_OUT1_NEXT_0_port, ID_EX_RF_OUT2_NEXT_31_port, 
      ID_EX_RF_OUT2_NEXT_30_port, ID_EX_RF_OUT2_NEXT_29_port, 
      ID_EX_RF_OUT2_NEXT_28_port, ID_EX_RF_OUT2_NEXT_27_port, 
      ID_EX_RF_OUT2_NEXT_26_port, ID_EX_RF_OUT2_NEXT_25_port, 
      ID_EX_RF_OUT2_NEXT_24_port, ID_EX_RF_OUT2_NEXT_23_port, 
      ID_EX_RF_OUT2_NEXT_22_port, ID_EX_RF_OUT2_NEXT_21_port, 
      ID_EX_RF_OUT2_NEXT_20_port, ID_EX_RF_OUT2_NEXT_19_port, 
      ID_EX_RF_OUT2_NEXT_18_port, ID_EX_RF_OUT2_NEXT_17_port, 
      ID_EX_RF_OUT2_NEXT_16_port, ID_EX_RF_OUT2_NEXT_15_port, 
      ID_EX_RF_OUT2_NEXT_14_port, ID_EX_RF_OUT2_NEXT_13_port, 
      ID_EX_RF_OUT2_NEXT_12_port, ID_EX_RF_OUT2_NEXT_11_port, 
      ID_EX_RF_OUT2_NEXT_10_port, ID_EX_RF_OUT2_NEXT_9_port, 
      ID_EX_RF_OUT2_NEXT_8_port, ID_EX_RF_OUT2_NEXT_7_port, 
      ID_EX_RF_OUT2_NEXT_6_port, ID_EX_RF_OUT2_NEXT_5_port, 
      ID_EX_RF_OUT2_NEXT_4_port, ID_EX_RF_OUT2_NEXT_3_port, 
      ID_EX_RF_OUT2_NEXT_2_port, ID_EX_RF_OUT2_NEXT_1_port, 
      ID_EX_RF_OUT2_NEXT_0_port, ID_EX_IMM_NEXT_31_port, ID_EX_IMM_NEXT_30_port
      , ID_EX_IMM_NEXT_29_port, ID_EX_IMM_NEXT_28_port, ID_EX_IMM_NEXT_27_port,
      ID_EX_IMM_NEXT_26_port, ID_EX_IMM_NEXT_25_port, ID_EX_IMM_NEXT_24_port, 
      ID_EX_IMM_NEXT_23_port, ID_EX_IMM_NEXT_22_port, ID_EX_IMM_NEXT_21_port, 
      ID_EX_IMM_NEXT_20_port, ID_EX_IMM_NEXT_19_port, ID_EX_IMM_NEXT_18_port, 
      ID_EX_IMM_NEXT_17_port, ID_EX_IMM_NEXT_16_port, ID_EX_IMM_NEXT_15_port, 
      ID_EX_IMM_NEXT_14_port, ID_EX_IMM_NEXT_13_port, ID_EX_IMM_NEXT_12_port, 
      ID_EX_IMM_NEXT_11_port, ID_EX_IMM_NEXT_10_port, ID_EX_IMM_NEXT_9_port, 
      ID_EX_IMM_NEXT_8_port, ID_EX_IMM_NEXT_7_port, ID_EX_IMM_NEXT_6_port, 
      ID_EX_IMM_NEXT_5_port, ID_EX_IMM_NEXT_4_port, ID_EX_IMM_NEXT_3_port, 
      ID_EX_IMM_NEXT_2_port, ID_EX_IMM_NEXT_1_port, ID_EX_IMM_NEXT_0_port, 
      EX_MEM_ALU_OUTPUT_NEXT_31_port, EX_MEM_ALU_OUTPUT_NEXT_30_port, 
      EX_MEM_ALU_OUTPUT_NEXT_29_port, EX_MEM_ALU_OUTPUT_NEXT_28_port, 
      EX_MEM_ALU_OUTPUT_NEXT_27_port, EX_MEM_ALU_OUTPUT_NEXT_26_port, 
      EX_MEM_ALU_OUTPUT_NEXT_25_port, EX_MEM_ALU_OUTPUT_NEXT_24_port, 
      EX_MEM_ALU_OUTPUT_NEXT_23_port, EX_MEM_ALU_OUTPUT_NEXT_22_port, 
      EX_MEM_ALU_OUTPUT_NEXT_21_port, EX_MEM_ALU_OUTPUT_NEXT_20_port, 
      EX_MEM_ALU_OUTPUT_NEXT_19_port, EX_MEM_ALU_OUTPUT_NEXT_18_port, 
      EX_MEM_ALU_OUTPUT_NEXT_17_port, EX_MEM_ALU_OUTPUT_NEXT_16_port, 
      EX_MEM_ALU_OUTPUT_NEXT_15_port, EX_MEM_ALU_OUTPUT_NEXT_14_port, 
      EX_MEM_ALU_OUTPUT_NEXT_13_port, EX_MEM_ALU_OUTPUT_NEXT_12_port, 
      EX_MEM_ALU_OUTPUT_NEXT_11_port, EX_MEM_ALU_OUTPUT_NEXT_10_port, 
      EX_MEM_ALU_OUTPUT_NEXT_9_port, EX_MEM_ALU_OUTPUT_NEXT_8_port, 
      EX_MEM_ALU_OUTPUT_NEXT_7_port, EX_MEM_ALU_OUTPUT_NEXT_6_port, 
      EX_MEM_ALU_OUTPUT_NEXT_5_port, EX_MEM_ALU_OUTPUT_NEXT_4_port, 
      EX_MEM_ALU_OUTPUT_NEXT_3_port, EX_MEM_ALU_OUTPUT_NEXT_2_port, 
      EX_MEM_ALU_OUTPUT_NEXT_1_port, EX_MEM_ALU_OUTPUT_NEXT_0_port, 
      EX_MEM_BRANCH_DETECT_NEXT, MEM_WB_DRAM_OUTPUT_NEXT_31_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_30_port, MEM_WB_DRAM_OUTPUT_NEXT_29_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_28_port, MEM_WB_DRAM_OUTPUT_NEXT_27_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_26_port, MEM_WB_DRAM_OUTPUT_NEXT_25_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_24_port, MEM_WB_DRAM_OUTPUT_NEXT_23_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_22_port, MEM_WB_DRAM_OUTPUT_NEXT_21_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_20_port, MEM_WB_DRAM_OUTPUT_NEXT_19_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_18_port, MEM_WB_DRAM_OUTPUT_NEXT_17_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_16_port, MEM_WB_DRAM_OUTPUT_NEXT_15_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_14_port, MEM_WB_DRAM_OUTPUT_NEXT_13_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_12_port, MEM_WB_DRAM_OUTPUT_NEXT_11_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_10_port, MEM_WB_DRAM_OUTPUT_NEXT_9_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_8_port, MEM_WB_DRAM_OUTPUT_NEXT_7_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_6_port, MEM_WB_DRAM_OUTPUT_NEXT_5_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_4_port, MEM_WB_DRAM_OUTPUT_NEXT_3_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_2_port, MEM_WB_DRAM_OUTPUT_NEXT_1_port, 
      MEM_WB_DRAM_OUTPUT_NEXT_0_port, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11,
      N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26
      , N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, 
      N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55
      , N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, 
      N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84
      , N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, 
      N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, 
      N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, 
      N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, 
      N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, 
      N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, 
      N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, 
      N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, 
      N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, 
      N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, 
      N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, 
      N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, 
      N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, 
      N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, 
      N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, 
      N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, 
      N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, 
      N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, 
      N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, 
      N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, 
      N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, 
      N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, 
      N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, 
      N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, 
      N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, 
      N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, 
      N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, 
      N411, N412, N413, N414, NPC_BUS_31_port, NPC_BUS_30_port, NPC_BUS_29_port
      , NPC_BUS_28_port, NPC_BUS_27_port, NPC_BUS_26_port, NPC_BUS_25_port, 
      NPC_BUS_24_port, NPC_BUS_23_port, NPC_BUS_22_port, NPC_BUS_21_port, 
      NPC_BUS_20_port, NPC_BUS_19_port, NPC_BUS_18_port, NPC_BUS_17_port, 
      NPC_BUS_16_port, NPC_BUS_15_port, NPC_BUS_14_port, NPC_BUS_13_port, 
      NPC_BUS_12_port, NPC_BUS_11_port, NPC_BUS_10_port, NPC_BUS_9_port, 
      NPC_BUS_8_port, NPC_BUS_7_port, NPC_BUS_6_port, NPC_BUS_5_port, 
      NPC_BUS_4_port, NPC_BUS_3_port, NPC_BUS_2_port, NPC_BUS_1_port, 
      NPC_BUS_0_port, ZERO_OUT, PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port,
      PC_BUS_28_port, PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, 
      PC_BUS_24_port, PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, 
      PC_BUS_20_port, PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, 
      PC_BUS_16_port, PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, 
      PC_BUS_12_port, PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, 
      PC_BUS_8_port, PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port
      , PC_BUS_3_port, PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, 
      JAL_MUX_OUT_31_port, JAL_MUX_OUT_30_port, JAL_MUX_OUT_29_port, 
      JAL_MUX_OUT_28_port, JAL_MUX_OUT_27_port, JAL_MUX_OUT_26_port, 
      JAL_MUX_OUT_25_port, JAL_MUX_OUT_24_port, JAL_MUX_OUT_23_port, 
      JAL_MUX_OUT_22_port, JAL_MUX_OUT_21_port, JAL_MUX_OUT_20_port, 
      JAL_MUX_OUT_19_port, JAL_MUX_OUT_18_port, JAL_MUX_OUT_17_port, 
      JAL_MUX_OUT_16_port, JAL_MUX_OUT_15_port, JAL_MUX_OUT_14_port, 
      JAL_MUX_OUT_13_port, JAL_MUX_OUT_12_port, JAL_MUX_OUT_11_port, 
      JAL_MUX_OUT_10_port, JAL_MUX_OUT_9_port, JAL_MUX_OUT_8_port, 
      JAL_MUX_OUT_7_port, JAL_MUX_OUT_6_port, JAL_MUX_OUT_5_port, 
      JAL_MUX_OUT_4_port, JAL_MUX_OUT_3_port, JAL_MUX_OUT_2_port, 
      JAL_MUX_OUT_1_port, JAL_MUX_OUT_0_port, RF_OUT1_31_port, RF_OUT1_30_port,
      RF_OUT1_29_port, RF_OUT1_28_port, RF_OUT1_27_port, RF_OUT1_26_port, 
      RF_OUT1_25_port, RF_OUT1_24_port, RF_OUT1_23_port, RF_OUT1_22_port, 
      RF_OUT1_21_port, RF_OUT1_20_port, RF_OUT1_19_port, RF_OUT1_18_port, 
      RF_OUT1_17_port, RF_OUT1_16_port, RF_OUT1_15_port, RF_OUT1_14_port, 
      RF_OUT1_13_port, RF_OUT1_12_port, RF_OUT1_11_port, RF_OUT1_10_port, 
      RF_OUT1_9_port, RF_OUT1_8_port, RF_OUT1_7_port, RF_OUT1_6_port, 
      RF_OUT1_5_port, RF_OUT1_4_port, RF_OUT1_3_port, RF_OUT1_2_port, 
      RF_OUT1_1_port, RF_OUT1_0_port, RF_OUT2_31_port, RF_OUT2_30_port, 
      RF_OUT2_29_port, RF_OUT2_28_port, RF_OUT2_27_port, RF_OUT2_26_port, 
      RF_OUT2_25_port, RF_OUT2_24_port, RF_OUT2_23_port, RF_OUT2_22_port, 
      RF_OUT2_21_port, RF_OUT2_20_port, RF_OUT2_19_port, RF_OUT2_18_port, 
      RF_OUT2_17_port, RF_OUT2_16_port, RF_OUT2_15_port, RF_OUT2_14_port, 
      RF_OUT2_13_port, RF_OUT2_12_port, RF_OUT2_11_port, RF_OUT2_10_port, 
      RF_OUT2_9_port, RF_OUT2_8_port, RF_OUT2_7_port, RF_OUT2_6_port, 
      RF_OUT2_5_port, RF_OUT2_4_port, RF_OUT2_3_port, RF_OUT2_2_port, 
      RF_OUT2_1_port, RF_OUT2_0_port, IMM_OUT_31_port, IMM_OUT_30_port, 
      IMM_OUT_29_port, IMM_OUT_28_port, IMM_OUT_27_port, IMM_OUT_26_port, 
      IMM_OUT_25_port, IMM_OUT_24_port, IMM_OUT_23_port, IMM_OUT_22_port, 
      IMM_OUT_21_port, IMM_OUT_20_port, IMM_OUT_19_port, IMM_OUT_18_port, 
      IMM_OUT_17_port, IMM_OUT_16_port, IMM_OUT_15_port, IMM_OUT_14_port, 
      IMM_OUT_13_port, IMM_OUT_12_port, IMM_OUT_11_port, IMM_OUT_10_port, 
      IMM_OUT_9_port, IMM_OUT_8_port, IMM_OUT_7_port, IMM_OUT_6_port, 
      IMM_OUT_5_port, IMM_OUT_4_port, IMM_OUT_3_port, IMM_OUT_2_port, 
      IMM_OUT_1_port, IMM_OUT_0_port, FORWARD_A_1_port, FORWARD_A_0_port, 
      ALU_PREOP1_31_port, ALU_PREOP1_30_port, ALU_PREOP1_29_port, 
      ALU_PREOP1_28_port, ALU_PREOP1_27_port, ALU_PREOP1_26_port, 
      ALU_PREOP1_25_port, ALU_PREOP1_24_port, ALU_PREOP1_23_port, 
      ALU_PREOP1_22_port, ALU_PREOP1_21_port, ALU_PREOP1_20_port, 
      ALU_PREOP1_19_port, ALU_PREOP1_18_port, ALU_PREOP1_17_port, 
      ALU_PREOP1_16_port, ALU_PREOP1_15_port, ALU_PREOP1_14_port, 
      ALU_PREOP1_13_port, ALU_PREOP1_12_port, ALU_PREOP1_11_port, 
      ALU_PREOP1_10_port, ALU_PREOP1_9_port, ALU_PREOP1_8_port, 
      ALU_PREOP1_7_port, ALU_PREOP1_6_port, ALU_PREOP1_5_port, 
      ALU_PREOP1_4_port, ALU_PREOP1_3_port, ALU_PREOP1_2_port, 
      ALU_PREOP1_1_port, ALU_PREOP1_0_port, FORWARD_B_1_port, FORWARD_B_0_port,
      ALU_PREOP2_31_port, ALU_PREOP2_30_port, ALU_PREOP2_29_port, 
      ALU_PREOP2_28_port, ALU_PREOP2_27_port, ALU_PREOP2_26_port, 
      ALU_PREOP2_25_port, ALU_PREOP2_24_port, ALU_PREOP2_23_port, 
      ALU_PREOP2_22_port, ALU_PREOP2_21_port, ALU_PREOP2_20_port, 
      ALU_PREOP2_19_port, ALU_PREOP2_18_port, ALU_PREOP2_17_port, 
      ALU_PREOP2_16_port, ALU_PREOP2_15_port, ALU_PREOP2_14_port, 
      ALU_PREOP2_13_port, ALU_PREOP2_12_port, ALU_PREOP2_11_port, 
      ALU_PREOP2_10_port, ALU_PREOP2_9_port, ALU_PREOP2_8_port, 
      ALU_PREOP2_7_port, ALU_PREOP2_6_port, ALU_PREOP2_5_port, 
      ALU_PREOP2_4_port, ALU_PREOP2_3_port, ALU_PREOP2_2_port, 
      ALU_PREOP2_1_port, ALU_PREOP2_0_port, ALU_OP1_31_port, ALU_OP1_30_port, 
      ALU_OP1_29_port, ALU_OP1_28_port, ALU_OP1_27_port, ALU_OP1_26_port, 
      ALU_OP1_25_port, ALU_OP1_24_port, ALU_OP1_23_port, ALU_OP1_22_port, 
      ALU_OP1_21_port, ALU_OP1_20_port, ALU_OP1_19_port, ALU_OP1_18_port, 
      ALU_OP1_17_port, ALU_OP1_16_port, ALU_OP1_15_port, ALU_OP1_14_port, 
      ALU_OP1_13_port, ALU_OP1_12_port, ALU_OP1_11_port, ALU_OP1_10_port, 
      ALU_OP1_9_port, ALU_OP1_8_port, ALU_OP1_7_port, ALU_OP1_6_port, 
      ALU_OP1_5_port, ALU_OP1_4_port, ALU_OP1_3_port, ALU_OP1_2_port, 
      ALU_OP1_1_port, ALU_OP1_0_port, ALU_OP2_31_port, ALU_OP2_30_port, 
      ALU_OP2_29_port, ALU_OP2_28_port, ALU_OP2_27_port, ALU_OP2_26_port, 
      ALU_OP2_25_port, ALU_OP2_24_port, ALU_OP2_23_port, ALU_OP2_22_port, 
      ALU_OP2_21_port, ALU_OP2_20_port, ALU_OP2_19_port, ALU_OP2_18_port, 
      ALU_OP2_17_port, ALU_OP2_16_port, ALU_OP2_15_port, ALU_OP2_14_port, 
      ALU_OP2_13_port, ALU_OP2_12_port, ALU_OP2_11_port, ALU_OP2_10_port, 
      ALU_OP2_9_port, ALU_OP2_8_port, ALU_OP2_7_port, ALU_OP2_6_port, 
      ALU_OP2_5_port, ALU_OP2_4_port, ALU_OP2_3_port, ALU_OP2_2_port, 
      ALU_OP2_1_port, ALU_OP2_0_port, ALU_OUTPUT_31_port, ALU_OUTPUT_30_port, 
      ALU_OUTPUT_29_port, ALU_OUTPUT_28_port, ALU_OUTPUT_27_port, 
      ALU_OUTPUT_26_port, ALU_OUTPUT_25_port, ALU_OUTPUT_24_port, 
      ALU_OUTPUT_23_port, ALU_OUTPUT_22_port, ALU_OUTPUT_21_port, 
      ALU_OUTPUT_20_port, ALU_OUTPUT_19_port, ALU_OUTPUT_18_port, 
      ALU_OUTPUT_17_port, ALU_OUTPUT_16_port, ALU_OUTPUT_15_port, 
      ALU_OUTPUT_14_port, ALU_OUTPUT_13_port, ALU_OUTPUT_12_port, 
      ALU_OUTPUT_11_port, ALU_OUTPUT_10_port, ALU_OUTPUT_9_port, 
      ALU_OUTPUT_8_port, ALU_OUTPUT_7_port, ALU_OUTPUT_6_port, 
      ALU_OUTPUT_5_port, ALU_OUTPUT_4_port, ALU_OUTPUT_3_port, 
      ALU_OUTPUT_2_port, ALU_OUTPUT_1_port, ALU_OUTPUT_0_port, BRANCH_DETECT, 
      WB_MUX_OUT_31_port, WB_MUX_OUT_30_port, WB_MUX_OUT_29_port, 
      WB_MUX_OUT_28_port, WB_MUX_OUT_27_port, WB_MUX_OUT_26_port, 
      WB_MUX_OUT_25_port, WB_MUX_OUT_24_port, WB_MUX_OUT_23_port, 
      WB_MUX_OUT_22_port, WB_MUX_OUT_21_port, WB_MUX_OUT_20_port, 
      WB_MUX_OUT_19_port, WB_MUX_OUT_18_port, WB_MUX_OUT_17_port, 
      WB_MUX_OUT_16_port, WB_MUX_OUT_15_port, WB_MUX_OUT_14_port, 
      WB_MUX_OUT_13_port, WB_MUX_OUT_12_port, WB_MUX_OUT_11_port, 
      WB_MUX_OUT_10_port, WB_MUX_OUT_9_port, WB_MUX_OUT_8_port, 
      WB_MUX_OUT_7_port, WB_MUX_OUT_6_port, WB_MUX_OUT_5_port, 
      WB_MUX_OUT_4_port, WB_MUX_OUT_3_port, WB_MUX_OUT_2_port, 
      WB_MUX_OUT_1_port, WB_MUX_OUT_0_port, n1, n2_port, n3_port, n4_port, 
      n5_port, n6_port, n7_port, n8_port, n9_port, n10_port, n11_port, n12_port
      , n13_port, n14_port, n15_port, n16_port, n17_port, n18_port, n19_port, 
      n20_port, n21_port, n22_port, n23_port, n24_port, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, 
      n62_port, n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, 
      n69_port, n70_port, n71_port, n72_port, n73_port, n74_port, n75_port, 
      n76_port, n77_port, n78_port, n79_port, n80_port, n81_port, n82_port, 
      n83_port, n84_port, n85_port, n86_port, n87_port, n88_port, n89_port, 
      n90_port, n91_port, n92_port, n93_port, n94_port, n95_port, n96_port, 
      n97_port, n98_port, n99_port, n100_port, n101_port, n102_port, n103_port,
      n104_port, n105_port, n106_port, n107_port, n108_port, n109_port, 
      n110_port, n111_port, n112_port, n113_port, n114_port, n115_port, 
      n116_port, n117_port, n118_port, n119_port, n120_port, n121_port, 
      n122_port, n123_port, n124_port, n125_port, n126_port, n127_port, 
      n128_port, n129_port, n130_port, n131_port, n132_port, n133_port, 
      n134_port, n135_port, n136_port, n137_port, n138_port, n139_port, 
      n140_port, n141_port, n142_port, n143_port, n144_port, n145_port, 
      n146_port, n147_port, n148_port, n149_port, n150_port, n151_port, 
      n152_port, n153_port, n154_port, n155_port, n156_port, n157_port, 
      n158_port, n159_port, n160_port, n161_port, n162_port, n163_port, 
      n164_port, n165_port, n166_port, n167_port, n168_port, n169_port, 
      n170_port, n171_port, n172_port, n173_port, n174_port, n175_port, 
      n176_port, n177_port, n178_port, n179_port, n180_port, n181_port, 
      n182_port, n183_port, n184_port, n185_port, n186_port, n187_port, n_1316,
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628 : std_logic;

begin
   IR_OUT <= ( IR_OUT_31_port, IR_OUT_30_port, IR_OUT_29_port, IR_OUT_28_port, 
      IR_OUT_27_port, IR_OUT_26_port, IR_OUT_25_port, IR_OUT_24_port, 
      IR_OUT_23_port, IR_OUT_22_port, IR_OUT_21_port, IR_OUT_20_port, 
      IR_OUT_19_port, IR_OUT_18_port, IR_OUT_17_port, IR_OUT_16_port, 
      IR_OUT_15_port, IR_OUT_14_port, IR_OUT_13_port, IR_OUT_12_port, 
      IR_OUT_11_port, IR_OUT_10_port, IR_OUT_9_port, IR_OUT_8_port, 
      IR_OUT_7_port, IR_OUT_6_port, IR_OUT_5_port, IR_OUT_4_port, IR_OUT_3_port
      , IR_OUT_2_port, IR_OUT_1_port, IR_OUT_0_port );
   PC_OUT <= ( PC_OUT_31_port, PC_OUT_30_port, PC_OUT_29_port, PC_OUT_28_port, 
      PC_OUT_27_port, PC_OUT_26_port, PC_OUT_25_port, PC_OUT_24_port, 
      PC_OUT_23_port, PC_OUT_22_port, PC_OUT_21_port, PC_OUT_20_port, 
      PC_OUT_19_port, PC_OUT_18_port, PC_OUT_17_port, PC_OUT_16_port, 
      PC_OUT_15_port, PC_OUT_14_port, PC_OUT_13_port, PC_OUT_12_port, 
      PC_OUT_11_port, PC_OUT_10_port, PC_OUT_9_port, PC_OUT_8_port, 
      PC_OUT_7_port, PC_OUT_6_port, PC_OUT_5_port, PC_OUT_4_port, PC_OUT_3_port
      , PC_OUT_2_port, PC_OUT_1_port, PC_OUT_0_port );
   ALU_OUT <= ( ALU_OUT_31_port, ALU_OUT_30_port, ALU_OUT_29_port, 
      ALU_OUT_28_port, ALU_OUT_27_port, ALU_OUT_26_port, ALU_OUT_25_port, 
      ALU_OUT_24_port, ALU_OUT_23_port, ALU_OUT_22_port, ALU_OUT_21_port, 
      ALU_OUT_20_port, ALU_OUT_19_port, ALU_OUT_18_port, ALU_OUT_17_port, 
      ALU_OUT_16_port, ALU_OUT_15_port, ALU_OUT_14_port, ALU_OUT_13_port, 
      ALU_OUT_12_port, ALU_OUT_11_port, ALU_OUT_10_port, ALU_OUT_9_port, 
      ALU_OUT_8_port, ALU_OUT_7_port, ALU_OUT_6_port, ALU_OUT_5_port, 
      ALU_OUT_4_port, ALU_OUT_3_port, ALU_OUT_2_port, ALU_OUT_1_port, 
      ALU_OUT_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n1 <= '0';
   IF_ID_IR_reg_31_inst : DFF_X1 port map( D => N65, CK => n10_port, Q => 
                           IF_ID_IR_31_port, QN => n_1316);
   IF_ID_IR_reg_30_inst : DFF_X1 port map( D => N64, CK => n10_port, Q => 
                           IF_ID_IR_30_port, QN => n_1317);
   IF_ID_IR_reg_29_inst : DFF_X1 port map( D => N63, CK => n10_port, Q => 
                           IF_ID_IR_29_port, QN => n_1318);
   IF_ID_IR_reg_28_inst : DFF_X1 port map( D => N62, CK => n10_port, Q => 
                           IF_ID_IR_28_port, QN => n_1319);
   IF_ID_IR_reg_27_inst : DFF_X1 port map( D => N61, CK => n10_port, Q => 
                           IF_ID_IR_27_port, QN => n_1320);
   IF_ID_IR_reg_26_inst : DFF_X1 port map( D => N60, CK => n10_port, Q => 
                           IF_ID_IR_26_port, QN => n_1321);
   IF_ID_IR_reg_25_inst : DFF_X1 port map( D => N59, CK => n10_port, Q => 
                           IF_ID_IR_25_port, QN => n_1322);
   IF_ID_IR_reg_24_inst : DFF_X1 port map( D => N58, CK => n10_port, Q => 
                           IF_ID_IR_24_port, QN => n_1323);
   IF_ID_IR_reg_23_inst : DFF_X1 port map( D => N57, CK => n10_port, Q => 
                           IF_ID_IR_23_port, QN => n_1324);
   IF_ID_IR_reg_22_inst : DFF_X1 port map( D => N56, CK => n10_port, Q => 
                           IF_ID_IR_22_port, QN => n_1325);
   IF_ID_IR_reg_21_inst : DFF_X1 port map( D => N55, CK => n10_port, Q => 
                           IF_ID_IR_21_port, QN => n_1326);
   IF_ID_IR_reg_20_inst : DFF_X1 port map( D => N54, CK => n10_port, Q => 
                           IF_ID_IR_20_port, QN => n_1327);
   IF_ID_IR_reg_19_inst : DFF_X1 port map( D => N53, CK => n10_port, Q => 
                           IF_ID_IR_19_port, QN => n_1328);
   IF_ID_IR_reg_18_inst : DFF_X1 port map( D => N52, CK => n10_port, Q => 
                           IF_ID_IR_18_port, QN => n_1329);
   IF_ID_IR_reg_17_inst : DFF_X1 port map( D => N51, CK => n10_port, Q => 
                           IF_ID_IR_17_port, QN => n_1330);
   IF_ID_IR_reg_16_inst : DFF_X1 port map( D => N50, CK => n10_port, Q => 
                           IF_ID_IR_16_port, QN => n_1331);
   IF_ID_IR_reg_15_inst : DFF_X1 port map( D => N49, CK => n10_port, Q => 
                           IF_ID_IR_15_port, QN => n_1332);
   IF_ID_IR_reg_14_inst : DFF_X1 port map( D => N48, CK => n10_port, Q => 
                           IF_ID_IR_14_port, QN => n_1333);
   IF_ID_IR_reg_13_inst : DFF_X1 port map( D => N47, CK => n10_port, Q => 
                           IF_ID_IR_13_port, QN => n_1334);
   IF_ID_IR_reg_12_inst : DFF_X1 port map( D => N46, CK => n10_port, Q => 
                           IF_ID_IR_12_port, QN => n_1335);
   IF_ID_IR_reg_11_inst : DFF_X1 port map( D => N45, CK => n10_port, Q => 
                           IF_ID_IR_11_port, QN => n_1336);
   IF_ID_IR_reg_10_inst : DFF_X1 port map( D => N44, CK => n10_port, Q => 
                           IF_ID_IR_10_port, QN => n_1337);
   IF_ID_IR_reg_9_inst : DFF_X1 port map( D => N43, CK => n10_port, Q => 
                           IF_ID_IR_9_port, QN => n_1338);
   IF_ID_IR_reg_8_inst : DFF_X1 port map( D => N42, CK => n10_port, Q => 
                           IF_ID_IR_8_port, QN => n_1339);
   IF_ID_IR_reg_7_inst : DFF_X1 port map( D => N41, CK => n10_port, Q => 
                           IF_ID_IR_7_port, QN => n_1340);
   IF_ID_IR_reg_6_inst : DFF_X1 port map( D => N40, CK => n10_port, Q => 
                           IF_ID_IR_6_port, QN => n_1341);
   IF_ID_IR_reg_5_inst : DFF_X1 port map( D => N39, CK => n10_port, Q => 
                           IF_ID_IR_5_port, QN => n_1342);
   IF_ID_IR_reg_4_inst : DFF_X1 port map( D => N38, CK => n10_port, Q => 
                           IF_ID_IR_4_port, QN => n_1343);
   IF_ID_IR_reg_3_inst : DFF_X1 port map( D => N37, CK => n10_port, Q => 
                           IF_ID_IR_3_port, QN => n_1344);
   IF_ID_IR_reg_2_inst : DFF_X1 port map( D => N36, CK => n10_port, Q => 
                           IF_ID_IR_2_port, QN => n_1345);
   IF_ID_IR_reg_1_inst : DFF_X1 port map( D => N35, CK => n10_port, Q => 
                           IF_ID_IR_1_port, QN => n_1346);
   IF_ID_IR_reg_0_inst : DFF_X1 port map( D => N34, CK => n10_port, Q => 
                           IF_ID_IR_0_port, QN => n_1347);
   ID_EX_RF_WE_reg : DFF_X1 port map( D => N98, CK => n11_port, Q => n_1348, QN
                           => n153_port);
   ID_EX_RS1_reg_4_inst : DFF_X1 port map( D => N103, CK => n10_port, Q => 
                           ID_EX_RS1_4_port, QN => n_1349);
   ID_EX_RS1_reg_3_inst : DFF_X1 port map( D => N102, CK => n10_port, Q => 
                           ID_EX_RS1_3_port, QN => n_1350);
   ID_EX_RS1_reg_2_inst : DFF_X1 port map( D => N101, CK => n10_port, Q => 
                           ID_EX_RS1_2_port, QN => n_1351);
   ID_EX_RS1_reg_1_inst : DFF_X1 port map( D => N100, CK => n10_port, Q => 
                           ID_EX_RS1_1_port, QN => n_1352);
   ID_EX_RS1_reg_0_inst : DFF_X1 port map( D => N99, CK => n10_port, Q => 
                           ID_EX_RS1_0_port, QN => n_1353);
   ID_EX_RS2_reg_4_inst : DFF_X1 port map( D => N108, CK => n10_port, Q => 
                           ID_EX_RS2_4_port, QN => n_1354);
   ID_EX_RS2_reg_3_inst : DFF_X1 port map( D => N107, CK => n10_port, Q => 
                           ID_EX_RS2_3_port, QN => n_1355);
   ID_EX_RS2_reg_2_inst : DFF_X1 port map( D => N106, CK => n10_port, Q => 
                           ID_EX_RS2_2_port, QN => n_1356);
   ID_EX_RS2_reg_1_inst : DFF_X1 port map( D => N105, CK => n10_port, Q => 
                           ID_EX_RS2_1_port, QN => n_1357);
   ID_EX_RS2_reg_0_inst : DFF_X1 port map( D => N104, CK => n10_port, Q => 
                           ID_EX_RS2_0_port, QN => n_1358);
   ID_EX_RD_reg_4_inst : DFF_X1 port map( D => N113, CK => n10_port, Q => 
                           n_1359, QN => n116_port);
   ID_EX_RD_reg_3_inst : DFF_X1 port map( D => N112, CK => n10_port, Q => 
                           n_1360, QN => n117_port);
   ID_EX_RD_reg_2_inst : DFF_X1 port map( D => N111, CK => n10_port, Q => 
                           n_1361, QN => n118_port);
   ID_EX_RD_reg_1_inst : DFF_X1 port map( D => N110, CK => n10_port, Q => 
                           n_1362, QN => n119_port);
   ID_EX_RD_reg_0_inst : DFF_X1 port map( D => N109, CK => n10_port, Q => 
                           n_1363, QN => n120_port);
   ID_EX_IMM_reg_31_inst : DFF_X1 port map( D => N209, CK => n10_port, Q => 
                           ID_EX_IMM_31_port, QN => n_1364);
   ID_EX_IMM_reg_30_inst : DFF_X1 port map( D => N208, CK => n10_port, Q => 
                           ID_EX_IMM_30_port, QN => n_1365);
   ID_EX_IMM_reg_29_inst : DFF_X1 port map( D => N207, CK => n10_port, Q => 
                           ID_EX_IMM_29_port, QN => n_1366);
   ID_EX_IMM_reg_28_inst : DFF_X1 port map( D => N206, CK => n10_port, Q => 
                           ID_EX_IMM_28_port, QN => n_1367);
   ID_EX_IMM_reg_27_inst : DFF_X1 port map( D => N205, CK => n10_port, Q => 
                           ID_EX_IMM_27_port, QN => n_1368);
   ID_EX_IMM_reg_26_inst : DFF_X1 port map( D => N204, CK => n10_port, Q => 
                           ID_EX_IMM_26_port, QN => n_1369);
   ID_EX_IMM_reg_25_inst : DFF_X1 port map( D => N203, CK => n10_port, Q => 
                           ID_EX_IMM_25_port, QN => n_1370);
   ID_EX_IMM_reg_24_inst : DFF_X1 port map( D => N202, CK => n10_port, Q => 
                           ID_EX_IMM_24_port, QN => n_1371);
   ID_EX_IMM_reg_23_inst : DFF_X1 port map( D => N201, CK => n10_port, Q => 
                           ID_EX_IMM_23_port, QN => n_1372);
   ID_EX_IMM_reg_22_inst : DFF_X1 port map( D => N200, CK => n10_port, Q => 
                           ID_EX_IMM_22_port, QN => n_1373);
   ID_EX_IMM_reg_21_inst : DFF_X1 port map( D => N199, CK => n10_port, Q => 
                           ID_EX_IMM_21_port, QN => n_1374);
   ID_EX_IMM_reg_20_inst : DFF_X1 port map( D => N198, CK => n10_port, Q => 
                           ID_EX_IMM_20_port, QN => n_1375);
   ID_EX_IMM_reg_19_inst : DFF_X1 port map( D => N197, CK => n10_port, Q => 
                           ID_EX_IMM_19_port, QN => n_1376);
   ID_EX_IMM_reg_18_inst : DFF_X1 port map( D => N196, CK => n10_port, Q => 
                           ID_EX_IMM_18_port, QN => n_1377);
   ID_EX_IMM_reg_17_inst : DFF_X1 port map( D => N195, CK => n10_port, Q => 
                           ID_EX_IMM_17_port, QN => n_1378);
   ID_EX_IMM_reg_16_inst : DFF_X1 port map( D => N194, CK => n9_port, Q => 
                           ID_EX_IMM_16_port, QN => n_1379);
   ID_EX_IMM_reg_15_inst : DFF_X1 port map( D => N193, CK => n10_port, Q => 
                           ID_EX_IMM_15_port, QN => n_1380);
   ID_EX_IMM_reg_14_inst : DFF_X1 port map( D => N192, CK => n10_port, Q => 
                           ID_EX_IMM_14_port, QN => n_1381);
   ID_EX_IMM_reg_13_inst : DFF_X1 port map( D => N191, CK => n10_port, Q => 
                           ID_EX_IMM_13_port, QN => n_1382);
   ID_EX_IMM_reg_12_inst : DFF_X1 port map( D => N190, CK => n10_port, Q => 
                           ID_EX_IMM_12_port, QN => n_1383);
   ID_EX_IMM_reg_11_inst : DFF_X1 port map( D => N189, CK => n10_port, Q => 
                           ID_EX_IMM_11_port, QN => n_1384);
   ID_EX_IMM_reg_10_inst : DFF_X1 port map( D => N188, CK => n10_port, Q => 
                           ID_EX_IMM_10_port, QN => n_1385);
   ID_EX_IMM_reg_9_inst : DFF_X1 port map( D => N187, CK => n10_port, Q => 
                           ID_EX_IMM_9_port, QN => n_1386);
   ID_EX_IMM_reg_8_inst : DFF_X1 port map( D => N186, CK => n10_port, Q => 
                           ID_EX_IMM_8_port, QN => n_1387);
   ID_EX_IMM_reg_7_inst : DFF_X1 port map( D => N185, CK => n10_port, Q => 
                           ID_EX_IMM_7_port, QN => n_1388);
   ID_EX_IMM_reg_6_inst : DFF_X1 port map( D => N184, CK => n10_port, Q => 
                           ID_EX_IMM_6_port, QN => n_1389);
   ID_EX_IMM_reg_5_inst : DFF_X1 port map( D => N183, CK => n10_port, Q => 
                           ID_EX_IMM_5_port, QN => n_1390);
   ID_EX_IMM_reg_4_inst : DFF_X1 port map( D => N182, CK => n10_port, Q => 
                           ID_EX_IMM_4_port, QN => n_1391);
   ID_EX_IMM_reg_3_inst : DFF_X1 port map( D => N181, CK => n10_port, Q => 
                           ID_EX_IMM_3_port, QN => n_1392);
   ID_EX_IMM_reg_2_inst : DFF_X1 port map( D => N180, CK => n10_port, Q => 
                           ID_EX_IMM_2_port, QN => n_1393);
   ID_EX_IMM_reg_1_inst : DFF_X1 port map( D => N179, CK => n10_port, Q => 
                           ID_EX_IMM_1_port, QN => n_1394);
   ID_EX_IMM_reg_0_inst : DFF_X1 port map( D => N178, CK => n10_port, Q => 
                           ID_EX_IMM_0_port, QN => n_1395);
   EX_MEM_RF_WE_reg : DFF_X1 port map( D => N242, CK => n11_port, Q => 
                           EX_MEM_RF_WE, QN => n83_port);
   EX_MEM_RD_reg_4_inst : DFF_X1 port map( D => N312, CK => n10_port, Q => 
                           EX_MEM_RD_4_port, QN => n46_port);
   EX_MEM_RD_reg_3_inst : DFF_X1 port map( D => N311, CK => n10_port, Q => 
                           EX_MEM_RD_3_port, QN => n47_port);
   EX_MEM_RD_reg_2_inst : DFF_X1 port map( D => N310, CK => n10_port, Q => 
                           EX_MEM_RD_2_port, QN => n48_port);
   EX_MEM_RD_reg_1_inst : DFF_X1 port map( D => N309, CK => n10_port, Q => 
                           EX_MEM_RD_1_port, QN => n49_port);
   EX_MEM_RD_reg_0_inst : DFF_X1 port map( D => N308, CK => n10_port, Q => 
                           EX_MEM_RD_0_port, QN => n50_port);
   MEM_WB_RF_WE_reg : DFF_X1 port map( D => N345, CK => n11_port, Q => 
                           MEM_WB_RF_WE, QN => n_1396);
   MEM_WB_DRAM_OUTPUT_reg_31_inst : DFF_X1 port map( D => N409, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_31_port, QN => n_1397);
   MEM_WB_DRAM_OUTPUT_reg_30_inst : DFF_X1 port map( D => N408, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_30_port, QN => n_1398);
   MEM_WB_DRAM_OUTPUT_reg_29_inst : DFF_X1 port map( D => N407, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_29_port, QN => n_1399);
   MEM_WB_DRAM_OUTPUT_reg_28_inst : DFF_X1 port map( D => N406, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_28_port, QN => n_1400);
   MEM_WB_DRAM_OUTPUT_reg_27_inst : DFF_X1 port map( D => N405, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_27_port, QN => n_1401);
   MEM_WB_DRAM_OUTPUT_reg_26_inst : DFF_X1 port map( D => N404, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_26_port, QN => n_1402);
   MEM_WB_DRAM_OUTPUT_reg_25_inst : DFF_X1 port map( D => N403, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_25_port, QN => n_1403);
   MEM_WB_DRAM_OUTPUT_reg_24_inst : DFF_X1 port map( D => N402, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_24_port, QN => n_1404);
   MEM_WB_DRAM_OUTPUT_reg_23_inst : DFF_X1 port map( D => N401, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_23_port, QN => n_1405);
   MEM_WB_DRAM_OUTPUT_reg_22_inst : DFF_X1 port map( D => N400, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_22_port, QN => n_1406);
   MEM_WB_DRAM_OUTPUT_reg_21_inst : DFF_X1 port map( D => N399, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_21_port, QN => n_1407);
   MEM_WB_DRAM_OUTPUT_reg_20_inst : DFF_X1 port map( D => N398, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_20_port, QN => n_1408);
   MEM_WB_DRAM_OUTPUT_reg_19_inst : DFF_X1 port map( D => N397, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_19_port, QN => n_1409);
   MEM_WB_DRAM_OUTPUT_reg_18_inst : DFF_X1 port map( D => N396, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_18_port, QN => n_1410);
   MEM_WB_DRAM_OUTPUT_reg_17_inst : DFF_X1 port map( D => N395, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_17_port, QN => n_1411);
   MEM_WB_DRAM_OUTPUT_reg_16_inst : DFF_X1 port map( D => N394, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_16_port, QN => n_1412);
   MEM_WB_DRAM_OUTPUT_reg_15_inst : DFF_X1 port map( D => N393, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_15_port, QN => n_1413);
   MEM_WB_DRAM_OUTPUT_reg_14_inst : DFF_X1 port map( D => N392, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_14_port, QN => n_1414);
   MEM_WB_DRAM_OUTPUT_reg_13_inst : DFF_X1 port map( D => N391, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_13_port, QN => n_1415);
   MEM_WB_DRAM_OUTPUT_reg_12_inst : DFF_X1 port map( D => N390, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_12_port, QN => n_1416);
   MEM_WB_DRAM_OUTPUT_reg_11_inst : DFF_X1 port map( D => N389, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_11_port, QN => n_1417);
   MEM_WB_DRAM_OUTPUT_reg_10_inst : DFF_X1 port map( D => N388, CK => n11_port,
                           Q => MEM_WB_DRAM_OUTPUT_10_port, QN => n_1418);
   MEM_WB_DRAM_OUTPUT_reg_9_inst : DFF_X1 port map( D => N387, CK => n11_port, 
                           Q => MEM_WB_DRAM_OUTPUT_9_port, QN => n_1419);
   MEM_WB_DRAM_OUTPUT_reg_8_inst : DFF_X1 port map( D => N386, CK => n11_port, 
                           Q => MEM_WB_DRAM_OUTPUT_8_port, QN => n_1420);
   MEM_WB_DRAM_OUTPUT_reg_7_inst : DFF_X1 port map( D => N385, CK => n11_port, 
                           Q => MEM_WB_DRAM_OUTPUT_7_port, QN => n_1421);
   MEM_WB_DRAM_OUTPUT_reg_6_inst : DFF_X1 port map( D => N384, CK => n11_port, 
                           Q => MEM_WB_DRAM_OUTPUT_6_port, QN => n_1422);
   MEM_WB_DRAM_OUTPUT_reg_5_inst : DFF_X1 port map( D => N383, CK => n11_port, 
                           Q => MEM_WB_DRAM_OUTPUT_5_port, QN => n_1423);
   MEM_WB_DRAM_OUTPUT_reg_4_inst : DFF_X1 port map( D => N382, CK => n11_port, 
                           Q => MEM_WB_DRAM_OUTPUT_4_port, QN => n_1424);
   MEM_WB_DRAM_OUTPUT_reg_3_inst : DFF_X1 port map( D => N381, CK => n11_port, 
                           Q => MEM_WB_DRAM_OUTPUT_3_port, QN => n_1425);
   MEM_WB_DRAM_OUTPUT_reg_2_inst : DFF_X1 port map( D => N380, CK => n11_port, 
                           Q => MEM_WB_DRAM_OUTPUT_2_port, QN => n_1426);
   MEM_WB_DRAM_OUTPUT_reg_1_inst : DFF_X1 port map( D => N379, CK => n11_port, 
                           Q => MEM_WB_DRAM_OUTPUT_1_port, QN => n_1427);
   MEM_WB_DRAM_OUTPUT_reg_0_inst : DFF_X1 port map( D => N378, CK => n9_port, Q
                           => MEM_WB_DRAM_OUTPUT_0_port, QN => n_1428);
   MEM_WB_RD_reg_4_inst : DFF_X1 port map( D => N414, CK => n10_port, Q => 
                           MEM_WB_RD_4_port, QN => n_1429);
   MEM_WB_RD_reg_3_inst : DFF_X1 port map( D => N413, CK => n10_port, Q => 
                           MEM_WB_RD_3_port, QN => n_1430);
   MEM_WB_RD_reg_2_inst : DFF_X1 port map( D => N412, CK => n10_port, Q => 
                           MEM_WB_RD_2_port, QN => n_1431);
   MEM_WB_RD_reg_1_inst : DFF_X1 port map( D => N411, CK => n10_port, Q => 
                           MEM_WB_RD_1_port, QN => n_1432);
   MEM_WB_RD_reg_0_inst : DFF_X1 port map( D => N410, CK => n10_port, Q => 
                           MEM_WB_RD_0_port, QN => n_1433);
   ID_EX_RF_OUT2_reg_0_inst : DFF_X1 port map( D => N146, CK => n11_port, Q => 
                           ID_EX_RF_OUT2_0_port, QN => n152_port);
   EX_MEM_RF_OUT2_reg_0_inst : DFF_X1 port map( D => N243, CK => n11_port, Q =>
                           DRAM_IN(0), QN => n_1434);
   ID_EX_RF_OUT2_reg_1_inst : DFF_X1 port map( D => N147, CK => n11_port, Q => 
                           ID_EX_RF_OUT2_1_port, QN => n151_port);
   EX_MEM_RF_OUT2_reg_1_inst : DFF_X1 port map( D => N244, CK => n9_port, Q => 
                           DRAM_IN(1), QN => n_1435);
   ID_EX_RF_OUT2_reg_2_inst : DFF_X1 port map( D => N148, CK => n10_port, Q => 
                           ID_EX_RF_OUT2_2_port, QN => n150_port);
   EX_MEM_RF_OUT2_reg_2_inst : DFF_X1 port map( D => N245, CK => n9_port, Q => 
                           DRAM_IN(2), QN => n_1436);
   ID_EX_RF_OUT2_reg_3_inst : DFF_X1 port map( D => N149, CK => n10_port, Q => 
                           ID_EX_RF_OUT2_3_port, QN => n149_port);
   EX_MEM_RF_OUT2_reg_3_inst : DFF_X1 port map( D => N246, CK => n9_port, Q => 
                           DRAM_IN(3), QN => n_1437);
   ID_EX_RF_OUT2_reg_4_inst : DFF_X1 port map( D => N150, CK => n11_port, Q => 
                           ID_EX_RF_OUT2_4_port, QN => n148_port);
   EX_MEM_RF_OUT2_reg_4_inst : DFF_X1 port map( D => N247, CK => n9_port, Q => 
                           DRAM_IN(4), QN => n_1438);
   ID_EX_RF_OUT2_reg_5_inst : DFF_X1 port map( D => N151, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_5_port, QN => n147_port);
   EX_MEM_RF_OUT2_reg_5_inst : DFF_X1 port map( D => N248, CK => n9_port, Q => 
                           DRAM_IN(5), QN => n_1439);
   ID_EX_RF_OUT2_reg_6_inst : DFF_X1 port map( D => N152, CK => n10_port, Q => 
                           ID_EX_RF_OUT2_6_port, QN => n146_port);
   EX_MEM_RF_OUT2_reg_6_inst : DFF_X1 port map( D => N249, CK => n9_port, Q => 
                           DRAM_IN(6), QN => n_1440);
   ID_EX_RF_OUT2_reg_7_inst : DFF_X1 port map( D => N153, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_7_port, QN => n145_port);
   EX_MEM_RF_OUT2_reg_7_inst : DFF_X1 port map( D => N250, CK => n9_port, Q => 
                           DRAM_IN(7), QN => n_1441);
   ID_EX_RF_OUT2_reg_8_inst : DFF_X1 port map( D => N154, CK => n11_port, Q => 
                           ID_EX_RF_OUT2_8_port, QN => n144_port);
   EX_MEM_RF_OUT2_reg_8_inst : DFF_X1 port map( D => N251, CK => n9_port, Q => 
                           DRAM_IN(8), QN => n_1442);
   ID_EX_RF_OUT2_reg_9_inst : DFF_X1 port map( D => N155, CK => n10_port, Q => 
                           ID_EX_RF_OUT2_9_port, QN => n143_port);
   EX_MEM_RF_OUT2_reg_9_inst : DFF_X1 port map( D => N252, CK => n9_port, Q => 
                           DRAM_IN(9), QN => n_1443);
   ID_EX_RF_OUT2_reg_10_inst : DFF_X1 port map( D => N156, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_10_port, QN => n142_port);
   EX_MEM_RF_OUT2_reg_10_inst : DFF_X1 port map( D => N253, CK => n9_port, Q =>
                           DRAM_IN(10), QN => n_1444);
   ID_EX_RF_OUT2_reg_11_inst : DFF_X1 port map( D => N157, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_11_port, QN => n141_port);
   EX_MEM_RF_OUT2_reg_11_inst : DFF_X1 port map( D => N254, CK => n9_port, Q =>
                           DRAM_IN(11), QN => n_1445);
   ID_EX_RF_OUT2_reg_12_inst : DFF_X1 port map( D => N158, CK => n11_port, Q =>
                           ID_EX_RF_OUT2_12_port, QN => n140_port);
   EX_MEM_RF_OUT2_reg_12_inst : DFF_X1 port map( D => N255, CK => n9_port, Q =>
                           DRAM_IN(12), QN => n_1446);
   ID_EX_RF_OUT2_reg_13_inst : DFF_X1 port map( D => N159, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_13_port, QN => n139_port);
   EX_MEM_RF_OUT2_reg_13_inst : DFF_X1 port map( D => N256, CK => n9_port, Q =>
                           DRAM_IN(13), QN => n_1447);
   ID_EX_RF_OUT2_reg_14_inst : DFF_X1 port map( D => N160, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_14_port, QN => n138_port);
   EX_MEM_RF_OUT2_reg_14_inst : DFF_X1 port map( D => N257, CK => n9_port, Q =>
                           DRAM_IN(14), QN => n_1448);
   ID_EX_RF_OUT2_reg_15_inst : DFF_X1 port map( D => N161, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_15_port, QN => n137_port);
   EX_MEM_RF_OUT2_reg_15_inst : DFF_X1 port map( D => N258, CK => n9_port, Q =>
                           DRAM_IN(15), QN => n_1449);
   ID_EX_RF_OUT2_reg_16_inst : DFF_X1 port map( D => N162, CK => n11_port, Q =>
                           ID_EX_RF_OUT2_16_port, QN => n136_port);
   EX_MEM_RF_OUT2_reg_16_inst : DFF_X1 port map( D => N259, CK => n9_port, Q =>
                           DRAM_IN(16), QN => n_1450);
   ID_EX_RF_OUT2_reg_17_inst : DFF_X1 port map( D => N163, CK => n10_port, Q =>
                           ID_EX_RF_OUT2_17_port, QN => n135_port);
   EX_MEM_RF_OUT2_reg_17_inst : DFF_X1 port map( D => N260, CK => n9_port, Q =>
                           DRAM_IN(17), QN => n_1451);
   ID_EX_RF_OUT2_reg_18_inst : DFF_X1 port map( D => N164, CK => n10_port, Q =>
                           ID_EX_RF_OUT2_18_port, QN => n134_port);
   EX_MEM_RF_OUT2_reg_18_inst : DFF_X1 port map( D => N261, CK => n9_port, Q =>
                           DRAM_IN(18), QN => n_1452);
   ID_EX_RF_OUT2_reg_19_inst : DFF_X1 port map( D => N165, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_19_port, QN => n133_port);
   EX_MEM_RF_OUT2_reg_19_inst : DFF_X1 port map( D => N262, CK => n9_port, Q =>
                           DRAM_IN(19), QN => n_1453);
   ID_EX_RF_OUT2_reg_20_inst : DFF_X1 port map( D => N166, CK => n11_port, Q =>
                           ID_EX_RF_OUT2_20_port, QN => n132_port);
   EX_MEM_RF_OUT2_reg_20_inst : DFF_X1 port map( D => N263, CK => n9_port, Q =>
                           DRAM_IN(20), QN => n_1454);
   ID_EX_RF_OUT2_reg_21_inst : DFF_X1 port map( D => N167, CK => n10_port, Q =>
                           ID_EX_RF_OUT2_21_port, QN => n131_port);
   EX_MEM_RF_OUT2_reg_21_inst : DFF_X1 port map( D => N264, CK => n9_port, Q =>
                           DRAM_IN(21), QN => n_1455);
   ID_EX_RF_OUT2_reg_22_inst : DFF_X1 port map( D => N168, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_22_port, QN => n130_port);
   EX_MEM_RF_OUT2_reg_22_inst : DFF_X1 port map( D => N265, CK => n9_port, Q =>
                           DRAM_IN(22), QN => n_1456);
   ID_EX_RF_OUT2_reg_23_inst : DFF_X1 port map( D => N169, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_23_port, QN => n129_port);
   EX_MEM_RF_OUT2_reg_23_inst : DFF_X1 port map( D => N266, CK => n9_port, Q =>
                           DRAM_IN(23), QN => n_1457);
   ID_EX_RF_OUT2_reg_24_inst : DFF_X1 port map( D => N170, CK => n11_port, Q =>
                           ID_EX_RF_OUT2_24_port, QN => n128_port);
   EX_MEM_RF_OUT2_reg_24_inst : DFF_X1 port map( D => N267, CK => n9_port, Q =>
                           DRAM_IN(24), QN => n_1458);
   ID_EX_RF_OUT2_reg_25_inst : DFF_X1 port map( D => N171, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_25_port, QN => n127_port);
   EX_MEM_RF_OUT2_reg_25_inst : DFF_X1 port map( D => N268, CK => n9_port, Q =>
                           DRAM_IN(25), QN => n_1459);
   ID_EX_RF_OUT2_reg_26_inst : DFF_X1 port map( D => N172, CK => n10_port, Q =>
                           ID_EX_RF_OUT2_26_port, QN => n126_port);
   EX_MEM_RF_OUT2_reg_26_inst : DFF_X1 port map( D => N269, CK => n9_port, Q =>
                           DRAM_IN(26), QN => n_1460);
   ID_EX_RF_OUT2_reg_27_inst : DFF_X1 port map( D => N173, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_27_port, QN => n125_port);
   EX_MEM_RF_OUT2_reg_27_inst : DFF_X1 port map( D => N270, CK => n9_port, Q =>
                           DRAM_IN(27), QN => n_1461);
   ID_EX_RF_OUT2_reg_28_inst : DFF_X1 port map( D => N174, CK => n11_port, Q =>
                           ID_EX_RF_OUT2_28_port, QN => n124_port);
   EX_MEM_RF_OUT2_reg_28_inst : DFF_X1 port map( D => N271, CK => n9_port, Q =>
                           DRAM_IN(28), QN => n_1462);
   ID_EX_RF_OUT2_reg_29_inst : DFF_X1 port map( D => N175, CK => n11_port, Q =>
                           ID_EX_RF_OUT2_29_port, QN => n123_port);
   EX_MEM_RF_OUT2_reg_29_inst : DFF_X1 port map( D => N272, CK => n9_port, Q =>
                           DRAM_IN(29), QN => n_1463);
   ID_EX_RF_OUT2_reg_30_inst : DFF_X1 port map( D => N176, CK => n11_port, Q =>
                           ID_EX_RF_OUT2_30_port, QN => n122_port);
   EX_MEM_RF_OUT2_reg_30_inst : DFF_X1 port map( D => N273, CK => n9_port, Q =>
                           DRAM_IN(30), QN => n_1464);
   ID_EX_RF_OUT2_reg_31_inst : DFF_X1 port map( D => N177, CK => n9_port, Q => 
                           ID_EX_RF_OUT2_31_port, QN => n121_port);
   EX_MEM_RF_OUT2_reg_31_inst : DFF_X1 port map( D => N274, CK => n9_port, Q =>
                           DRAM_IN(31), QN => n_1465);
   ID_EX_RF_OUT1_reg_0_inst : DFF_X1 port map( D => N114, CK => n10_port, Q => 
                           ID_EX_RF_OUT1_0_port, QN => n_1466);
   ID_EX_RF_OUT1_reg_1_inst : DFF_X1 port map( D => N115, CK => n10_port, Q => 
                           ID_EX_RF_OUT1_1_port, QN => n_1467);
   ID_EX_RF_OUT1_reg_2_inst : DFF_X1 port map( D => N116, CK => n10_port, Q => 
                           ID_EX_RF_OUT1_2_port, QN => n_1468);
   ID_EX_RF_OUT1_reg_3_inst : DFF_X1 port map( D => N117, CK => n10_port, Q => 
                           ID_EX_RF_OUT1_3_port, QN => n_1469);
   ID_EX_RF_OUT1_reg_4_inst : DFF_X1 port map( D => N118, CK => n10_port, Q => 
                           ID_EX_RF_OUT1_4_port, QN => n_1470);
   ID_EX_RF_OUT1_reg_5_inst : DFF_X1 port map( D => N119, CK => n9_port, Q => 
                           ID_EX_RF_OUT1_5_port, QN => n_1471);
   ID_EX_RF_OUT1_reg_6_inst : DFF_X1 port map( D => N120, CK => n10_port, Q => 
                           ID_EX_RF_OUT1_6_port, QN => n_1472);
   ID_EX_RF_OUT1_reg_7_inst : DFF_X1 port map( D => N121, CK => n10_port, Q => 
                           ID_EX_RF_OUT1_7_port, QN => n_1473);
   ID_EX_RF_OUT1_reg_8_inst : DFF_X1 port map( D => N122, CK => n10_port, Q => 
                           ID_EX_RF_OUT1_8_port, QN => n_1474);
   ID_EX_RF_OUT1_reg_9_inst : DFF_X1 port map( D => N123, CK => n10_port, Q => 
                           ID_EX_RF_OUT1_9_port, QN => n_1475);
   ID_EX_RF_OUT1_reg_10_inst : DFF_X1 port map( D => N124, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_10_port, QN => n_1476);
   ID_EX_RF_OUT1_reg_11_inst : DFF_X1 port map( D => N125, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_11_port, QN => n_1477);
   ID_EX_RF_OUT1_reg_12_inst : DFF_X1 port map( D => N126, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_12_port, QN => n_1478);
   ID_EX_RF_OUT1_reg_13_inst : DFF_X1 port map( D => N127, CK => n9_port, Q => 
                           ID_EX_RF_OUT1_13_port, QN => n_1479);
   ID_EX_RF_OUT1_reg_14_inst : DFF_X1 port map( D => N128, CK => n9_port, Q => 
                           ID_EX_RF_OUT1_14_port, QN => n_1480);
   ID_EX_RF_OUT1_reg_15_inst : DFF_X1 port map( D => N129, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_15_port, QN => n_1481);
   ID_EX_RF_OUT1_reg_16_inst : DFF_X1 port map( D => N130, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_16_port, QN => n_1482);
   ID_EX_RF_OUT1_reg_17_inst : DFF_X1 port map( D => N131, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_17_port, QN => n_1483);
   ID_EX_RF_OUT1_reg_18_inst : DFF_X1 port map( D => N132, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_18_port, QN => n_1484);
   ID_EX_RF_OUT1_reg_19_inst : DFF_X1 port map( D => N133, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_19_port, QN => n_1485);
   ID_EX_RF_OUT1_reg_20_inst : DFF_X1 port map( D => N134, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_20_port, QN => n_1486);
   ID_EX_RF_OUT1_reg_21_inst : DFF_X1 port map( D => N135, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_21_port, QN => n_1487);
   ID_EX_RF_OUT1_reg_22_inst : DFF_X1 port map( D => N136, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_22_port, QN => n_1488);
   ID_EX_RF_OUT1_reg_23_inst : DFF_X1 port map( D => N137, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_23_port, QN => n_1489);
   ID_EX_RF_OUT1_reg_24_inst : DFF_X1 port map( D => N138, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_24_port, QN => n_1490);
   ID_EX_RF_OUT1_reg_25_inst : DFF_X1 port map( D => N139, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_25_port, QN => n_1491);
   ID_EX_RF_OUT1_reg_26_inst : DFF_X1 port map( D => N140, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_26_port, QN => n_1492);
   ID_EX_RF_OUT1_reg_27_inst : DFF_X1 port map( D => N141, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_27_port, QN => n_1493);
   ID_EX_RF_OUT1_reg_28_inst : DFF_X1 port map( D => N142, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_28_port, QN => n_1494);
   ID_EX_RF_OUT1_reg_29_inst : DFF_X1 port map( D => N143, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_29_port, QN => n_1495);
   ID_EX_RF_OUT1_reg_30_inst : DFF_X1 port map( D => N144, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_30_port, QN => n_1496);
   ID_EX_RF_OUT1_reg_31_inst : DFF_X1 port map( D => N145, CK => n10_port, Q =>
                           ID_EX_RF_OUT1_31_port, QN => n_1497);
   EX_MEM_BRANCH_DETECT_reg : DFF_X1 port map( D => N307, CK => n10_port, Q => 
                           EX_MEM_BRANCH_DETECT, QN => n_1498);
   EX_MEM_ALU_OUTPUT_reg_0_inst : DFF_X1 port map( D => N275, CK => n11_port, Q
                           => ALU_OUT_0_port, QN => n82_port);
   MEM_WB_ALU_OUTPUT_reg_0_inst : DFF_X1 port map( D => N346, CK => n11_port, Q
                           => MEM_WB_ALU_OUTPUT_0_port, QN => n_1499);
   EX_MEM_ALU_OUTPUT_reg_1_inst : DFF_X1 port map( D => N276, CK => n10_port, Q
                           => ALU_OUT_1_port, QN => n81_port);
   MEM_WB_ALU_OUTPUT_reg_1_inst : DFF_X1 port map( D => N347, CK => n9_port, Q 
                           => MEM_WB_ALU_OUTPUT_1_port, QN => n_1500);
   EX_MEM_ALU_OUTPUT_reg_2_inst : DFF_X1 port map( D => N277, CK => n10_port, Q
                           => ALU_OUT_2_port, QN => n80_port);
   MEM_WB_ALU_OUTPUT_reg_2_inst : DFF_X1 port map( D => N348, CK => n10_port, Q
                           => MEM_WB_ALU_OUTPUT_2_port, QN => n_1501);
   EX_MEM_ALU_OUTPUT_reg_3_inst : DFF_X1 port map( D => N278, CK => n10_port, Q
                           => ALU_OUT_3_port, QN => n79_port);
   MEM_WB_ALU_OUTPUT_reg_3_inst : DFF_X1 port map( D => N349, CK => n10_port, Q
                           => MEM_WB_ALU_OUTPUT_3_port, QN => n_1502);
   EX_MEM_ALU_OUTPUT_reg_4_inst : DFF_X1 port map( D => N279, CK => n11_port, Q
                           => ALU_OUT_4_port, QN => n78_port);
   MEM_WB_ALU_OUTPUT_reg_4_inst : DFF_X1 port map( D => N350, CK => n11_port, Q
                           => MEM_WB_ALU_OUTPUT_4_port, QN => n_1503);
   EX_MEM_ALU_OUTPUT_reg_5_inst : DFF_X1 port map( D => N280, CK => n9_port, Q 
                           => ALU_OUT_5_port, QN => n77_port);
   MEM_WB_ALU_OUTPUT_reg_5_inst : DFF_X1 port map( D => N351, CK => n9_port, Q 
                           => MEM_WB_ALU_OUTPUT_5_port, QN => n_1504);
   EX_MEM_ALU_OUTPUT_reg_6_inst : DFF_X1 port map( D => N281, CK => n10_port, Q
                           => ALU_OUT_6_port, QN => n76_port);
   MEM_WB_ALU_OUTPUT_reg_6_inst : DFF_X1 port map( D => N352, CK => n10_port, Q
                           => MEM_WB_ALU_OUTPUT_6_port, QN => n_1505);
   EX_MEM_ALU_OUTPUT_reg_7_inst : DFF_X1 port map( D => N282, CK => n10_port, Q
                           => ALU_OUT_7_port, QN => n75_port);
   MEM_WB_ALU_OUTPUT_reg_7_inst : DFF_X1 port map( D => N353, CK => n10_port, Q
                           => MEM_WB_ALU_OUTPUT_7_port, QN => n_1506);
   EX_MEM_ALU_OUTPUT_reg_8_inst : DFF_X1 port map( D => N283, CK => n11_port, Q
                           => ALU_OUT_8_port, QN => n74_port);
   MEM_WB_ALU_OUTPUT_reg_8_inst : DFF_X1 port map( D => N354, CK => n11_port, Q
                           => MEM_WB_ALU_OUTPUT_8_port, QN => n_1507);
   EX_MEM_ALU_OUTPUT_reg_9_inst : DFF_X1 port map( D => N284, CK => n10_port, Q
                           => ALU_OUT_9_port, QN => n73_port);
   MEM_WB_ALU_OUTPUT_reg_9_inst : DFF_X1 port map( D => N355, CK => n10_port, Q
                           => MEM_WB_ALU_OUTPUT_9_port, QN => n_1508);
   EX_MEM_ALU_OUTPUT_reg_10_inst : DFF_X1 port map( D => N285, CK => n10_port, 
                           Q => ALU_OUT_10_port, QN => n72_port);
   MEM_WB_ALU_OUTPUT_reg_10_inst : DFF_X1 port map( D => N356, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_10_port, QN => n_1509);
   EX_MEM_ALU_OUTPUT_reg_11_inst : DFF_X1 port map( D => N286, CK => n10_port, 
                           Q => ALU_OUT_11_port, QN => n71_port);
   MEM_WB_ALU_OUTPUT_reg_11_inst : DFF_X1 port map( D => N357, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_11_port, QN => n_1510);
   EX_MEM_ALU_OUTPUT_reg_12_inst : DFF_X1 port map( D => N287, CK => n11_port, 
                           Q => ALU_OUT_12_port, QN => n70_port);
   MEM_WB_ALU_OUTPUT_reg_12_inst : DFF_X1 port map( D => N358, CK => n11_port, 
                           Q => MEM_WB_ALU_OUTPUT_12_port, QN => n_1511);
   EX_MEM_ALU_OUTPUT_reg_13_inst : DFF_X1 port map( D => N288, CK => n9_port, Q
                           => ALU_OUT_13_port, QN => n69_port);
   MEM_WB_ALU_OUTPUT_reg_13_inst : DFF_X1 port map( D => N359, CK => n9_port, Q
                           => MEM_WB_ALU_OUTPUT_13_port, QN => n_1512);
   EX_MEM_ALU_OUTPUT_reg_14_inst : DFF_X1 port map( D => N289, CK => n9_port, Q
                           => ALU_OUT_14_port, QN => n68_port);
   MEM_WB_ALU_OUTPUT_reg_14_inst : DFF_X1 port map( D => N360, CK => n9_port, Q
                           => MEM_WB_ALU_OUTPUT_14_port, QN => n_1513);
   EX_MEM_ALU_OUTPUT_reg_15_inst : DFF_X1 port map( D => N290, CK => n10_port, 
                           Q => ALU_OUT_15_port, QN => n67_port);
   MEM_WB_ALU_OUTPUT_reg_15_inst : DFF_X1 port map( D => N361, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_15_port, QN => n_1514);
   EX_MEM_ALU_OUTPUT_reg_16_inst : DFF_X1 port map( D => N291, CK => n11_port, 
                           Q => ALU_OUT_16_port, QN => n66_port);
   MEM_WB_ALU_OUTPUT_reg_16_inst : DFF_X1 port map( D => N362, CK => n11_port, 
                           Q => MEM_WB_ALU_OUTPUT_16_port, QN => n_1515);
   EX_MEM_ALU_OUTPUT_reg_17_inst : DFF_X1 port map( D => N292, CK => n10_port, 
                           Q => ALU_OUT_17_port, QN => n65_port);
   MEM_WB_ALU_OUTPUT_reg_17_inst : DFF_X1 port map( D => N363, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_17_port, QN => n_1516);
   EX_MEM_ALU_OUTPUT_reg_18_inst : DFF_X1 port map( D => N293, CK => n10_port, 
                           Q => ALU_OUT_18_port, QN => n64_port);
   MEM_WB_ALU_OUTPUT_reg_18_inst : DFF_X1 port map( D => N364, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_18_port, QN => n_1517);
   EX_MEM_ALU_OUTPUT_reg_19_inst : DFF_X1 port map( D => N294, CK => n10_port, 
                           Q => ALU_OUT_19_port, QN => n63_port);
   MEM_WB_ALU_OUTPUT_reg_19_inst : DFF_X1 port map( D => N365, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_19_port, QN => n_1518);
   EX_MEM_ALU_OUTPUT_reg_20_inst : DFF_X1 port map( D => N295, CK => n11_port, 
                           Q => ALU_OUT_20_port, QN => n62_port);
   MEM_WB_ALU_OUTPUT_reg_20_inst : DFF_X1 port map( D => N366, CK => n11_port, 
                           Q => MEM_WB_ALU_OUTPUT_20_port, QN => n_1519);
   EX_MEM_ALU_OUTPUT_reg_21_inst : DFF_X1 port map( D => N296, CK => n10_port, 
                           Q => ALU_OUT_21_port, QN => n61_port);
   MEM_WB_ALU_OUTPUT_reg_21_inst : DFF_X1 port map( D => N367, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_21_port, QN => n_1520);
   EX_MEM_ALU_OUTPUT_reg_22_inst : DFF_X1 port map( D => N297, CK => n10_port, 
                           Q => ALU_OUT_22_port, QN => n60_port);
   MEM_WB_ALU_OUTPUT_reg_22_inst : DFF_X1 port map( D => N368, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_22_port, QN => n_1521);
   EX_MEM_ALU_OUTPUT_reg_23_inst : DFF_X1 port map( D => N298, CK => n10_port, 
                           Q => ALU_OUT_23_port, QN => n59_port);
   MEM_WB_ALU_OUTPUT_reg_23_inst : DFF_X1 port map( D => N369, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_23_port, QN => n_1522);
   EX_MEM_ALU_OUTPUT_reg_24_inst : DFF_X1 port map( D => N299, CK => n11_port, 
                           Q => ALU_OUT_24_port, QN => n58_port);
   MEM_WB_ALU_OUTPUT_reg_24_inst : DFF_X1 port map( D => N370, CK => n11_port, 
                           Q => MEM_WB_ALU_OUTPUT_24_port, QN => n_1523);
   EX_MEM_ALU_OUTPUT_reg_25_inst : DFF_X1 port map( D => N300, CK => n10_port, 
                           Q => ALU_OUT_25_port, QN => n57_port);
   MEM_WB_ALU_OUTPUT_reg_25_inst : DFF_X1 port map( D => N371, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_25_port, QN => n_1524);
   EX_MEM_ALU_OUTPUT_reg_26_inst : DFF_X1 port map( D => N301, CK => n10_port, 
                           Q => ALU_OUT_26_port, QN => n56_port);
   MEM_WB_ALU_OUTPUT_reg_26_inst : DFF_X1 port map( D => N372, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_26_port, QN => n_1525);
   EX_MEM_ALU_OUTPUT_reg_27_inst : DFF_X1 port map( D => N302, CK => n10_port, 
                           Q => ALU_OUT_27_port, QN => n55_port);
   MEM_WB_ALU_OUTPUT_reg_27_inst : DFF_X1 port map( D => N373, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_27_port, QN => n_1526);
   EX_MEM_ALU_OUTPUT_reg_28_inst : DFF_X1 port map( D => N303, CK => n11_port, 
                           Q => ALU_OUT_28_port, QN => n54_port);
   MEM_WB_ALU_OUTPUT_reg_28_inst : DFF_X1 port map( D => N374, CK => n11_port, 
                           Q => MEM_WB_ALU_OUTPUT_28_port, QN => n_1527);
   EX_MEM_ALU_OUTPUT_reg_29_inst : DFF_X1 port map( D => N304, CK => n11_port, 
                           Q => ALU_OUT_29_port, QN => n53_port);
   MEM_WB_ALU_OUTPUT_reg_29_inst : DFF_X1 port map( D => N375, CK => n11_port, 
                           Q => MEM_WB_ALU_OUTPUT_29_port, QN => n_1528);
   EX_MEM_ALU_OUTPUT_reg_30_inst : DFF_X1 port map( D => N305, CK => n11_port, 
                           Q => ALU_OUT_30_port, QN => n52_port);
   MEM_WB_ALU_OUTPUT_reg_30_inst : DFF_X1 port map( D => N376, CK => n11_port, 
                           Q => MEM_WB_ALU_OUTPUT_30_port, QN => n_1529);
   EX_MEM_ALU_OUTPUT_reg_31_inst : DFF_X1 port map( D => N306, CK => n10_port, 
                           Q => ALU_OUT_31_port, QN => n51_port);
   IF_ID_NPC_reg_0_inst : DFF_X1 port map( D => N2, CK => n10_port, Q => n_1530
                           , QN => n45_port);
   ID_EX_NPC_reg_0_inst : DFF_X1 port map( D => N66, CK => n10_port, Q => 
                           ID_EX_NPC_0_port, QN => n185_port);
   EX_MEM_NPC_reg_0_inst : DFF_X1 port map( D => N210, CK => n10_port, Q => 
                           n_1531, QN => n115_port);
   MEM_WB_NPC_reg_0_inst : DFF_X1 port map( D => N313, CK => n10_port, Q => 
                           MEM_WB_NPC_0_port, QN => n_1532);
   IF_ID_NPC_reg_1_inst : DFF_X1 port map( D => N3, CK => n10_port, Q => n_1533
                           , QN => n44_port);
   ID_EX_NPC_reg_1_inst : DFF_X1 port map( D => N67, CK => n10_port, Q => 
                           ID_EX_NPC_1_port, QN => n184_port);
   EX_MEM_NPC_reg_1_inst : DFF_X1 port map( D => N211, CK => n9_port, Q => 
                           n_1534, QN => n114_port);
   MEM_WB_NPC_reg_1_inst : DFF_X1 port map( D => N314, CK => n9_port, Q => 
                           MEM_WB_NPC_1_port, QN => n_1535);
   IF_ID_NPC_reg_2_inst : DFF_X1 port map( D => N4, CK => n10_port, Q => n_1536
                           , QN => n43_port);
   ID_EX_NPC_reg_2_inst : DFF_X1 port map( D => N68, CK => n10_port, Q => 
                           ID_EX_NPC_2_port, QN => n183_port);
   EX_MEM_NPC_reg_2_inst : DFF_X1 port map( D => N212, CK => n10_port, Q => 
                           n_1537, QN => n113_port);
   MEM_WB_NPC_reg_2_inst : DFF_X1 port map( D => N315, CK => n10_port, Q => 
                           MEM_WB_NPC_2_port, QN => n_1538);
   IF_ID_NPC_reg_3_inst : DFF_X1 port map( D => N5, CK => n10_port, Q => n_1539
                           , QN => n42_port);
   ID_EX_NPC_reg_3_inst : DFF_X1 port map( D => N69, CK => n10_port, Q => 
                           ID_EX_NPC_3_port, QN => n182_port);
   EX_MEM_NPC_reg_3_inst : DFF_X1 port map( D => N213, CK => n10_port, Q => 
                           n_1540, QN => n112_port);
   MEM_WB_NPC_reg_3_inst : DFF_X1 port map( D => N316, CK => n10_port, Q => 
                           MEM_WB_NPC_3_port, QN => n_1541);
   IF_ID_NPC_reg_4_inst : DFF_X1 port map( D => N6, CK => n10_port, Q => n_1542
                           , QN => n41_port);
   ID_EX_NPC_reg_4_inst : DFF_X1 port map( D => N70, CK => n10_port, Q => 
                           ID_EX_NPC_4_port, QN => n181_port);
   EX_MEM_NPC_reg_4_inst : DFF_X1 port map( D => N214, CK => n10_port, Q => 
                           n_1543, QN => n111_port);
   MEM_WB_NPC_reg_4_inst : DFF_X1 port map( D => N317, CK => n10_port, Q => 
                           MEM_WB_NPC_4_port, QN => n_1544);
   IF_ID_NPC_reg_5_inst : DFF_X1 port map( D => N7, CK => n9_port, Q => n_1545,
                           QN => n40_port);
   ID_EX_NPC_reg_5_inst : DFF_X1 port map( D => N71, CK => n9_port, Q => 
                           ID_EX_NPC_5_port, QN => n180_port);
   EX_MEM_NPC_reg_5_inst : DFF_X1 port map( D => N215, CK => n9_port, Q => 
                           n_1546, QN => n110_port);
   MEM_WB_NPC_reg_5_inst : DFF_X1 port map( D => N318, CK => n9_port, Q => 
                           MEM_WB_NPC_5_port, QN => n_1547);
   IF_ID_NPC_reg_6_inst : DFF_X1 port map( D => N8, CK => n9_port, Q => n_1548,
                           QN => n39_port);
   ID_EX_NPC_reg_6_inst : DFF_X1 port map( D => N72, CK => n9_port, Q => 
                           ID_EX_NPC_6_port, QN => n179_port);
   EX_MEM_NPC_reg_6_inst : DFF_X1 port map( D => N216, CK => n9_port, Q => 
                           n_1549, QN => n109_port);
   MEM_WB_NPC_reg_6_inst : DFF_X1 port map( D => N319, CK => n9_port, Q => 
                           MEM_WB_NPC_6_port, QN => n_1550);
   IF_ID_NPC_reg_7_inst : DFF_X1 port map( D => N9, CK => n9_port, Q => n_1551,
                           QN => n38_port);
   ID_EX_NPC_reg_7_inst : DFF_X1 port map( D => N73, CK => n9_port, Q => 
                           ID_EX_NPC_7_port, QN => n178_port);
   EX_MEM_NPC_reg_7_inst : DFF_X1 port map( D => N217, CK => n9_port, Q => 
                           n_1552, QN => n108_port);
   MEM_WB_NPC_reg_7_inst : DFF_X1 port map( D => N320, CK => n9_port, Q => 
                           MEM_WB_NPC_7_port, QN => n_1553);
   IF_ID_NPC_reg_8_inst : DFF_X1 port map( D => N10, CK => n9_port, Q => n_1554
                           , QN => n37_port);
   ID_EX_NPC_reg_8_inst : DFF_X1 port map( D => N74, CK => n9_port, Q => 
                           ID_EX_NPC_8_port, QN => n177_port);
   EX_MEM_NPC_reg_8_inst : DFF_X1 port map( D => N218, CK => n9_port, Q => 
                           n_1555, QN => n107_port);
   MEM_WB_NPC_reg_8_inst : DFF_X1 port map( D => N321, CK => n9_port, Q => 
                           MEM_WB_NPC_8_port, QN => n_1556);
   IF_ID_NPC_reg_9_inst : DFF_X1 port map( D => N11, CK => n9_port, Q => n_1557
                           , QN => n36_port);
   ID_EX_NPC_reg_9_inst : DFF_X1 port map( D => N75, CK => n9_port, Q => 
                           ID_EX_NPC_9_port, QN => n176_port);
   EX_MEM_NPC_reg_9_inst : DFF_X1 port map( D => N219, CK => n9_port, Q => 
                           n_1558, QN => n106_port);
   MEM_WB_NPC_reg_9_inst : DFF_X1 port map( D => N322, CK => n9_port, Q => 
                           MEM_WB_NPC_9_port, QN => n_1559);
   IF_ID_NPC_reg_10_inst : DFF_X1 port map( D => N12, CK => n9_port, Q => 
                           n_1560, QN => n35_port);
   ID_EX_NPC_reg_10_inst : DFF_X1 port map( D => N76, CK => n9_port, Q => 
                           ID_EX_NPC_10_port, QN => n175_port);
   EX_MEM_NPC_reg_10_inst : DFF_X1 port map( D => N220, CK => n9_port, Q => 
                           n_1561, QN => n105_port);
   MEM_WB_NPC_reg_10_inst : DFF_X1 port map( D => N323, CK => n9_port, Q => 
                           MEM_WB_NPC_10_port, QN => n_1562);
   IF_ID_NPC_reg_11_inst : DFF_X1 port map( D => N13, CK => n9_port, Q => 
                           n_1563, QN => n34_port);
   ID_EX_NPC_reg_11_inst : DFF_X1 port map( D => N77, CK => n9_port, Q => 
                           ID_EX_NPC_11_port, QN => n174_port);
   EX_MEM_NPC_reg_11_inst : DFF_X1 port map( D => N221, CK => n9_port, Q => 
                           n_1564, QN => n104_port);
   MEM_WB_NPC_reg_11_inst : DFF_X1 port map( D => N324, CK => n9_port, Q => 
                           MEM_WB_NPC_11_port, QN => n_1565);
   IF_ID_NPC_reg_12_inst : DFF_X1 port map( D => N14, CK => n9_port, Q => 
                           n_1566, QN => n33_port);
   ID_EX_NPC_reg_12_inst : DFF_X1 port map( D => N78, CK => n9_port, Q => 
                           ID_EX_NPC_12_port, QN => n173_port);
   EX_MEM_NPC_reg_12_inst : DFF_X1 port map( D => N222, CK => n9_port, Q => 
                           n_1567, QN => n103_port);
   MEM_WB_NPC_reg_12_inst : DFF_X1 port map( D => N325, CK => n9_port, Q => 
                           MEM_WB_NPC_12_port, QN => n_1568);
   IF_ID_NPC_reg_13_inst : DFF_X1 port map( D => N15, CK => n9_port, Q => 
                           n_1569, QN => n32_port);
   ID_EX_NPC_reg_13_inst : DFF_X1 port map( D => N79, CK => n9_port, Q => 
                           ID_EX_NPC_13_port, QN => n172_port);
   EX_MEM_NPC_reg_13_inst : DFF_X1 port map( D => N223, CK => n9_port, Q => 
                           n_1570, QN => n102_port);
   MEM_WB_NPC_reg_13_inst : DFF_X1 port map( D => N326, CK => n9_port, Q => 
                           MEM_WB_NPC_13_port, QN => n_1571);
   IF_ID_NPC_reg_14_inst : DFF_X1 port map( D => N16, CK => n9_port, Q => 
                           n_1572, QN => n31_port);
   ID_EX_NPC_reg_14_inst : DFF_X1 port map( D => N80, CK => n9_port, Q => 
                           ID_EX_NPC_14_port, QN => n171_port);
   EX_MEM_NPC_reg_14_inst : DFF_X1 port map( D => N224, CK => n9_port, Q => 
                           n_1573, QN => n101_port);
   MEM_WB_NPC_reg_14_inst : DFF_X1 port map( D => N327, CK => n9_port, Q => 
                           MEM_WB_NPC_14_port, QN => n_1574);
   IF_ID_NPC_reg_15_inst : DFF_X1 port map( D => N17, CK => n9_port, Q => 
                           n_1575, QN => n30_port);
   ID_EX_NPC_reg_15_inst : DFF_X1 port map( D => N81, CK => n9_port, Q => 
                           ID_EX_NPC_15_port, QN => n170_port);
   EX_MEM_NPC_reg_15_inst : DFF_X1 port map( D => N225, CK => n9_port, Q => 
                           n_1576, QN => n100_port);
   MEM_WB_NPC_reg_15_inst : DFF_X1 port map( D => N328, CK => n9_port, Q => 
                           MEM_WB_NPC_15_port, QN => n_1577);
   IF_ID_NPC_reg_16_inst : DFF_X1 port map( D => N18, CK => n9_port, Q => 
                           n_1578, QN => n29_port);
   ID_EX_NPC_reg_16_inst : DFF_X1 port map( D => N82, CK => n9_port, Q => 
                           ID_EX_NPC_16_port, QN => n169_port);
   EX_MEM_NPC_reg_16_inst : DFF_X1 port map( D => N226, CK => n9_port, Q => 
                           n_1579, QN => n99_port);
   MEM_WB_NPC_reg_16_inst : DFF_X1 port map( D => N329, CK => n9_port, Q => 
                           MEM_WB_NPC_16_port, QN => n_1580);
   IF_ID_NPC_reg_17_inst : DFF_X1 port map( D => N19, CK => n9_port, Q => 
                           n_1581, QN => n28_port);
   ID_EX_NPC_reg_17_inst : DFF_X1 port map( D => N83, CK => n9_port, Q => 
                           ID_EX_NPC_17_port, QN => n168_port);
   EX_MEM_NPC_reg_17_inst : DFF_X1 port map( D => N227, CK => n9_port, Q => 
                           n_1582, QN => n98_port);
   MEM_WB_NPC_reg_17_inst : DFF_X1 port map( D => N330, CK => n9_port, Q => 
                           MEM_WB_NPC_17_port, QN => n_1583);
   IF_ID_NPC_reg_18_inst : DFF_X1 port map( D => N20, CK => n9_port, Q => 
                           n_1584, QN => n27_port);
   ID_EX_NPC_reg_18_inst : DFF_X1 port map( D => N84, CK => n9_port, Q => 
                           ID_EX_NPC_18_port, QN => n167_port);
   EX_MEM_NPC_reg_18_inst : DFF_X1 port map( D => N228, CK => n9_port, Q => 
                           n_1585, QN => n97_port);
   MEM_WB_NPC_reg_18_inst : DFF_X1 port map( D => N331, CK => n9_port, Q => 
                           MEM_WB_NPC_18_port, QN => n_1586);
   IF_ID_NPC_reg_19_inst : DFF_X1 port map( D => N21, CK => n9_port, Q => 
                           n_1587, QN => n26_port);
   ID_EX_NPC_reg_19_inst : DFF_X1 port map( D => N85, CK => n9_port, Q => 
                           ID_EX_NPC_19_port, QN => n166_port);
   EX_MEM_NPC_reg_19_inst : DFF_X1 port map( D => N229, CK => n9_port, Q => 
                           n_1588, QN => n96_port);
   MEM_WB_NPC_reg_19_inst : DFF_X1 port map( D => N332, CK => n9_port, Q => 
                           MEM_WB_NPC_19_port, QN => n_1589);
   IF_ID_NPC_reg_20_inst : DFF_X1 port map( D => N22, CK => n9_port, Q => 
                           n_1590, QN => n25_port);
   ID_EX_NPC_reg_20_inst : DFF_X1 port map( D => N86, CK => n9_port, Q => 
                           ID_EX_NPC_20_port, QN => n165_port);
   EX_MEM_NPC_reg_20_inst : DFF_X1 port map( D => N230, CK => n9_port, Q => 
                           n_1591, QN => n95_port);
   MEM_WB_NPC_reg_20_inst : DFF_X1 port map( D => N333, CK => n9_port, Q => 
                           MEM_WB_NPC_20_port, QN => n_1592);
   IF_ID_NPC_reg_21_inst : DFF_X1 port map( D => N23, CK => n9_port, Q => 
                           n_1593, QN => n24_port);
   ID_EX_NPC_reg_21_inst : DFF_X1 port map( D => N87, CK => n9_port, Q => 
                           ID_EX_NPC_21_port, QN => n164_port);
   EX_MEM_NPC_reg_21_inst : DFF_X1 port map( D => N231, CK => n9_port, Q => 
                           n_1594, QN => n94_port);
   MEM_WB_NPC_reg_21_inst : DFF_X1 port map( D => N334, CK => n9_port, Q => 
                           MEM_WB_NPC_21_port, QN => n_1595);
   IF_ID_NPC_reg_22_inst : DFF_X1 port map( D => N24, CK => n9_port, Q => 
                           n_1596, QN => n23_port);
   ID_EX_NPC_reg_22_inst : DFF_X1 port map( D => N88, CK => n9_port, Q => 
                           ID_EX_NPC_22_port, QN => n163_port);
   EX_MEM_NPC_reg_22_inst : DFF_X1 port map( D => N232, CK => n9_port, Q => 
                           n_1597, QN => n93_port);
   MEM_WB_NPC_reg_22_inst : DFF_X1 port map( D => N335, CK => n9_port, Q => 
                           MEM_WB_NPC_22_port, QN => n_1598);
   IF_ID_NPC_reg_23_inst : DFF_X1 port map( D => N25, CK => n9_port, Q => 
                           n_1599, QN => n22_port);
   ID_EX_NPC_reg_23_inst : DFF_X1 port map( D => N89, CK => n9_port, Q => 
                           ID_EX_NPC_23_port, QN => n162_port);
   EX_MEM_NPC_reg_23_inst : DFF_X1 port map( D => N233, CK => n9_port, Q => 
                           n_1600, QN => n92_port);
   MEM_WB_NPC_reg_23_inst : DFF_X1 port map( D => N336, CK => n9_port, Q => 
                           MEM_WB_NPC_23_port, QN => n_1601);
   IF_ID_NPC_reg_24_inst : DFF_X1 port map( D => N26, CK => n9_port, Q => 
                           n_1602, QN => n21_port);
   ID_EX_NPC_reg_24_inst : DFF_X1 port map( D => N90, CK => n9_port, Q => 
                           ID_EX_NPC_24_port, QN => n161_port);
   EX_MEM_NPC_reg_24_inst : DFF_X1 port map( D => N234, CK => n9_port, Q => 
                           n_1603, QN => n91_port);
   MEM_WB_NPC_reg_24_inst : DFF_X1 port map( D => N337, CK => n9_port, Q => 
                           MEM_WB_NPC_24_port, QN => n_1604);
   IF_ID_NPC_reg_25_inst : DFF_X1 port map( D => N27, CK => n9_port, Q => 
                           n_1605, QN => n20_port);
   ID_EX_NPC_reg_25_inst : DFF_X1 port map( D => N91, CK => n9_port, Q => 
                           ID_EX_NPC_25_port, QN => n160_port);
   EX_MEM_NPC_reg_25_inst : DFF_X1 port map( D => N235, CK => n9_port, Q => 
                           n_1606, QN => n90_port);
   MEM_WB_NPC_reg_25_inst : DFF_X1 port map( D => N338, CK => n9_port, Q => 
                           MEM_WB_NPC_25_port, QN => n_1607);
   IF_ID_NPC_reg_26_inst : DFF_X1 port map( D => N28, CK => n9_port, Q => 
                           n_1608, QN => n19_port);
   ID_EX_NPC_reg_26_inst : DFF_X1 port map( D => N92, CK => n9_port, Q => 
                           ID_EX_NPC_26_port, QN => n159_port);
   EX_MEM_NPC_reg_26_inst : DFF_X1 port map( D => N236, CK => n9_port, Q => 
                           n_1609, QN => n89_port);
   MEM_WB_NPC_reg_26_inst : DFF_X1 port map( D => N339, CK => n9_port, Q => 
                           MEM_WB_NPC_26_port, QN => n_1610);
   IF_ID_NPC_reg_27_inst : DFF_X1 port map( D => N29, CK => n9_port, Q => 
                           n_1611, QN => n18_port);
   ID_EX_NPC_reg_27_inst : DFF_X1 port map( D => N93, CK => n9_port, Q => 
                           ID_EX_NPC_27_port, QN => n158_port);
   EX_MEM_NPC_reg_27_inst : DFF_X1 port map( D => N237, CK => n9_port, Q => 
                           n_1612, QN => n88_port);
   MEM_WB_NPC_reg_27_inst : DFF_X1 port map( D => N340, CK => n9_port, Q => 
                           MEM_WB_NPC_27_port, QN => n_1613);
   IF_ID_NPC_reg_28_inst : DFF_X1 port map( D => N30, CK => n9_port, Q => 
                           n_1614, QN => n17_port);
   ID_EX_NPC_reg_28_inst : DFF_X1 port map( D => N94, CK => n9_port, Q => 
                           ID_EX_NPC_28_port, QN => n157_port);
   EX_MEM_NPC_reg_28_inst : DFF_X1 port map( D => N238, CK => n9_port, Q => 
                           n_1615, QN => n87_port);
   MEM_WB_NPC_reg_28_inst : DFF_X1 port map( D => N341, CK => n9_port, Q => 
                           MEM_WB_NPC_28_port, QN => n_1616);
   IF_ID_NPC_reg_29_inst : DFF_X1 port map( D => N31, CK => n9_port, Q => 
                           n_1617, QN => n16_port);
   ID_EX_NPC_reg_29_inst : DFF_X1 port map( D => N95, CK => n9_port, Q => 
                           ID_EX_NPC_29_port, QN => n156_port);
   EX_MEM_NPC_reg_29_inst : DFF_X1 port map( D => N239, CK => n9_port, Q => 
                           n_1618, QN => n86_port);
   MEM_WB_NPC_reg_29_inst : DFF_X1 port map( D => N342, CK => n9_port, Q => 
                           MEM_WB_NPC_29_port, QN => n_1619);
   IF_ID_NPC_reg_30_inst : DFF_X1 port map( D => N32, CK => n9_port, Q => 
                           n_1620, QN => n15_port);
   ID_EX_NPC_reg_30_inst : DFF_X1 port map( D => N96, CK => n9_port, Q => 
                           ID_EX_NPC_30_port, QN => n155_port);
   EX_MEM_NPC_reg_30_inst : DFF_X1 port map( D => N240, CK => n9_port, Q => 
                           n_1621, QN => n85_port);
   MEM_WB_NPC_reg_30_inst : DFF_X1 port map( D => N343, CK => n9_port, Q => 
                           MEM_WB_NPC_30_port, QN => n_1622);
   IF_ID_NPC_reg_31_inst : DFF_X1 port map( D => N33, CK => n9_port, Q => 
                           n_1623, QN => n14_port);
   ID_EX_NPC_reg_31_inst : DFF_X1 port map( D => N97, CK => n9_port, Q => 
                           ID_EX_NPC_31_port, QN => n154_port);
   EX_MEM_NPC_reg_31_inst : DFF_X1 port map( D => N241, CK => n9_port, Q => 
                           n_1624, QN => n84_port);
   MEM_WB_NPC_reg_31_inst : DFF_X1 port map( D => N344, CK => n9_port, Q => 
                           MEM_WB_NPC_31_port, QN => n_1625);
   MEM_WB_ALU_OUTPUT_reg_31_inst : DFF_X1 port map( D => N377, CK => n10_port, 
                           Q => MEM_WB_ALU_OUTPUT_31_port, QN => n_1626);
   PROGRAM_COUNTER : FFDR_N32 port map( CLK => n9_port, RST => RST, EN => 
                           PC_LATCH_EN, REGIN(31) => PC_BUS_31_port, REGIN(30) 
                           => PC_BUS_30_port, REGIN(29) => PC_BUS_29_port, 
                           REGIN(28) => PC_BUS_28_port, REGIN(27) => 
                           PC_BUS_27_port, REGIN(26) => PC_BUS_26_port, 
                           REGIN(25) => PC_BUS_25_port, REGIN(24) => 
                           PC_BUS_24_port, REGIN(23) => PC_BUS_23_port, 
                           REGIN(22) => PC_BUS_22_port, REGIN(21) => 
                           PC_BUS_21_port, REGIN(20) => PC_BUS_20_port, 
                           REGIN(19) => PC_BUS_19_port, REGIN(18) => 
                           PC_BUS_18_port, REGIN(17) => PC_BUS_17_port, 
                           REGIN(16) => PC_BUS_16_port, REGIN(15) => 
                           PC_BUS_15_port, REGIN(14) => PC_BUS_14_port, 
                           REGIN(13) => PC_BUS_13_port, REGIN(12) => 
                           PC_BUS_12_port, REGIN(11) => PC_BUS_11_port, 
                           REGIN(10) => PC_BUS_10_port, REGIN(9) => 
                           PC_BUS_9_port, REGIN(8) => PC_BUS_8_port, REGIN(7) 
                           => PC_BUS_7_port, REGIN(6) => PC_BUS_6_port, 
                           REGIN(5) => PC_BUS_5_port, REGIN(4) => PC_BUS_4_port
                           , REGIN(3) => PC_BUS_3_port, REGIN(2) => 
                           PC_BUS_2_port, REGIN(1) => PC_BUS_1_port, REGIN(0) 
                           => PC_BUS_0_port, REGOUT(31) => PC_OUT_31_port, 
                           REGOUT(30) => PC_OUT_30_port, REGOUT(29) => 
                           PC_OUT_29_port, REGOUT(28) => PC_OUT_28_port, 
                           REGOUT(27) => PC_OUT_27_port, REGOUT(26) => 
                           PC_OUT_26_port, REGOUT(25) => PC_OUT_25_port, 
                           REGOUT(24) => PC_OUT_24_port, REGOUT(23) => 
                           PC_OUT_23_port, REGOUT(22) => PC_OUT_22_port, 
                           REGOUT(21) => PC_OUT_21_port, REGOUT(20) => 
                           PC_OUT_20_port, REGOUT(19) => PC_OUT_19_port, 
                           REGOUT(18) => PC_OUT_18_port, REGOUT(17) => 
                           PC_OUT_17_port, REGOUT(16) => PC_OUT_16_port, 
                           REGOUT(15) => PC_OUT_15_port, REGOUT(14) => 
                           PC_OUT_14_port, REGOUT(13) => PC_OUT_13_port, 
                           REGOUT(12) => PC_OUT_12_port, REGOUT(11) => 
                           PC_OUT_11_port, REGOUT(10) => PC_OUT_10_port, 
                           REGOUT(9) => PC_OUT_9_port, REGOUT(8) => 
                           PC_OUT_8_port, REGOUT(7) => PC_OUT_7_port, REGOUT(6)
                           => PC_OUT_6_port, REGOUT(5) => PC_OUT_5_port, 
                           REGOUT(4) => PC_OUT_4_port, REGOUT(3) => 
                           PC_OUT_3_port, REGOUT(2) => PC_OUT_2_port, REGOUT(1)
                           => PC_OUT_1_port, REGOUT(0) => PC_OUT_0_port);
   PC_MUX : MUX21_N32_4 port map( A(31) => NPC_BUS_31_port, A(30) => 
                           NPC_BUS_30_port, A(29) => NPC_BUS_29_port, A(28) => 
                           NPC_BUS_28_port, A(27) => NPC_BUS_27_port, A(26) => 
                           NPC_BUS_26_port, A(25) => NPC_BUS_25_port, A(24) => 
                           NPC_BUS_24_port, A(23) => NPC_BUS_23_port, A(22) => 
                           NPC_BUS_22_port, A(21) => NPC_BUS_21_port, A(20) => 
                           NPC_BUS_20_port, A(19) => NPC_BUS_19_port, A(18) => 
                           NPC_BUS_18_port, A(17) => NPC_BUS_17_port, A(16) => 
                           NPC_BUS_16_port, A(15) => NPC_BUS_15_port, A(14) => 
                           NPC_BUS_14_port, A(13) => NPC_BUS_13_port, A(12) => 
                           NPC_BUS_12_port, A(11) => NPC_BUS_11_port, A(10) => 
                           NPC_BUS_10_port, A(9) => NPC_BUS_9_port, A(8) => 
                           NPC_BUS_8_port, A(7) => NPC_BUS_7_port, A(6) => 
                           NPC_BUS_6_port, A(5) => NPC_BUS_5_port, A(4) => 
                           NPC_BUS_4_port, A(3) => NPC_BUS_3_port, A(2) => 
                           NPC_BUS_2_port, A(1) => NPC_BUS_1_port, A(0) => 
                           NPC_BUS_0_port, B(31) => ALU_OUT_31_port, B(30) => 
                           ALU_OUT_30_port, B(29) => ALU_OUT_29_port, B(28) => 
                           ALU_OUT_28_port, B(27) => ALU_OUT_27_port, B(26) => 
                           ALU_OUT_26_port, B(25) => ALU_OUT_25_port, B(24) => 
                           ALU_OUT_24_port, B(23) => ALU_OUT_23_port, B(22) => 
                           ALU_OUT_22_port, B(21) => ALU_OUT_21_port, B(20) => 
                           ALU_OUT_20_port, B(19) => ALU_OUT_19_port, B(18) => 
                           ALU_OUT_18_port, B(17) => ALU_OUT_17_port, B(16) => 
                           ALU_OUT_16_port, B(15) => ALU_OUT_15_port, B(14) => 
                           ALU_OUT_14_port, B(13) => ALU_OUT_13_port, B(12) => 
                           ALU_OUT_12_port, B(11) => ALU_OUT_11_port, B(10) => 
                           ALU_OUT_10_port, B(9) => ALU_OUT_9_port, B(8) => 
                           ALU_OUT_8_port, B(7) => ALU_OUT_7_port, B(6) => 
                           ALU_OUT_6_port, B(5) => ALU_OUT_5_port, B(4) => 
                           ALU_OUT_4_port, B(3) => ALU_OUT_3_port, B(2) => 
                           ALU_OUT_2_port, B(1) => ALU_OUT_1_port, B(0) => 
                           ALU_OUT_0_port, S => n187_port, Y(31) => 
                           PC_BUS_31_port, Y(30) => PC_BUS_30_port, Y(29) => 
                           PC_BUS_29_port, Y(28) => PC_BUS_28_port, Y(27) => 
                           PC_BUS_27_port, Y(26) => PC_BUS_26_port, Y(25) => 
                           PC_BUS_25_port, Y(24) => PC_BUS_24_port, Y(23) => 
                           PC_BUS_23_port, Y(22) => PC_BUS_22_port, Y(21) => 
                           PC_BUS_21_port, Y(20) => PC_BUS_20_port, Y(19) => 
                           PC_BUS_19_port, Y(18) => PC_BUS_18_port, Y(17) => 
                           PC_BUS_17_port, Y(16) => PC_BUS_16_port, Y(15) => 
                           PC_BUS_15_port, Y(14) => PC_BUS_14_port, Y(13) => 
                           PC_BUS_13_port, Y(12) => PC_BUS_12_port, Y(11) => 
                           PC_BUS_11_port, Y(10) => PC_BUS_10_port, Y(9) => 
                           PC_BUS_9_port, Y(8) => PC_BUS_8_port, Y(7) => 
                           PC_BUS_7_port, Y(6) => PC_BUS_6_port, Y(5) => 
                           PC_BUS_5_port, Y(4) => PC_BUS_4_port, Y(3) => 
                           PC_BUS_3_port, Y(2) => PC_BUS_2_port, Y(1) => 
                           PC_BUS_1_port, Y(0) => PC_BUS_0_port);
   NEXT_PROGRAM_COUNTER : LDR_N32_6 port map( RST => RST, EN => NPC_LATCH_EN, 
                           REGIN(31) => PC_BUS_31_port, REGIN(30) => 
                           PC_BUS_30_port, REGIN(29) => PC_BUS_29_port, 
                           REGIN(28) => PC_BUS_28_port, REGIN(27) => 
                           PC_BUS_27_port, REGIN(26) => PC_BUS_26_port, 
                           REGIN(25) => PC_BUS_25_port, REGIN(24) => 
                           PC_BUS_24_port, REGIN(23) => PC_BUS_23_port, 
                           REGIN(22) => PC_BUS_22_port, REGIN(21) => 
                           PC_BUS_21_port, REGIN(20) => PC_BUS_20_port, 
                           REGIN(19) => PC_BUS_19_port, REGIN(18) => 
                           PC_BUS_18_port, REGIN(17) => PC_BUS_17_port, 
                           REGIN(16) => PC_BUS_16_port, REGIN(15) => 
                           PC_BUS_15_port, REGIN(14) => PC_BUS_14_port, 
                           REGIN(13) => PC_BUS_13_port, REGIN(12) => 
                           PC_BUS_12_port, REGIN(11) => PC_BUS_11_port, 
                           REGIN(10) => PC_BUS_10_port, REGIN(9) => 
                           PC_BUS_9_port, REGIN(8) => PC_BUS_8_port, REGIN(7) 
                           => PC_BUS_7_port, REGIN(6) => PC_BUS_6_port, 
                           REGIN(5) => PC_BUS_5_port, REGIN(4) => PC_BUS_4_port
                           , REGIN(3) => PC_BUS_3_port, REGIN(2) => 
                           PC_BUS_2_port, REGIN(1) => PC_BUS_1_port, REGIN(0) 
                           => PC_BUS_0_port, REGOUT(31) => 
                           IF_ID_NPC_NEXT_31_port, REGOUT(30) => 
                           IF_ID_NPC_NEXT_30_port, REGOUT(29) => 
                           IF_ID_NPC_NEXT_29_port, REGOUT(28) => 
                           IF_ID_NPC_NEXT_28_port, REGOUT(27) => 
                           IF_ID_NPC_NEXT_27_port, REGOUT(26) => 
                           IF_ID_NPC_NEXT_26_port, REGOUT(25) => 
                           IF_ID_NPC_NEXT_25_port, REGOUT(24) => 
                           IF_ID_NPC_NEXT_24_port, REGOUT(23) => 
                           IF_ID_NPC_NEXT_23_port, REGOUT(22) => 
                           IF_ID_NPC_NEXT_22_port, REGOUT(21) => 
                           IF_ID_NPC_NEXT_21_port, REGOUT(20) => 
                           IF_ID_NPC_NEXT_20_port, REGOUT(19) => 
                           IF_ID_NPC_NEXT_19_port, REGOUT(18) => 
                           IF_ID_NPC_NEXT_18_port, REGOUT(17) => 
                           IF_ID_NPC_NEXT_17_port, REGOUT(16) => 
                           IF_ID_NPC_NEXT_16_port, REGOUT(15) => 
                           IF_ID_NPC_NEXT_15_port, REGOUT(14) => 
                           IF_ID_NPC_NEXT_14_port, REGOUT(13) => 
                           IF_ID_NPC_NEXT_13_port, REGOUT(12) => 
                           IF_ID_NPC_NEXT_12_port, REGOUT(11) => 
                           IF_ID_NPC_NEXT_11_port, REGOUT(10) => 
                           IF_ID_NPC_NEXT_10_port, REGOUT(9) => 
                           IF_ID_NPC_NEXT_9_port, REGOUT(8) => 
                           IF_ID_NPC_NEXT_8_port, REGOUT(7) => 
                           IF_ID_NPC_NEXT_7_port, REGOUT(6) => 
                           IF_ID_NPC_NEXT_6_port, REGOUT(5) => 
                           IF_ID_NPC_NEXT_5_port, REGOUT(4) => 
                           IF_ID_NPC_NEXT_4_port, REGOUT(3) => 
                           IF_ID_NPC_NEXT_3_port, REGOUT(2) => 
                           IF_ID_NPC_NEXT_2_port, REGOUT(1) => 
                           IF_ID_NPC_NEXT_1_port, REGOUT(0) => 
                           IF_ID_NPC_NEXT_0_port);
   INSTRUCTION_REGISTER : LDR_N32_5 port map( RST => RST, EN => IR_LATCH_EN, 
                           REGIN(31) => IR_IN(31), REGIN(30) => IR_IN(30), 
                           REGIN(29) => IR_IN(29), REGIN(28) => IR_IN(28), 
                           REGIN(27) => IR_IN(27), REGIN(26) => IR_IN(26), 
                           REGIN(25) => IR_IN(25), REGIN(24) => IR_IN(24), 
                           REGIN(23) => IR_IN(23), REGIN(22) => IR_IN(22), 
                           REGIN(21) => IR_IN(21), REGIN(20) => IR_IN(20), 
                           REGIN(19) => IR_IN(19), REGIN(18) => IR_IN(18), 
                           REGIN(17) => IR_IN(17), REGIN(16) => IR_IN(16), 
                           REGIN(15) => IR_IN(15), REGIN(14) => IR_IN(14), 
                           REGIN(13) => IR_IN(13), REGIN(12) => IR_IN(12), 
                           REGIN(11) => IR_IN(11), REGIN(10) => IR_IN(10), 
                           REGIN(9) => IR_IN(9), REGIN(8) => IR_IN(8), REGIN(7)
                           => IR_IN(7), REGIN(6) => IR_IN(6), REGIN(5) => 
                           IR_IN(5), REGIN(4) => IR_IN(4), REGIN(3) => IR_IN(3)
                           , REGIN(2) => IR_IN(2), REGIN(1) => IR_IN(1), 
                           REGIN(0) => IR_IN(0), REGOUT(31) => IR_OUT_31_port, 
                           REGOUT(30) => IR_OUT_30_port, REGOUT(29) => 
                           IR_OUT_29_port, REGOUT(28) => IR_OUT_28_port, 
                           REGOUT(27) => IR_OUT_27_port, REGOUT(26) => 
                           IR_OUT_26_port, REGOUT(25) => IR_OUT_25_port, 
                           REGOUT(24) => IR_OUT_24_port, REGOUT(23) => 
                           IR_OUT_23_port, REGOUT(22) => IR_OUT_22_port, 
                           REGOUT(21) => IR_OUT_21_port, REGOUT(20) => 
                           IR_OUT_20_port, REGOUT(19) => IR_OUT_19_port, 
                           REGOUT(18) => IR_OUT_18_port, REGOUT(17) => 
                           IR_OUT_17_port, REGOUT(16) => IR_OUT_16_port, 
                           REGOUT(15) => IR_OUT_15_port, REGOUT(14) => 
                           IR_OUT_14_port, REGOUT(13) => IR_OUT_13_port, 
                           REGOUT(12) => IR_OUT_12_port, REGOUT(11) => 
                           IR_OUT_11_port, REGOUT(10) => IR_OUT_10_port, 
                           REGOUT(9) => IR_OUT_9_port, REGOUT(8) => 
                           IR_OUT_8_port, REGOUT(7) => IR_OUT_7_port, REGOUT(6)
                           => IR_OUT_6_port, REGOUT(5) => IR_OUT_5_port, 
                           REGOUT(4) => IR_OUT_4_port, REGOUT(3) => 
                           IR_OUT_3_port, REGOUT(2) => IR_OUT_2_port, REGOUT(1)
                           => IR_OUT_1_port, REGOUT(0) => IR_OUT_0_port);
   REGISTER_FILE : RF_N32_NA5 port map( RST => RST, EN => X_Logic1_port, EN_RD1
                           => X_Logic1_port, EN_RD2 => X_Logic1_port, EN_WR => 
                           MEM_WB_RF_WE, ADD_RD1(4) => ID_EX_RS1_NEXT_4_port, 
                           ADD_RD1(3) => ID_EX_RS1_NEXT_3_port, ADD_RD1(2) => 
                           ID_EX_RS1_NEXT_2_port, ADD_RD1(1) => 
                           ID_EX_RS1_NEXT_1_port, ADD_RD1(0) => 
                           ID_EX_RS1_NEXT_0_port, ADD_RD2(4) => 
                           ID_EX_RS2_NEXT_4_port, ADD_RD2(3) => 
                           ID_EX_RS2_NEXT_3_port, ADD_RD2(2) => 
                           ID_EX_RS2_NEXT_2_port, ADD_RD2(1) => 
                           ID_EX_RS2_NEXT_1_port, ADD_RD2(0) => 
                           ID_EX_RS2_NEXT_0_port, ADD_WR(4) => MEM_WB_RD_4_port
                           , ADD_WR(3) => MEM_WB_RD_3_port, ADD_WR(2) => 
                           MEM_WB_RD_2_port, ADD_WR(1) => MEM_WB_RD_1_port, 
                           ADD_WR(0) => MEM_WB_RD_0_port, DATAIN(31) => 
                           JAL_MUX_OUT_31_port, DATAIN(30) => 
                           JAL_MUX_OUT_30_port, DATAIN(29) => 
                           JAL_MUX_OUT_29_port, DATAIN(28) => 
                           JAL_MUX_OUT_28_port, DATAIN(27) => 
                           JAL_MUX_OUT_27_port, DATAIN(26) => 
                           JAL_MUX_OUT_26_port, DATAIN(25) => 
                           JAL_MUX_OUT_25_port, DATAIN(24) => 
                           JAL_MUX_OUT_24_port, DATAIN(23) => 
                           JAL_MUX_OUT_23_port, DATAIN(22) => 
                           JAL_MUX_OUT_22_port, DATAIN(21) => 
                           JAL_MUX_OUT_21_port, DATAIN(20) => 
                           JAL_MUX_OUT_20_port, DATAIN(19) => 
                           JAL_MUX_OUT_19_port, DATAIN(18) => 
                           JAL_MUX_OUT_18_port, DATAIN(17) => 
                           JAL_MUX_OUT_17_port, DATAIN(16) => 
                           JAL_MUX_OUT_16_port, DATAIN(15) => 
                           JAL_MUX_OUT_15_port, DATAIN(14) => 
                           JAL_MUX_OUT_14_port, DATAIN(13) => 
                           JAL_MUX_OUT_13_port, DATAIN(12) => 
                           JAL_MUX_OUT_12_port, DATAIN(11) => 
                           JAL_MUX_OUT_11_port, DATAIN(10) => 
                           JAL_MUX_OUT_10_port, DATAIN(9) => JAL_MUX_OUT_9_port
                           , DATAIN(8) => JAL_MUX_OUT_8_port, DATAIN(7) => 
                           JAL_MUX_OUT_7_port, DATAIN(6) => JAL_MUX_OUT_6_port,
                           DATAIN(5) => JAL_MUX_OUT_5_port, DATAIN(4) => 
                           JAL_MUX_OUT_4_port, DATAIN(3) => JAL_MUX_OUT_3_port,
                           DATAIN(2) => JAL_MUX_OUT_2_port, DATAIN(1) => 
                           JAL_MUX_OUT_1_port, DATAIN(0) => JAL_MUX_OUT_0_port,
                           OUT1(31) => RF_OUT1_31_port, OUT1(30) => 
                           RF_OUT1_30_port, OUT1(29) => RF_OUT1_29_port, 
                           OUT1(28) => RF_OUT1_28_port, OUT1(27) => 
                           RF_OUT1_27_port, OUT1(26) => RF_OUT1_26_port, 
                           OUT1(25) => RF_OUT1_25_port, OUT1(24) => 
                           RF_OUT1_24_port, OUT1(23) => RF_OUT1_23_port, 
                           OUT1(22) => RF_OUT1_22_port, OUT1(21) => 
                           RF_OUT1_21_port, OUT1(20) => RF_OUT1_20_port, 
                           OUT1(19) => RF_OUT1_19_port, OUT1(18) => 
                           RF_OUT1_18_port, OUT1(17) => RF_OUT1_17_port, 
                           OUT1(16) => RF_OUT1_16_port, OUT1(15) => 
                           RF_OUT1_15_port, OUT1(14) => RF_OUT1_14_port, 
                           OUT1(13) => RF_OUT1_13_port, OUT1(12) => 
                           RF_OUT1_12_port, OUT1(11) => RF_OUT1_11_port, 
                           OUT1(10) => RF_OUT1_10_port, OUT1(9) => 
                           RF_OUT1_9_port, OUT1(8) => RF_OUT1_8_port, OUT1(7) 
                           => RF_OUT1_7_port, OUT1(6) => RF_OUT1_6_port, 
                           OUT1(5) => RF_OUT1_5_port, OUT1(4) => RF_OUT1_4_port
                           , OUT1(3) => RF_OUT1_3_port, OUT1(2) => 
                           RF_OUT1_2_port, OUT1(1) => RF_OUT1_1_port, OUT1(0) 
                           => RF_OUT1_0_port, OUT2(31) => RF_OUT2_31_port, 
                           OUT2(30) => RF_OUT2_30_port, OUT2(29) => 
                           RF_OUT2_29_port, OUT2(28) => RF_OUT2_28_port, 
                           OUT2(27) => RF_OUT2_27_port, OUT2(26) => 
                           RF_OUT2_26_port, OUT2(25) => RF_OUT2_25_port, 
                           OUT2(24) => RF_OUT2_24_port, OUT2(23) => 
                           RF_OUT2_23_port, OUT2(22) => RF_OUT2_22_port, 
                           OUT2(21) => RF_OUT2_21_port, OUT2(20) => 
                           RF_OUT2_20_port, OUT2(19) => RF_OUT2_19_port, 
                           OUT2(18) => RF_OUT2_18_port, OUT2(17) => 
                           RF_OUT2_17_port, OUT2(16) => RF_OUT2_16_port, 
                           OUT2(15) => RF_OUT2_15_port, OUT2(14) => 
                           RF_OUT2_14_port, OUT2(13) => RF_OUT2_13_port, 
                           OUT2(12) => RF_OUT2_12_port, OUT2(11) => 
                           RF_OUT2_11_port, OUT2(10) => RF_OUT2_10_port, 
                           OUT2(9) => RF_OUT2_9_port, OUT2(8) => RF_OUT2_8_port
                           , OUT2(7) => RF_OUT2_7_port, OUT2(6) => 
                           RF_OUT2_6_port, OUT2(5) => RF_OUT2_5_port, OUT2(4) 
                           => RF_OUT2_4_port, OUT2(3) => RF_OUT2_3_port, 
                           OUT2(2) => RF_OUT2_2_port, OUT2(1) => RF_OUT2_1_port
                           , OUT2(0) => RF_OUT2_0_port);
   SIGN_EXTEND : SIGNEX_N32_OPC6_REG5 port map( INSTR(31) => IF_ID_IR_31_port, 
                           INSTR(30) => IF_ID_IR_30_port, INSTR(29) => 
                           IF_ID_IR_29_port, INSTR(28) => IF_ID_IR_28_port, 
                           INSTR(27) => IF_ID_IR_27_port, INSTR(26) => 
                           IF_ID_IR_26_port, INSTR(25) => IF_ID_IR_25_port, 
                           INSTR(24) => IF_ID_IR_24_port, INSTR(23) => 
                           IF_ID_IR_23_port, INSTR(22) => IF_ID_IR_22_port, 
                           INSTR(21) => IF_ID_IR_21_port, INSTR(20) => 
                           IF_ID_IR_20_port, INSTR(19) => IF_ID_IR_19_port, 
                           INSTR(18) => IF_ID_IR_18_port, INSTR(17) => 
                           IF_ID_IR_17_port, INSTR(16) => IF_ID_IR_16_port, 
                           INSTR(15) => IF_ID_IR_15_port, INSTR(14) => 
                           IF_ID_IR_14_port, INSTR(13) => IF_ID_IR_13_port, 
                           INSTR(12) => IF_ID_IR_12_port, INSTR(11) => 
                           IF_ID_IR_11_port, INSTR(10) => IF_ID_IR_10_port, 
                           INSTR(9) => IF_ID_IR_9_port, INSTR(8) => 
                           IF_ID_IR_8_port, INSTR(7) => IF_ID_IR_7_port, 
                           INSTR(6) => IF_ID_IR_6_port, INSTR(5) => 
                           IF_ID_IR_5_port, INSTR(4) => IF_ID_IR_4_port, 
                           INSTR(3) => IF_ID_IR_3_port, INSTR(2) => 
                           IF_ID_IR_2_port, INSTR(1) => IF_ID_IR_1_port, 
                           INSTR(0) => IF_ID_IR_0_port, IMM(31) => 
                           IMM_OUT_31_port, IMM(30) => IMM_OUT_30_port, IMM(29)
                           => IMM_OUT_29_port, IMM(28) => IMM_OUT_28_port, 
                           IMM(27) => IMM_OUT_27_port, IMM(26) => 
                           IMM_OUT_26_port, IMM(25) => IMM_OUT_25_port, IMM(24)
                           => IMM_OUT_24_port, IMM(23) => IMM_OUT_23_port, 
                           IMM(22) => IMM_OUT_22_port, IMM(21) => 
                           IMM_OUT_21_port, IMM(20) => IMM_OUT_20_port, IMM(19)
                           => IMM_OUT_19_port, IMM(18) => IMM_OUT_18_port, 
                           IMM(17) => IMM_OUT_17_port, IMM(16) => 
                           IMM_OUT_16_port, IMM(15) => IMM_OUT_15_port, IMM(14)
                           => IMM_OUT_14_port, IMM(13) => IMM_OUT_13_port, 
                           IMM(12) => IMM_OUT_12_port, IMM(11) => 
                           IMM_OUT_11_port, IMM(10) => IMM_OUT_10_port, IMM(9) 
                           => IMM_OUT_9_port, IMM(8) => IMM_OUT_8_port, IMM(7) 
                           => IMM_OUT_7_port, IMM(6) => IMM_OUT_6_port, IMM(5) 
                           => IMM_OUT_5_port, IMM(4) => IMM_OUT_4_port, IMM(3) 
                           => IMM_OUT_3_port, IMM(2) => IMM_OUT_2_port, IMM(1) 
                           => IMM_OUT_1_port, IMM(0) => IMM_OUT_0_port);
   REGISTER_ADDRESSER : REGADDR_N32_OPC6_REG5 port map( INSTR(31) => 
                           IF_ID_IR_31_port, INSTR(30) => IF_ID_IR_30_port, 
                           INSTR(29) => IF_ID_IR_29_port, INSTR(28) => 
                           IF_ID_IR_28_port, INSTR(27) => IF_ID_IR_27_port, 
                           INSTR(26) => IF_ID_IR_26_port, INSTR(25) => 
                           IF_ID_IR_25_port, INSTR(24) => IF_ID_IR_24_port, 
                           INSTR(23) => IF_ID_IR_23_port, INSTR(22) => 
                           IF_ID_IR_22_port, INSTR(21) => IF_ID_IR_21_port, 
                           INSTR(20) => IF_ID_IR_20_port, INSTR(19) => 
                           IF_ID_IR_19_port, INSTR(18) => IF_ID_IR_18_port, 
                           INSTR(17) => IF_ID_IR_17_port, INSTR(16) => 
                           IF_ID_IR_16_port, INSTR(15) => IF_ID_IR_15_port, 
                           INSTR(14) => IF_ID_IR_14_port, INSTR(13) => 
                           IF_ID_IR_13_port, INSTR(12) => IF_ID_IR_12_port, 
                           INSTR(11) => IF_ID_IR_11_port, INSTR(10) => 
                           IF_ID_IR_10_port, INSTR(9) => IF_ID_IR_9_port, 
                           INSTR(8) => IF_ID_IR_8_port, INSTR(7) => 
                           IF_ID_IR_7_port, INSTR(6) => IF_ID_IR_6_port, 
                           INSTR(5) => IF_ID_IR_5_port, INSTR(4) => 
                           IF_ID_IR_4_port, INSTR(3) => IF_ID_IR_3_port, 
                           INSTR(2) => IF_ID_IR_2_port, INSTR(1) => 
                           IF_ID_IR_1_port, INSTR(0) => IF_ID_IR_0_port, RS1(4)
                           => ID_EX_RS1_NEXT_4_port, RS1(3) => 
                           ID_EX_RS1_NEXT_3_port, RS1(2) => 
                           ID_EX_RS1_NEXT_2_port, RS1(1) => 
                           ID_EX_RS1_NEXT_1_port, RS1(0) => 
                           ID_EX_RS1_NEXT_0_port, RS2(4) => 
                           ID_EX_RS2_NEXT_4_port, RS2(3) => 
                           ID_EX_RS2_NEXT_3_port, RS2(2) => 
                           ID_EX_RS2_NEXT_2_port, RS2(1) => 
                           ID_EX_RS2_NEXT_1_port, RS2(0) => 
                           ID_EX_RS2_NEXT_0_port, RD(4) => ID_EX_RD_NEXT_4_port
                           , RD(3) => ID_EX_RD_NEXT_3_port, RD(2) => 
                           ID_EX_RD_NEXT_2_port, RD(1) => ID_EX_RD_NEXT_1_port,
                           RD(0) => ID_EX_RD_NEXT_0_port);
   LATCH_RF1 : LDR_N32_4 port map( RST => RST, EN => RegA_LATCH_EN, REGIN(31) 
                           => RF_OUT1_31_port, REGIN(30) => RF_OUT1_30_port, 
                           REGIN(29) => RF_OUT1_29_port, REGIN(28) => 
                           RF_OUT1_28_port, REGIN(27) => RF_OUT1_27_port, 
                           REGIN(26) => RF_OUT1_26_port, REGIN(25) => 
                           RF_OUT1_25_port, REGIN(24) => RF_OUT1_24_port, 
                           REGIN(23) => RF_OUT1_23_port, REGIN(22) => 
                           RF_OUT1_22_port, REGIN(21) => RF_OUT1_21_port, 
                           REGIN(20) => RF_OUT1_20_port, REGIN(19) => 
                           RF_OUT1_19_port, REGIN(18) => RF_OUT1_18_port, 
                           REGIN(17) => RF_OUT1_17_port, REGIN(16) => 
                           RF_OUT1_16_port, REGIN(15) => RF_OUT1_15_port, 
                           REGIN(14) => RF_OUT1_14_port, REGIN(13) => 
                           RF_OUT1_13_port, REGIN(12) => RF_OUT1_12_port, 
                           REGIN(11) => RF_OUT1_11_port, REGIN(10) => 
                           RF_OUT1_10_port, REGIN(9) => RF_OUT1_9_port, 
                           REGIN(8) => RF_OUT1_8_port, REGIN(7) => 
                           RF_OUT1_7_port, REGIN(6) => RF_OUT1_6_port, REGIN(5)
                           => RF_OUT1_5_port, REGIN(4) => RF_OUT1_4_port, 
                           REGIN(3) => RF_OUT1_3_port, REGIN(2) => 
                           RF_OUT1_2_port, REGIN(1) => RF_OUT1_1_port, REGIN(0)
                           => RF_OUT1_0_port, REGOUT(31) => 
                           ID_EX_RF_OUT1_NEXT_31_port, REGOUT(30) => 
                           ID_EX_RF_OUT1_NEXT_30_port, REGOUT(29) => 
                           ID_EX_RF_OUT1_NEXT_29_port, REGOUT(28) => 
                           ID_EX_RF_OUT1_NEXT_28_port, REGOUT(27) => 
                           ID_EX_RF_OUT1_NEXT_27_port, REGOUT(26) => 
                           ID_EX_RF_OUT1_NEXT_26_port, REGOUT(25) => 
                           ID_EX_RF_OUT1_NEXT_25_port, REGOUT(24) => 
                           ID_EX_RF_OUT1_NEXT_24_port, REGOUT(23) => 
                           ID_EX_RF_OUT1_NEXT_23_port, REGOUT(22) => 
                           ID_EX_RF_OUT1_NEXT_22_port, REGOUT(21) => 
                           ID_EX_RF_OUT1_NEXT_21_port, REGOUT(20) => 
                           ID_EX_RF_OUT1_NEXT_20_port, REGOUT(19) => 
                           ID_EX_RF_OUT1_NEXT_19_port, REGOUT(18) => 
                           ID_EX_RF_OUT1_NEXT_18_port, REGOUT(17) => 
                           ID_EX_RF_OUT1_NEXT_17_port, REGOUT(16) => 
                           ID_EX_RF_OUT1_NEXT_16_port, REGOUT(15) => 
                           ID_EX_RF_OUT1_NEXT_15_port, REGOUT(14) => 
                           ID_EX_RF_OUT1_NEXT_14_port, REGOUT(13) => 
                           ID_EX_RF_OUT1_NEXT_13_port, REGOUT(12) => 
                           ID_EX_RF_OUT1_NEXT_12_port, REGOUT(11) => 
                           ID_EX_RF_OUT1_NEXT_11_port, REGOUT(10) => 
                           ID_EX_RF_OUT1_NEXT_10_port, REGOUT(9) => 
                           ID_EX_RF_OUT1_NEXT_9_port, REGOUT(8) => 
                           ID_EX_RF_OUT1_NEXT_8_port, REGOUT(7) => 
                           ID_EX_RF_OUT1_NEXT_7_port, REGOUT(6) => 
                           ID_EX_RF_OUT1_NEXT_6_port, REGOUT(5) => 
                           ID_EX_RF_OUT1_NEXT_5_port, REGOUT(4) => 
                           ID_EX_RF_OUT1_NEXT_4_port, REGOUT(3) => 
                           ID_EX_RF_OUT1_NEXT_3_port, REGOUT(2) => 
                           ID_EX_RF_OUT1_NEXT_2_port, REGOUT(1) => 
                           ID_EX_RF_OUT1_NEXT_1_port, REGOUT(0) => 
                           ID_EX_RF_OUT1_NEXT_0_port);
   LATCH_RF2 : LDR_N32_3 port map( RST => RST, EN => RegB_LATCH_EN, REGIN(31) 
                           => RF_OUT2_31_port, REGIN(30) => RF_OUT2_30_port, 
                           REGIN(29) => RF_OUT2_29_port, REGIN(28) => 
                           RF_OUT2_28_port, REGIN(27) => RF_OUT2_27_port, 
                           REGIN(26) => RF_OUT2_26_port, REGIN(25) => 
                           RF_OUT2_25_port, REGIN(24) => RF_OUT2_24_port, 
                           REGIN(23) => RF_OUT2_23_port, REGIN(22) => 
                           RF_OUT2_22_port, REGIN(21) => RF_OUT2_21_port, 
                           REGIN(20) => RF_OUT2_20_port, REGIN(19) => 
                           RF_OUT2_19_port, REGIN(18) => RF_OUT2_18_port, 
                           REGIN(17) => RF_OUT2_17_port, REGIN(16) => 
                           RF_OUT2_16_port, REGIN(15) => RF_OUT2_15_port, 
                           REGIN(14) => RF_OUT2_14_port, REGIN(13) => 
                           RF_OUT2_13_port, REGIN(12) => RF_OUT2_12_port, 
                           REGIN(11) => RF_OUT2_11_port, REGIN(10) => 
                           RF_OUT2_10_port, REGIN(9) => RF_OUT2_9_port, 
                           REGIN(8) => RF_OUT2_8_port, REGIN(7) => 
                           RF_OUT2_7_port, REGIN(6) => RF_OUT2_6_port, REGIN(5)
                           => RF_OUT2_5_port, REGIN(4) => RF_OUT2_4_port, 
                           REGIN(3) => RF_OUT2_3_port, REGIN(2) => 
                           RF_OUT2_2_port, REGIN(1) => RF_OUT2_1_port, REGIN(0)
                           => RF_OUT2_0_port, REGOUT(31) => 
                           ID_EX_RF_OUT2_NEXT_31_port, REGOUT(30) => 
                           ID_EX_RF_OUT2_NEXT_30_port, REGOUT(29) => 
                           ID_EX_RF_OUT2_NEXT_29_port, REGOUT(28) => 
                           ID_EX_RF_OUT2_NEXT_28_port, REGOUT(27) => 
                           ID_EX_RF_OUT2_NEXT_27_port, REGOUT(26) => 
                           ID_EX_RF_OUT2_NEXT_26_port, REGOUT(25) => 
                           ID_EX_RF_OUT2_NEXT_25_port, REGOUT(24) => 
                           ID_EX_RF_OUT2_NEXT_24_port, REGOUT(23) => 
                           ID_EX_RF_OUT2_NEXT_23_port, REGOUT(22) => 
                           ID_EX_RF_OUT2_NEXT_22_port, REGOUT(21) => 
                           ID_EX_RF_OUT2_NEXT_21_port, REGOUT(20) => 
                           ID_EX_RF_OUT2_NEXT_20_port, REGOUT(19) => 
                           ID_EX_RF_OUT2_NEXT_19_port, REGOUT(18) => 
                           ID_EX_RF_OUT2_NEXT_18_port, REGOUT(17) => 
                           ID_EX_RF_OUT2_NEXT_17_port, REGOUT(16) => 
                           ID_EX_RF_OUT2_NEXT_16_port, REGOUT(15) => 
                           ID_EX_RF_OUT2_NEXT_15_port, REGOUT(14) => 
                           ID_EX_RF_OUT2_NEXT_14_port, REGOUT(13) => 
                           ID_EX_RF_OUT2_NEXT_13_port, REGOUT(12) => 
                           ID_EX_RF_OUT2_NEXT_12_port, REGOUT(11) => 
                           ID_EX_RF_OUT2_NEXT_11_port, REGOUT(10) => 
                           ID_EX_RF_OUT2_NEXT_10_port, REGOUT(9) => 
                           ID_EX_RF_OUT2_NEXT_9_port, REGOUT(8) => 
                           ID_EX_RF_OUT2_NEXT_8_port, REGOUT(7) => 
                           ID_EX_RF_OUT2_NEXT_7_port, REGOUT(6) => 
                           ID_EX_RF_OUT2_NEXT_6_port, REGOUT(5) => 
                           ID_EX_RF_OUT2_NEXT_5_port, REGOUT(4) => 
                           ID_EX_RF_OUT2_NEXT_4_port, REGOUT(3) => 
                           ID_EX_RF_OUT2_NEXT_3_port, REGOUT(2) => 
                           ID_EX_RF_OUT2_NEXT_2_port, REGOUT(1) => 
                           ID_EX_RF_OUT2_NEXT_1_port, REGOUT(0) => 
                           ID_EX_RF_OUT2_NEXT_0_port);
   LATCH_IMM : LDR_N32_2 port map( RST => RST, EN => RegIMM_LATCH_EN, REGIN(31)
                           => IMM_OUT_31_port, REGIN(30) => IMM_OUT_30_port, 
                           REGIN(29) => IMM_OUT_29_port, REGIN(28) => 
                           IMM_OUT_28_port, REGIN(27) => IMM_OUT_27_port, 
                           REGIN(26) => IMM_OUT_26_port, REGIN(25) => 
                           IMM_OUT_25_port, REGIN(24) => IMM_OUT_24_port, 
                           REGIN(23) => IMM_OUT_23_port, REGIN(22) => 
                           IMM_OUT_22_port, REGIN(21) => IMM_OUT_21_port, 
                           REGIN(20) => IMM_OUT_20_port, REGIN(19) => 
                           IMM_OUT_19_port, REGIN(18) => IMM_OUT_18_port, 
                           REGIN(17) => IMM_OUT_17_port, REGIN(16) => 
                           IMM_OUT_16_port, REGIN(15) => IMM_OUT_15_port, 
                           REGIN(14) => IMM_OUT_14_port, REGIN(13) => 
                           IMM_OUT_13_port, REGIN(12) => IMM_OUT_12_port, 
                           REGIN(11) => IMM_OUT_11_port, REGIN(10) => 
                           IMM_OUT_10_port, REGIN(9) => IMM_OUT_9_port, 
                           REGIN(8) => IMM_OUT_8_port, REGIN(7) => 
                           IMM_OUT_7_port, REGIN(6) => IMM_OUT_6_port, REGIN(5)
                           => IMM_OUT_5_port, REGIN(4) => IMM_OUT_4_port, 
                           REGIN(3) => IMM_OUT_3_port, REGIN(2) => 
                           IMM_OUT_2_port, REGIN(1) => IMM_OUT_1_port, REGIN(0)
                           => IMM_OUT_0_port, REGOUT(31) => 
                           ID_EX_IMM_NEXT_31_port, REGOUT(30) => 
                           ID_EX_IMM_NEXT_30_port, REGOUT(29) => 
                           ID_EX_IMM_NEXT_29_port, REGOUT(28) => 
                           ID_EX_IMM_NEXT_28_port, REGOUT(27) => 
                           ID_EX_IMM_NEXT_27_port, REGOUT(26) => 
                           ID_EX_IMM_NEXT_26_port, REGOUT(25) => 
                           ID_EX_IMM_NEXT_25_port, REGOUT(24) => 
                           ID_EX_IMM_NEXT_24_port, REGOUT(23) => 
                           ID_EX_IMM_NEXT_23_port, REGOUT(22) => 
                           ID_EX_IMM_NEXT_22_port, REGOUT(21) => 
                           ID_EX_IMM_NEXT_21_port, REGOUT(20) => 
                           ID_EX_IMM_NEXT_20_port, REGOUT(19) => 
                           ID_EX_IMM_NEXT_19_port, REGOUT(18) => 
                           ID_EX_IMM_NEXT_18_port, REGOUT(17) => 
                           ID_EX_IMM_NEXT_17_port, REGOUT(16) => 
                           ID_EX_IMM_NEXT_16_port, REGOUT(15) => 
                           ID_EX_IMM_NEXT_15_port, REGOUT(14) => 
                           ID_EX_IMM_NEXT_14_port, REGOUT(13) => 
                           ID_EX_IMM_NEXT_13_port, REGOUT(12) => 
                           ID_EX_IMM_NEXT_12_port, REGOUT(11) => 
                           ID_EX_IMM_NEXT_11_port, REGOUT(10) => 
                           ID_EX_IMM_NEXT_10_port, REGOUT(9) => 
                           ID_EX_IMM_NEXT_9_port, REGOUT(8) => 
                           ID_EX_IMM_NEXT_8_port, REGOUT(7) => 
                           ID_EX_IMM_NEXT_7_port, REGOUT(6) => 
                           ID_EX_IMM_NEXT_6_port, REGOUT(5) => 
                           ID_EX_IMM_NEXT_5_port, REGOUT(4) => 
                           ID_EX_IMM_NEXT_4_port, REGOUT(3) => 
                           ID_EX_IMM_NEXT_3_port, REGOUT(2) => 
                           ID_EX_IMM_NEXT_2_port, REGOUT(1) => 
                           ID_EX_IMM_NEXT_1_port, REGOUT(0) => 
                           ID_EX_IMM_NEXT_0_port);
   ALU_PRE_MUX1 : MUX41_N32_1 port map( A(31) => ID_EX_RF_OUT1_31_port, A(30) 
                           => ID_EX_RF_OUT1_30_port, A(29) => 
                           ID_EX_RF_OUT1_29_port, A(28) => 
                           ID_EX_RF_OUT1_28_port, A(27) => 
                           ID_EX_RF_OUT1_27_port, A(26) => 
                           ID_EX_RF_OUT1_26_port, A(25) => 
                           ID_EX_RF_OUT1_25_port, A(24) => 
                           ID_EX_RF_OUT1_24_port, A(23) => 
                           ID_EX_RF_OUT1_23_port, A(22) => 
                           ID_EX_RF_OUT1_22_port, A(21) => 
                           ID_EX_RF_OUT1_21_port, A(20) => 
                           ID_EX_RF_OUT1_20_port, A(19) => 
                           ID_EX_RF_OUT1_19_port, A(18) => 
                           ID_EX_RF_OUT1_18_port, A(17) => 
                           ID_EX_RF_OUT1_17_port, A(16) => 
                           ID_EX_RF_OUT1_16_port, A(15) => 
                           ID_EX_RF_OUT1_15_port, A(14) => 
                           ID_EX_RF_OUT1_14_port, A(13) => 
                           ID_EX_RF_OUT1_13_port, A(12) => 
                           ID_EX_RF_OUT1_12_port, A(11) => 
                           ID_EX_RF_OUT1_11_port, A(10) => 
                           ID_EX_RF_OUT1_10_port, A(9) => ID_EX_RF_OUT1_9_port,
                           A(8) => ID_EX_RF_OUT1_8_port, A(7) => 
                           ID_EX_RF_OUT1_7_port, A(6) => ID_EX_RF_OUT1_6_port, 
                           A(5) => ID_EX_RF_OUT1_5_port, A(4) => 
                           ID_EX_RF_OUT1_4_port, A(3) => ID_EX_RF_OUT1_3_port, 
                           A(2) => ID_EX_RF_OUT1_2_port, A(1) => 
                           ID_EX_RF_OUT1_1_port, A(0) => ID_EX_RF_OUT1_0_port, 
                           B(31) => ALU_OUT_31_port, B(30) => ALU_OUT_30_port, 
                           B(29) => ALU_OUT_29_port, B(28) => ALU_OUT_28_port, 
                           B(27) => ALU_OUT_27_port, B(26) => ALU_OUT_26_port, 
                           B(25) => ALU_OUT_25_port, B(24) => ALU_OUT_24_port, 
                           B(23) => ALU_OUT_23_port, B(22) => ALU_OUT_22_port, 
                           B(21) => ALU_OUT_21_port, B(20) => ALU_OUT_20_port, 
                           B(19) => ALU_OUT_19_port, B(18) => ALU_OUT_18_port, 
                           B(17) => ALU_OUT_17_port, B(16) => ALU_OUT_16_port, 
                           B(15) => ALU_OUT_15_port, B(14) => ALU_OUT_14_port, 
                           B(13) => ALU_OUT_13_port, B(12) => ALU_OUT_12_port, 
                           B(11) => ALU_OUT_11_port, B(10) => ALU_OUT_10_port, 
                           B(9) => ALU_OUT_9_port, B(8) => ALU_OUT_8_port, B(7)
                           => ALU_OUT_7_port, B(6) => ALU_OUT_6_port, B(5) => 
                           ALU_OUT_5_port, B(4) => ALU_OUT_4_port, B(3) => 
                           ALU_OUT_3_port, B(2) => ALU_OUT_2_port, B(1) => 
                           ALU_OUT_1_port, B(0) => ALU_OUT_0_port, C(31) => 
                           JAL_MUX_OUT_31_port, C(30) => JAL_MUX_OUT_30_port, 
                           C(29) => JAL_MUX_OUT_29_port, C(28) => 
                           JAL_MUX_OUT_28_port, C(27) => JAL_MUX_OUT_27_port, 
                           C(26) => JAL_MUX_OUT_26_port, C(25) => 
                           JAL_MUX_OUT_25_port, C(24) => JAL_MUX_OUT_24_port, 
                           C(23) => JAL_MUX_OUT_23_port, C(22) => 
                           JAL_MUX_OUT_22_port, C(21) => JAL_MUX_OUT_21_port, 
                           C(20) => JAL_MUX_OUT_20_port, C(19) => 
                           JAL_MUX_OUT_19_port, C(18) => JAL_MUX_OUT_18_port, 
                           C(17) => JAL_MUX_OUT_17_port, C(16) => 
                           JAL_MUX_OUT_16_port, C(15) => JAL_MUX_OUT_15_port, 
                           C(14) => JAL_MUX_OUT_14_port, C(13) => 
                           JAL_MUX_OUT_13_port, C(12) => JAL_MUX_OUT_12_port, 
                           C(11) => JAL_MUX_OUT_11_port, C(10) => 
                           JAL_MUX_OUT_10_port, C(9) => JAL_MUX_OUT_9_port, 
                           C(8) => JAL_MUX_OUT_8_port, C(7) => 
                           JAL_MUX_OUT_7_port, C(6) => JAL_MUX_OUT_6_port, C(5)
                           => JAL_MUX_OUT_5_port, C(4) => JAL_MUX_OUT_4_port, 
                           C(3) => JAL_MUX_OUT_3_port, C(2) => 
                           JAL_MUX_OUT_2_port, C(1) => JAL_MUX_OUT_1_port, C(0)
                           => JAL_MUX_OUT_0_port, D(31) => X_Logic0_port, D(30)
                           => X_Logic0_port, D(29) => X_Logic0_port, D(28) => 
                           X_Logic0_port, D(27) => X_Logic0_port, D(26) => 
                           X_Logic0_port, D(25) => X_Logic0_port, D(24) => 
                           X_Logic0_port, D(23) => X_Logic0_port, D(22) => 
                           X_Logic0_port, D(21) => X_Logic0_port, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, S(1) => FORWARD_A_1_port, S(0) => 
                           FORWARD_A_0_port, Y(31) => ALU_PREOP1_31_port, Y(30)
                           => ALU_PREOP1_30_port, Y(29) => ALU_PREOP1_29_port, 
                           Y(28) => ALU_PREOP1_28_port, Y(27) => 
                           ALU_PREOP1_27_port, Y(26) => ALU_PREOP1_26_port, 
                           Y(25) => ALU_PREOP1_25_port, Y(24) => 
                           ALU_PREOP1_24_port, Y(23) => ALU_PREOP1_23_port, 
                           Y(22) => ALU_PREOP1_22_port, Y(21) => 
                           ALU_PREOP1_21_port, Y(20) => ALU_PREOP1_20_port, 
                           Y(19) => ALU_PREOP1_19_port, Y(18) => 
                           ALU_PREOP1_18_port, Y(17) => ALU_PREOP1_17_port, 
                           Y(16) => ALU_PREOP1_16_port, Y(15) => 
                           ALU_PREOP1_15_port, Y(14) => ALU_PREOP1_14_port, 
                           Y(13) => ALU_PREOP1_13_port, Y(12) => 
                           ALU_PREOP1_12_port, Y(11) => ALU_PREOP1_11_port, 
                           Y(10) => ALU_PREOP1_10_port, Y(9) => 
                           ALU_PREOP1_9_port, Y(8) => ALU_PREOP1_8_port, Y(7) 
                           => ALU_PREOP1_7_port, Y(6) => ALU_PREOP1_6_port, 
                           Y(5) => ALU_PREOP1_5_port, Y(4) => ALU_PREOP1_4_port
                           , Y(3) => ALU_PREOP1_3_port, Y(2) => 
                           ALU_PREOP1_2_port, Y(1) => ALU_PREOP1_1_port, Y(0) 
                           => ALU_PREOP1_0_port);
   ALU_PRE_MUX2 : MUX41_N32_0 port map( A(31) => ID_EX_RF_OUT2_31_port, A(30) 
                           => ID_EX_RF_OUT2_30_port, A(29) => 
                           ID_EX_RF_OUT2_29_port, A(28) => 
                           ID_EX_RF_OUT2_28_port, A(27) => 
                           ID_EX_RF_OUT2_27_port, A(26) => 
                           ID_EX_RF_OUT2_26_port, A(25) => 
                           ID_EX_RF_OUT2_25_port, A(24) => 
                           ID_EX_RF_OUT2_24_port, A(23) => 
                           ID_EX_RF_OUT2_23_port, A(22) => 
                           ID_EX_RF_OUT2_22_port, A(21) => 
                           ID_EX_RF_OUT2_21_port, A(20) => 
                           ID_EX_RF_OUT2_20_port, A(19) => 
                           ID_EX_RF_OUT2_19_port, A(18) => 
                           ID_EX_RF_OUT2_18_port, A(17) => 
                           ID_EX_RF_OUT2_17_port, A(16) => 
                           ID_EX_RF_OUT2_16_port, A(15) => 
                           ID_EX_RF_OUT2_15_port, A(14) => 
                           ID_EX_RF_OUT2_14_port, A(13) => 
                           ID_EX_RF_OUT2_13_port, A(12) => 
                           ID_EX_RF_OUT2_12_port, A(11) => 
                           ID_EX_RF_OUT2_11_port, A(10) => 
                           ID_EX_RF_OUT2_10_port, A(9) => ID_EX_RF_OUT2_9_port,
                           A(8) => ID_EX_RF_OUT2_8_port, A(7) => 
                           ID_EX_RF_OUT2_7_port, A(6) => ID_EX_RF_OUT2_6_port, 
                           A(5) => ID_EX_RF_OUT2_5_port, A(4) => 
                           ID_EX_RF_OUT2_4_port, A(3) => ID_EX_RF_OUT2_3_port, 
                           A(2) => ID_EX_RF_OUT2_2_port, A(1) => 
                           ID_EX_RF_OUT2_1_port, A(0) => ID_EX_RF_OUT2_0_port, 
                           B(31) => ALU_OUT_31_port, B(30) => ALU_OUT_30_port, 
                           B(29) => ALU_OUT_29_port, B(28) => ALU_OUT_28_port, 
                           B(27) => ALU_OUT_27_port, B(26) => ALU_OUT_26_port, 
                           B(25) => ALU_OUT_25_port, B(24) => ALU_OUT_24_port, 
                           B(23) => ALU_OUT_23_port, B(22) => ALU_OUT_22_port, 
                           B(21) => ALU_OUT_21_port, B(20) => ALU_OUT_20_port, 
                           B(19) => ALU_OUT_19_port, B(18) => ALU_OUT_18_port, 
                           B(17) => ALU_OUT_17_port, B(16) => ALU_OUT_16_port, 
                           B(15) => ALU_OUT_15_port, B(14) => ALU_OUT_14_port, 
                           B(13) => ALU_OUT_13_port, B(12) => ALU_OUT_12_port, 
                           B(11) => ALU_OUT_11_port, B(10) => ALU_OUT_10_port, 
                           B(9) => ALU_OUT_9_port, B(8) => ALU_OUT_8_port, B(7)
                           => ALU_OUT_7_port, B(6) => ALU_OUT_6_port, B(5) => 
                           ALU_OUT_5_port, B(4) => ALU_OUT_4_port, B(3) => 
                           ALU_OUT_3_port, B(2) => ALU_OUT_2_port, B(1) => 
                           ALU_OUT_1_port, B(0) => ALU_OUT_0_port, C(31) => 
                           JAL_MUX_OUT_31_port, C(30) => JAL_MUX_OUT_30_port, 
                           C(29) => JAL_MUX_OUT_29_port, C(28) => 
                           JAL_MUX_OUT_28_port, C(27) => JAL_MUX_OUT_27_port, 
                           C(26) => JAL_MUX_OUT_26_port, C(25) => 
                           JAL_MUX_OUT_25_port, C(24) => JAL_MUX_OUT_24_port, 
                           C(23) => JAL_MUX_OUT_23_port, C(22) => 
                           JAL_MUX_OUT_22_port, C(21) => JAL_MUX_OUT_21_port, 
                           C(20) => JAL_MUX_OUT_20_port, C(19) => 
                           JAL_MUX_OUT_19_port, C(18) => JAL_MUX_OUT_18_port, 
                           C(17) => JAL_MUX_OUT_17_port, C(16) => 
                           JAL_MUX_OUT_16_port, C(15) => JAL_MUX_OUT_15_port, 
                           C(14) => JAL_MUX_OUT_14_port, C(13) => 
                           JAL_MUX_OUT_13_port, C(12) => JAL_MUX_OUT_12_port, 
                           C(11) => JAL_MUX_OUT_11_port, C(10) => 
                           JAL_MUX_OUT_10_port, C(9) => JAL_MUX_OUT_9_port, 
                           C(8) => JAL_MUX_OUT_8_port, C(7) => 
                           JAL_MUX_OUT_7_port, C(6) => JAL_MUX_OUT_6_port, C(5)
                           => JAL_MUX_OUT_5_port, C(4) => JAL_MUX_OUT_4_port, 
                           C(3) => JAL_MUX_OUT_3_port, C(2) => 
                           JAL_MUX_OUT_2_port, C(1) => JAL_MUX_OUT_1_port, C(0)
                           => JAL_MUX_OUT_0_port, D(31) => X_Logic0_port, D(30)
                           => X_Logic0_port, D(29) => X_Logic0_port, D(28) => 
                           X_Logic0_port, D(27) => X_Logic0_port, D(26) => 
                           X_Logic0_port, D(25) => X_Logic0_port, D(24) => 
                           X_Logic0_port, D(23) => X_Logic0_port, D(22) => 
                           X_Logic0_port, D(21) => X_Logic0_port, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, S(1) => FORWARD_B_1_port, S(0) => 
                           FORWARD_B_0_port, Y(31) => ALU_PREOP2_31_port, Y(30)
                           => ALU_PREOP2_30_port, Y(29) => ALU_PREOP2_29_port, 
                           Y(28) => ALU_PREOP2_28_port, Y(27) => 
                           ALU_PREOP2_27_port, Y(26) => ALU_PREOP2_26_port, 
                           Y(25) => ALU_PREOP2_25_port, Y(24) => 
                           ALU_PREOP2_24_port, Y(23) => ALU_PREOP2_23_port, 
                           Y(22) => ALU_PREOP2_22_port, Y(21) => 
                           ALU_PREOP2_21_port, Y(20) => ALU_PREOP2_20_port, 
                           Y(19) => ALU_PREOP2_19_port, Y(18) => 
                           ALU_PREOP2_18_port, Y(17) => ALU_PREOP2_17_port, 
                           Y(16) => ALU_PREOP2_16_port, Y(15) => 
                           ALU_PREOP2_15_port, Y(14) => ALU_PREOP2_14_port, 
                           Y(13) => ALU_PREOP2_13_port, Y(12) => 
                           ALU_PREOP2_12_port, Y(11) => ALU_PREOP2_11_port, 
                           Y(10) => ALU_PREOP2_10_port, Y(9) => 
                           ALU_PREOP2_9_port, Y(8) => ALU_PREOP2_8_port, Y(7) 
                           => ALU_PREOP2_7_port, Y(6) => ALU_PREOP2_6_port, 
                           Y(5) => ALU_PREOP2_5_port, Y(4) => ALU_PREOP2_4_port
                           , Y(3) => ALU_PREOP2_3_port, Y(2) => 
                           ALU_PREOP2_2_port, Y(1) => ALU_PREOP2_1_port, Y(0) 
                           => ALU_PREOP2_0_port);
   ALU_MUX1 : MUX21_N32_3 port map( A(31) => ALU_PREOP1_31_port, A(30) => 
                           ALU_PREOP1_30_port, A(29) => ALU_PREOP1_29_port, 
                           A(28) => ALU_PREOP1_28_port, A(27) => 
                           ALU_PREOP1_27_port, A(26) => ALU_PREOP1_26_port, 
                           A(25) => ALU_PREOP1_25_port, A(24) => 
                           ALU_PREOP1_24_port, A(23) => ALU_PREOP1_23_port, 
                           A(22) => ALU_PREOP1_22_port, A(21) => 
                           ALU_PREOP1_21_port, A(20) => ALU_PREOP1_20_port, 
                           A(19) => ALU_PREOP1_19_port, A(18) => 
                           ALU_PREOP1_18_port, A(17) => ALU_PREOP1_17_port, 
                           A(16) => ALU_PREOP1_16_port, A(15) => 
                           ALU_PREOP1_15_port, A(14) => ALU_PREOP1_14_port, 
                           A(13) => ALU_PREOP1_13_port, A(12) => 
                           ALU_PREOP1_12_port, A(11) => ALU_PREOP1_11_port, 
                           A(10) => ALU_PREOP1_10_port, A(9) => 
                           ALU_PREOP1_9_port, A(8) => ALU_PREOP1_8_port, A(7) 
                           => ALU_PREOP1_7_port, A(6) => ALU_PREOP1_6_port, 
                           A(5) => ALU_PREOP1_5_port, A(4) => ALU_PREOP1_4_port
                           , A(3) => ALU_PREOP1_3_port, A(2) => 
                           ALU_PREOP1_2_port, A(1) => ALU_PREOP1_1_port, A(0) 
                           => ALU_PREOP1_0_port, B(31) => ID_EX_NPC_31_port, 
                           B(30) => ID_EX_NPC_30_port, B(29) => 
                           ID_EX_NPC_29_port, B(28) => ID_EX_NPC_28_port, B(27)
                           => ID_EX_NPC_27_port, B(26) => ID_EX_NPC_26_port, 
                           B(25) => ID_EX_NPC_25_port, B(24) => 
                           ID_EX_NPC_24_port, B(23) => ID_EX_NPC_23_port, B(22)
                           => ID_EX_NPC_22_port, B(21) => ID_EX_NPC_21_port, 
                           B(20) => ID_EX_NPC_20_port, B(19) => 
                           ID_EX_NPC_19_port, B(18) => ID_EX_NPC_18_port, B(17)
                           => ID_EX_NPC_17_port, B(16) => ID_EX_NPC_16_port, 
                           B(15) => ID_EX_NPC_15_port, B(14) => 
                           ID_EX_NPC_14_port, B(13) => ID_EX_NPC_13_port, B(12)
                           => ID_EX_NPC_12_port, B(11) => ID_EX_NPC_11_port, 
                           B(10) => ID_EX_NPC_10_port, B(9) => ID_EX_NPC_9_port
                           , B(8) => ID_EX_NPC_8_port, B(7) => ID_EX_NPC_7_port
                           , B(6) => ID_EX_NPC_6_port, B(5) => ID_EX_NPC_5_port
                           , B(4) => ID_EX_NPC_4_port, B(3) => ID_EX_NPC_3_port
                           , B(2) => ID_EX_NPC_2_port, B(1) => ID_EX_NPC_1_port
                           , B(0) => ID_EX_NPC_0_port, S => MUXA_SEL, Y(31) => 
                           ALU_OP1_31_port, Y(30) => ALU_OP1_30_port, Y(29) => 
                           ALU_OP1_29_port, Y(28) => ALU_OP1_28_port, Y(27) => 
                           ALU_OP1_27_port, Y(26) => ALU_OP1_26_port, Y(25) => 
                           ALU_OP1_25_port, Y(24) => ALU_OP1_24_port, Y(23) => 
                           ALU_OP1_23_port, Y(22) => ALU_OP1_22_port, Y(21) => 
                           ALU_OP1_21_port, Y(20) => ALU_OP1_20_port, Y(19) => 
                           ALU_OP1_19_port, Y(18) => ALU_OP1_18_port, Y(17) => 
                           ALU_OP1_17_port, Y(16) => ALU_OP1_16_port, Y(15) => 
                           ALU_OP1_15_port, Y(14) => ALU_OP1_14_port, Y(13) => 
                           ALU_OP1_13_port, Y(12) => ALU_OP1_12_port, Y(11) => 
                           ALU_OP1_11_port, Y(10) => ALU_OP1_10_port, Y(9) => 
                           ALU_OP1_9_port, Y(8) => ALU_OP1_8_port, Y(7) => 
                           ALU_OP1_7_port, Y(6) => ALU_OP1_6_port, Y(5) => 
                           ALU_OP1_5_port, Y(4) => ALU_OP1_4_port, Y(3) => 
                           ALU_OP1_3_port, Y(2) => ALU_OP1_2_port, Y(1) => 
                           ALU_OP1_1_port, Y(0) => ALU_OP1_0_port);
   ALU_MUX2 : MUX21_N32_2 port map( A(31) => ALU_PREOP2_31_port, A(30) => 
                           ALU_PREOP2_30_port, A(29) => ALU_PREOP2_29_port, 
                           A(28) => ALU_PREOP2_28_port, A(27) => 
                           ALU_PREOP2_27_port, A(26) => ALU_PREOP2_26_port, 
                           A(25) => ALU_PREOP2_25_port, A(24) => 
                           ALU_PREOP2_24_port, A(23) => ALU_PREOP2_23_port, 
                           A(22) => ALU_PREOP2_22_port, A(21) => 
                           ALU_PREOP2_21_port, A(20) => ALU_PREOP2_20_port, 
                           A(19) => ALU_PREOP2_19_port, A(18) => 
                           ALU_PREOP2_18_port, A(17) => ALU_PREOP2_17_port, 
                           A(16) => ALU_PREOP2_16_port, A(15) => 
                           ALU_PREOP2_15_port, A(14) => ALU_PREOP2_14_port, 
                           A(13) => ALU_PREOP2_13_port, A(12) => 
                           ALU_PREOP2_12_port, A(11) => ALU_PREOP2_11_port, 
                           A(10) => ALU_PREOP2_10_port, A(9) => 
                           ALU_PREOP2_9_port, A(8) => ALU_PREOP2_8_port, A(7) 
                           => ALU_PREOP2_7_port, A(6) => ALU_PREOP2_6_port, 
                           A(5) => ALU_PREOP2_5_port, A(4) => ALU_PREOP2_4_port
                           , A(3) => ALU_PREOP2_3_port, A(2) => 
                           ALU_PREOP2_2_port, A(1) => ALU_PREOP2_1_port, A(0) 
                           => ALU_PREOP2_0_port, B(31) => ID_EX_IMM_31_port, 
                           B(30) => ID_EX_IMM_30_port, B(29) => 
                           ID_EX_IMM_29_port, B(28) => ID_EX_IMM_28_port, B(27)
                           => ID_EX_IMM_27_port, B(26) => ID_EX_IMM_26_port, 
                           B(25) => ID_EX_IMM_25_port, B(24) => 
                           ID_EX_IMM_24_port, B(23) => ID_EX_IMM_23_port, B(22)
                           => ID_EX_IMM_22_port, B(21) => ID_EX_IMM_21_port, 
                           B(20) => ID_EX_IMM_20_port, B(19) => 
                           ID_EX_IMM_19_port, B(18) => ID_EX_IMM_18_port, B(17)
                           => ID_EX_IMM_17_port, B(16) => ID_EX_IMM_16_port, 
                           B(15) => ID_EX_IMM_15_port, B(14) => 
                           ID_EX_IMM_14_port, B(13) => ID_EX_IMM_13_port, B(12)
                           => ID_EX_IMM_12_port, B(11) => ID_EX_IMM_11_port, 
                           B(10) => ID_EX_IMM_10_port, B(9) => ID_EX_IMM_9_port
                           , B(8) => ID_EX_IMM_8_port, B(7) => ID_EX_IMM_7_port
                           , B(6) => ID_EX_IMM_6_port, B(5) => ID_EX_IMM_5_port
                           , B(4) => ID_EX_IMM_4_port, B(3) => ID_EX_IMM_3_port
                           , B(2) => ID_EX_IMM_2_port, B(1) => ID_EX_IMM_1_port
                           , B(0) => ID_EX_IMM_0_port, S => MUXB_SEL, Y(31) => 
                           ALU_OP2_31_port, Y(30) => ALU_OP2_30_port, Y(29) => 
                           ALU_OP2_29_port, Y(28) => ALU_OP2_28_port, Y(27) => 
                           ALU_OP2_27_port, Y(26) => ALU_OP2_26_port, Y(25) => 
                           ALU_OP2_25_port, Y(24) => ALU_OP2_24_port, Y(23) => 
                           ALU_OP2_23_port, Y(22) => ALU_OP2_22_port, Y(21) => 
                           ALU_OP2_21_port, Y(20) => ALU_OP2_20_port, Y(19) => 
                           ALU_OP2_19_port, Y(18) => ALU_OP2_18_port, Y(17) => 
                           ALU_OP2_17_port, Y(16) => ALU_OP2_16_port, Y(15) => 
                           ALU_OP2_15_port, Y(14) => ALU_OP2_14_port, Y(13) => 
                           ALU_OP2_13_port, Y(12) => ALU_OP2_12_port, Y(11) => 
                           ALU_OP2_11_port, Y(10) => ALU_OP2_10_port, Y(9) => 
                           ALU_OP2_9_port, Y(8) => ALU_OP2_8_port, Y(7) => 
                           ALU_OP2_7_port, Y(6) => ALU_OP2_6_port, Y(5) => 
                           ALU_OP2_5_port, Y(4) => ALU_OP2_4_port, Y(3) => 
                           ALU_OP2_3_port, Y(2) => ALU_OP2_2_port, Y(1) => 
                           ALU_OP2_1_port, Y(0) => ALU_OP2_0_port);
   ARITHMETIC_LOGIC_UNIT : ALU_N32_NB8 port map( OP1(31) => ALU_OP1_31_port, 
                           OP1(30) => ALU_OP1_30_port, OP1(29) => 
                           ALU_OP1_29_port, OP1(28) => ALU_OP1_28_port, OP1(27)
                           => ALU_OP1_27_port, OP1(26) => ALU_OP1_26_port, 
                           OP1(25) => ALU_OP1_25_port, OP1(24) => 
                           ALU_OP1_24_port, OP1(23) => ALU_OP1_23_port, OP1(22)
                           => ALU_OP1_22_port, OP1(21) => ALU_OP1_21_port, 
                           OP1(20) => ALU_OP1_20_port, OP1(19) => 
                           ALU_OP1_19_port, OP1(18) => ALU_OP1_18_port, OP1(17)
                           => ALU_OP1_17_port, OP1(16) => ALU_OP1_16_port, 
                           OP1(15) => ALU_OP1_15_port, OP1(14) => 
                           ALU_OP1_14_port, OP1(13) => ALU_OP1_13_port, OP1(12)
                           => ALU_OP1_12_port, OP1(11) => ALU_OP1_11_port, 
                           OP1(10) => ALU_OP1_10_port, OP1(9) => ALU_OP1_9_port
                           , OP1(8) => ALU_OP1_8_port, OP1(7) => ALU_OP1_7_port
                           , OP1(6) => ALU_OP1_6_port, OP1(5) => ALU_OP1_5_port
                           , OP1(4) => ALU_OP1_4_port, OP1(3) => ALU_OP1_3_port
                           , OP1(2) => ALU_OP1_2_port, OP1(1) => ALU_OP1_1_port
                           , OP1(0) => ALU_OP1_0_port, OP2(31) => 
                           ALU_OP2_31_port, OP2(30) => ALU_OP2_30_port, OP2(29)
                           => ALU_OP2_29_port, OP2(28) => ALU_OP2_28_port, 
                           OP2(27) => ALU_OP2_27_port, OP2(26) => 
                           ALU_OP2_26_port, OP2(25) => ALU_OP2_25_port, OP2(24)
                           => ALU_OP2_24_port, OP2(23) => ALU_OP2_23_port, 
                           OP2(22) => ALU_OP2_22_port, OP2(21) => 
                           ALU_OP2_21_port, OP2(20) => ALU_OP2_20_port, OP2(19)
                           => ALU_OP2_19_port, OP2(18) => ALU_OP2_18_port, 
                           OP2(17) => ALU_OP2_17_port, OP2(16) => 
                           ALU_OP2_16_port, OP2(15) => ALU_OP2_15_port, OP2(14)
                           => ALU_OP2_14_port, OP2(13) => ALU_OP2_13_port, 
                           OP2(12) => ALU_OP2_12_port, OP2(11) => 
                           ALU_OP2_11_port, OP2(10) => ALU_OP2_10_port, OP2(9) 
                           => ALU_OP2_9_port, OP2(8) => ALU_OP2_8_port, OP2(7) 
                           => ALU_OP2_7_port, OP2(6) => ALU_OP2_6_port, OP2(5) 
                           => ALU_OP2_5_port, OP2(4) => ALU_OP2_4_port, OP2(3) 
                           => ALU_OP2_3_port, OP2(2) => ALU_OP2_2_port, OP2(1) 
                           => ALU_OP2_1_port, OP2(0) => ALU_OP2_0_port, OPC(0) 
                           => ALU_OPCODE(0), OPC(1) => ALU_OPCODE(1), OPC(2) =>
                           ALU_OPCODE(2), OPC(3) => ALU_OPCODE(3), OPC(4) => 
                           ALU_OPCODE(4), OPC(5) => ALU_OPCODE(5), OPC(6) => 
                           ALU_OPCODE(6), Y(31) => ALU_OUTPUT_31_port, Y(30) =>
                           ALU_OUTPUT_30_port, Y(29) => ALU_OUTPUT_29_port, 
                           Y(28) => ALU_OUTPUT_28_port, Y(27) => 
                           ALU_OUTPUT_27_port, Y(26) => ALU_OUTPUT_26_port, 
                           Y(25) => ALU_OUTPUT_25_port, Y(24) => 
                           ALU_OUTPUT_24_port, Y(23) => ALU_OUTPUT_23_port, 
                           Y(22) => ALU_OUTPUT_22_port, Y(21) => 
                           ALU_OUTPUT_21_port, Y(20) => ALU_OUTPUT_20_port, 
                           Y(19) => ALU_OUTPUT_19_port, Y(18) => 
                           ALU_OUTPUT_18_port, Y(17) => ALU_OUTPUT_17_port, 
                           Y(16) => ALU_OUTPUT_16_port, Y(15) => 
                           ALU_OUTPUT_15_port, Y(14) => ALU_OUTPUT_14_port, 
                           Y(13) => ALU_OUTPUT_13_port, Y(12) => 
                           ALU_OUTPUT_12_port, Y(11) => ALU_OUTPUT_11_port, 
                           Y(10) => ALU_OUTPUT_10_port, Y(9) => 
                           ALU_OUTPUT_9_port, Y(8) => ALU_OUTPUT_8_port, Y(7) 
                           => ALU_OUTPUT_7_port, Y(6) => ALU_OUTPUT_6_port, 
                           Y(5) => ALU_OUTPUT_5_port, Y(4) => ALU_OUTPUT_4_port
                           , Y(3) => ALU_OUTPUT_3_port, Y(2) => 
                           ALU_OUTPUT_2_port, Y(1) => ALU_OUTPUT_1_port, Y(0) 
                           => ALU_OUTPUT_0_port, Z => n_1627);
   BRANCH_MUX : MUX21_L_320 port map( A => ZERO_OUT, B => n186_port, S => 
                           EQ_COND, Y => BRANCH_DETECT);
   Z_DETECTOR : ZERO_DETECTOR_N32_1 port map( A(31) => ALU_PREOP1_31_port, 
                           A(30) => ALU_PREOP1_30_port, A(29) => 
                           ALU_PREOP1_29_port, A(28) => ALU_PREOP1_28_port, 
                           A(27) => ALU_PREOP1_27_port, A(26) => 
                           ALU_PREOP1_26_port, A(25) => ALU_PREOP1_25_port, 
                           A(24) => ALU_PREOP1_24_port, A(23) => 
                           ALU_PREOP1_23_port, A(22) => ALU_PREOP1_22_port, 
                           A(21) => ALU_PREOP1_21_port, A(20) => 
                           ALU_PREOP1_20_port, A(19) => ALU_PREOP1_19_port, 
                           A(18) => ALU_PREOP1_18_port, A(17) => 
                           ALU_PREOP1_17_port, A(16) => ALU_PREOP1_16_port, 
                           A(15) => ALU_PREOP1_15_port, A(14) => 
                           ALU_PREOP1_14_port, A(13) => ALU_PREOP1_13_port, 
                           A(12) => ALU_PREOP1_12_port, A(11) => 
                           ALU_PREOP1_11_port, A(10) => ALU_PREOP1_10_port, 
                           A(9) => ALU_PREOP1_9_port, A(8) => ALU_PREOP1_8_port
                           , A(7) => ALU_PREOP1_7_port, A(6) => 
                           ALU_PREOP1_6_port, A(5) => ALU_PREOP1_5_port, A(4) 
                           => ALU_PREOP1_4_port, A(3) => ALU_PREOP1_3_port, 
                           A(2) => ALU_PREOP1_2_port, A(1) => ALU_PREOP1_1_port
                           , A(0) => ALU_PREOP1_0_port, Y => ZERO_OUT);
   FORWARDING_UNIT : FU_N5 port map( RS1(4) => ID_EX_RS1_4_port, RS1(3) => 
                           ID_EX_RS1_3_port, RS1(2) => ID_EX_RS1_2_port, RS1(1)
                           => ID_EX_RS1_1_port, RS1(0) => ID_EX_RS1_0_port, 
                           RS2(4) => ID_EX_RS2_4_port, RS2(3) => 
                           ID_EX_RS2_3_port, RS2(2) => ID_EX_RS2_2_port, RS2(1)
                           => ID_EX_RS2_1_port, RS2(0) => ID_EX_RS2_0_port, 
                           RD_MEM(4) => EX_MEM_RD_4_port, RD_MEM(3) => 
                           EX_MEM_RD_3_port, RD_MEM(2) => EX_MEM_RD_2_port, 
                           RD_MEM(1) => EX_MEM_RD_1_port, RD_MEM(0) => 
                           EX_MEM_RD_0_port, RD_WB(4) => MEM_WB_RD_4_port, 
                           RD_WB(3) => MEM_WB_RD_3_port, RD_WB(2) => 
                           MEM_WB_RD_2_port, RD_WB(1) => MEM_WB_RD_1_port, 
                           RD_WB(0) => MEM_WB_RD_0_port, RF_WE_MEM => 
                           EX_MEM_RF_WE, RF_WE_WB => MEM_WB_RF_WE, FORWARD_A(1)
                           => FORWARD_A_1_port, FORWARD_A(0) => 
                           FORWARD_A_0_port, FORWARD_B(1) => FORWARD_B_1_port, 
                           FORWARD_B(0) => FORWARD_B_0_port);
   LATCH_ALUOUT : LDR_N32_1 port map( RST => RST, EN => ALU_OUTREG_EN, 
                           REGIN(31) => ALU_OUTPUT_31_port, REGIN(30) => 
                           ALU_OUTPUT_30_port, REGIN(29) => ALU_OUTPUT_29_port,
                           REGIN(28) => ALU_OUTPUT_28_port, REGIN(27) => 
                           ALU_OUTPUT_27_port, REGIN(26) => ALU_OUTPUT_26_port,
                           REGIN(25) => ALU_OUTPUT_25_port, REGIN(24) => 
                           ALU_OUTPUT_24_port, REGIN(23) => ALU_OUTPUT_23_port,
                           REGIN(22) => ALU_OUTPUT_22_port, REGIN(21) => 
                           ALU_OUTPUT_21_port, REGIN(20) => ALU_OUTPUT_20_port,
                           REGIN(19) => ALU_OUTPUT_19_port, REGIN(18) => 
                           ALU_OUTPUT_18_port, REGIN(17) => ALU_OUTPUT_17_port,
                           REGIN(16) => ALU_OUTPUT_16_port, REGIN(15) => 
                           ALU_OUTPUT_15_port, REGIN(14) => ALU_OUTPUT_14_port,
                           REGIN(13) => ALU_OUTPUT_13_port, REGIN(12) => 
                           ALU_OUTPUT_12_port, REGIN(11) => ALU_OUTPUT_11_port,
                           REGIN(10) => ALU_OUTPUT_10_port, REGIN(9) => 
                           ALU_OUTPUT_9_port, REGIN(8) => ALU_OUTPUT_8_port, 
                           REGIN(7) => ALU_OUTPUT_7_port, REGIN(6) => 
                           ALU_OUTPUT_6_port, REGIN(5) => ALU_OUTPUT_5_port, 
                           REGIN(4) => ALU_OUTPUT_4_port, REGIN(3) => 
                           ALU_OUTPUT_3_port, REGIN(2) => ALU_OUTPUT_2_port, 
                           REGIN(1) => ALU_OUTPUT_1_port, REGIN(0) => 
                           ALU_OUTPUT_0_port, REGOUT(31) => 
                           EX_MEM_ALU_OUTPUT_NEXT_31_port, REGOUT(30) => 
                           EX_MEM_ALU_OUTPUT_NEXT_30_port, REGOUT(29) => 
                           EX_MEM_ALU_OUTPUT_NEXT_29_port, REGOUT(28) => 
                           EX_MEM_ALU_OUTPUT_NEXT_28_port, REGOUT(27) => 
                           EX_MEM_ALU_OUTPUT_NEXT_27_port, REGOUT(26) => 
                           EX_MEM_ALU_OUTPUT_NEXT_26_port, REGOUT(25) => 
                           EX_MEM_ALU_OUTPUT_NEXT_25_port, REGOUT(24) => 
                           EX_MEM_ALU_OUTPUT_NEXT_24_port, REGOUT(23) => 
                           EX_MEM_ALU_OUTPUT_NEXT_23_port, REGOUT(22) => 
                           EX_MEM_ALU_OUTPUT_NEXT_22_port, REGOUT(21) => 
                           EX_MEM_ALU_OUTPUT_NEXT_21_port, REGOUT(20) => 
                           EX_MEM_ALU_OUTPUT_NEXT_20_port, REGOUT(19) => 
                           EX_MEM_ALU_OUTPUT_NEXT_19_port, REGOUT(18) => 
                           EX_MEM_ALU_OUTPUT_NEXT_18_port, REGOUT(17) => 
                           EX_MEM_ALU_OUTPUT_NEXT_17_port, REGOUT(16) => 
                           EX_MEM_ALU_OUTPUT_NEXT_16_port, REGOUT(15) => 
                           EX_MEM_ALU_OUTPUT_NEXT_15_port, REGOUT(14) => 
                           EX_MEM_ALU_OUTPUT_NEXT_14_port, REGOUT(13) => 
                           EX_MEM_ALU_OUTPUT_NEXT_13_port, REGOUT(12) => 
                           EX_MEM_ALU_OUTPUT_NEXT_12_port, REGOUT(11) => 
                           EX_MEM_ALU_OUTPUT_NEXT_11_port, REGOUT(10) => 
                           EX_MEM_ALU_OUTPUT_NEXT_10_port, REGOUT(9) => 
                           EX_MEM_ALU_OUTPUT_NEXT_9_port, REGOUT(8) => 
                           EX_MEM_ALU_OUTPUT_NEXT_8_port, REGOUT(7) => 
                           EX_MEM_ALU_OUTPUT_NEXT_7_port, REGOUT(6) => 
                           EX_MEM_ALU_OUTPUT_NEXT_6_port, REGOUT(5) => 
                           EX_MEM_ALU_OUTPUT_NEXT_5_port, REGOUT(4) => 
                           EX_MEM_ALU_OUTPUT_NEXT_4_port, REGOUT(3) => 
                           EX_MEM_ALU_OUTPUT_NEXT_3_port, REGOUT(2) => 
                           EX_MEM_ALU_OUTPUT_NEXT_2_port, REGOUT(1) => 
                           EX_MEM_ALU_OUTPUT_NEXT_1_port, REGOUT(0) => 
                           EX_MEM_ALU_OUTPUT_NEXT_0_port);
   LATCH_BRANCH : LD_224 port map( RST => RST, EN => ALU_OUTREG_EN, D => 
                           BRANCH_DETECT, Q => EX_MEM_BRANCH_DETECT_NEXT);
   LATCH_LMD : LDR_N32_0 port map( RST => RST, EN => LMD_LATCH_EN, REGIN(31) =>
                           DRAM_OUT(31), REGIN(30) => DRAM_OUT(30), REGIN(29) 
                           => DRAM_OUT(29), REGIN(28) => DRAM_OUT(28), 
                           REGIN(27) => DRAM_OUT(27), REGIN(26) => DRAM_OUT(26)
                           , REGIN(25) => DRAM_OUT(25), REGIN(24) => 
                           DRAM_OUT(24), REGIN(23) => DRAM_OUT(23), REGIN(22) 
                           => DRAM_OUT(22), REGIN(21) => DRAM_OUT(21), 
                           REGIN(20) => DRAM_OUT(20), REGIN(19) => DRAM_OUT(19)
                           , REGIN(18) => DRAM_OUT(18), REGIN(17) => 
                           DRAM_OUT(17), REGIN(16) => DRAM_OUT(16), REGIN(15) 
                           => DRAM_OUT(15), REGIN(14) => DRAM_OUT(14), 
                           REGIN(13) => DRAM_OUT(13), REGIN(12) => DRAM_OUT(12)
                           , REGIN(11) => DRAM_OUT(11), REGIN(10) => 
                           DRAM_OUT(10), REGIN(9) => DRAM_OUT(9), REGIN(8) => 
                           DRAM_OUT(8), REGIN(7) => DRAM_OUT(7), REGIN(6) => 
                           DRAM_OUT(6), REGIN(5) => DRAM_OUT(5), REGIN(4) => 
                           DRAM_OUT(4), REGIN(3) => DRAM_OUT(3), REGIN(2) => 
                           DRAM_OUT(2), REGIN(1) => DRAM_OUT(1), REGIN(0) => 
                           DRAM_OUT(0), REGOUT(31) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_31_port, REGOUT(30) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_30_port, REGOUT(29) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_29_port, REGOUT(28) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_28_port, REGOUT(27) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_27_port, REGOUT(26) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_26_port, REGOUT(25) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_25_port, REGOUT(24) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_24_port, REGOUT(23) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_23_port, REGOUT(22) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_22_port, REGOUT(21) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_21_port, REGOUT(20) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_20_port, REGOUT(19) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_19_port, REGOUT(18) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_18_port, REGOUT(17) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_17_port, REGOUT(16) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_16_port, REGOUT(15) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_15_port, REGOUT(14) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_14_port, REGOUT(13) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_13_port, REGOUT(12) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_12_port, REGOUT(11) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_11_port, REGOUT(10) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_10_port, REGOUT(9) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_9_port, REGOUT(8) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_8_port, REGOUT(7) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_7_port, REGOUT(6) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_6_port, REGOUT(5) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_5_port, REGOUT(4) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_4_port, REGOUT(3) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_3_port, REGOUT(2) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_2_port, REGOUT(1) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_1_port, REGOUT(0) => 
                           MEM_WB_DRAM_OUTPUT_NEXT_0_port);
   WB_MUX : MUX21_N32_1 port map( A(31) => MEM_WB_DRAM_OUTPUT_31_port, A(30) =>
                           MEM_WB_DRAM_OUTPUT_30_port, A(29) => 
                           MEM_WB_DRAM_OUTPUT_29_port, A(28) => 
                           MEM_WB_DRAM_OUTPUT_28_port, A(27) => 
                           MEM_WB_DRAM_OUTPUT_27_port, A(26) => 
                           MEM_WB_DRAM_OUTPUT_26_port, A(25) => 
                           MEM_WB_DRAM_OUTPUT_25_port, A(24) => 
                           MEM_WB_DRAM_OUTPUT_24_port, A(23) => 
                           MEM_WB_DRAM_OUTPUT_23_port, A(22) => 
                           MEM_WB_DRAM_OUTPUT_22_port, A(21) => 
                           MEM_WB_DRAM_OUTPUT_21_port, A(20) => 
                           MEM_WB_DRAM_OUTPUT_20_port, A(19) => 
                           MEM_WB_DRAM_OUTPUT_19_port, A(18) => 
                           MEM_WB_DRAM_OUTPUT_18_port, A(17) => 
                           MEM_WB_DRAM_OUTPUT_17_port, A(16) => 
                           MEM_WB_DRAM_OUTPUT_16_port, A(15) => 
                           MEM_WB_DRAM_OUTPUT_15_port, A(14) => 
                           MEM_WB_DRAM_OUTPUT_14_port, A(13) => 
                           MEM_WB_DRAM_OUTPUT_13_port, A(12) => 
                           MEM_WB_DRAM_OUTPUT_12_port, A(11) => 
                           MEM_WB_DRAM_OUTPUT_11_port, A(10) => 
                           MEM_WB_DRAM_OUTPUT_10_port, A(9) => 
                           MEM_WB_DRAM_OUTPUT_9_port, A(8) => 
                           MEM_WB_DRAM_OUTPUT_8_port, A(7) => 
                           MEM_WB_DRAM_OUTPUT_7_port, A(6) => 
                           MEM_WB_DRAM_OUTPUT_6_port, A(5) => 
                           MEM_WB_DRAM_OUTPUT_5_port, A(4) => 
                           MEM_WB_DRAM_OUTPUT_4_port, A(3) => 
                           MEM_WB_DRAM_OUTPUT_3_port, A(2) => 
                           MEM_WB_DRAM_OUTPUT_2_port, A(1) => 
                           MEM_WB_DRAM_OUTPUT_1_port, A(0) => 
                           MEM_WB_DRAM_OUTPUT_0_port, B(31) => 
                           MEM_WB_ALU_OUTPUT_31_port, B(30) => 
                           MEM_WB_ALU_OUTPUT_30_port, B(29) => 
                           MEM_WB_ALU_OUTPUT_29_port, B(28) => 
                           MEM_WB_ALU_OUTPUT_28_port, B(27) => 
                           MEM_WB_ALU_OUTPUT_27_port, B(26) => 
                           MEM_WB_ALU_OUTPUT_26_port, B(25) => 
                           MEM_WB_ALU_OUTPUT_25_port, B(24) => 
                           MEM_WB_ALU_OUTPUT_24_port, B(23) => 
                           MEM_WB_ALU_OUTPUT_23_port, B(22) => 
                           MEM_WB_ALU_OUTPUT_22_port, B(21) => 
                           MEM_WB_ALU_OUTPUT_21_port, B(20) => 
                           MEM_WB_ALU_OUTPUT_20_port, B(19) => 
                           MEM_WB_ALU_OUTPUT_19_port, B(18) => 
                           MEM_WB_ALU_OUTPUT_18_port, B(17) => 
                           MEM_WB_ALU_OUTPUT_17_port, B(16) => 
                           MEM_WB_ALU_OUTPUT_16_port, B(15) => 
                           MEM_WB_ALU_OUTPUT_15_port, B(14) => 
                           MEM_WB_ALU_OUTPUT_14_port, B(13) => 
                           MEM_WB_ALU_OUTPUT_13_port, B(12) => 
                           MEM_WB_ALU_OUTPUT_12_port, B(11) => 
                           MEM_WB_ALU_OUTPUT_11_port, B(10) => 
                           MEM_WB_ALU_OUTPUT_10_port, B(9) => 
                           MEM_WB_ALU_OUTPUT_9_port, B(8) => 
                           MEM_WB_ALU_OUTPUT_8_port, B(7) => 
                           MEM_WB_ALU_OUTPUT_7_port, B(6) => 
                           MEM_WB_ALU_OUTPUT_6_port, B(5) => 
                           MEM_WB_ALU_OUTPUT_5_port, B(4) => 
                           MEM_WB_ALU_OUTPUT_4_port, B(3) => 
                           MEM_WB_ALU_OUTPUT_3_port, B(2) => 
                           MEM_WB_ALU_OUTPUT_2_port, B(1) => 
                           MEM_WB_ALU_OUTPUT_1_port, B(0) => 
                           MEM_WB_ALU_OUTPUT_0_port, S => WB_MUX_SEL, Y(31) => 
                           WB_MUX_OUT_31_port, Y(30) => WB_MUX_OUT_30_port, 
                           Y(29) => WB_MUX_OUT_29_port, Y(28) => 
                           WB_MUX_OUT_28_port, Y(27) => WB_MUX_OUT_27_port, 
                           Y(26) => WB_MUX_OUT_26_port, Y(25) => 
                           WB_MUX_OUT_25_port, Y(24) => WB_MUX_OUT_24_port, 
                           Y(23) => WB_MUX_OUT_23_port, Y(22) => 
                           WB_MUX_OUT_22_port, Y(21) => WB_MUX_OUT_21_port, 
                           Y(20) => WB_MUX_OUT_20_port, Y(19) => 
                           WB_MUX_OUT_19_port, Y(18) => WB_MUX_OUT_18_port, 
                           Y(17) => WB_MUX_OUT_17_port, Y(16) => 
                           WB_MUX_OUT_16_port, Y(15) => WB_MUX_OUT_15_port, 
                           Y(14) => WB_MUX_OUT_14_port, Y(13) => 
                           WB_MUX_OUT_13_port, Y(12) => WB_MUX_OUT_12_port, 
                           Y(11) => WB_MUX_OUT_11_port, Y(10) => 
                           WB_MUX_OUT_10_port, Y(9) => WB_MUX_OUT_9_port, Y(8) 
                           => WB_MUX_OUT_8_port, Y(7) => WB_MUX_OUT_7_port, 
                           Y(6) => WB_MUX_OUT_6_port, Y(5) => WB_MUX_OUT_5_port
                           , Y(4) => WB_MUX_OUT_4_port, Y(3) => 
                           WB_MUX_OUT_3_port, Y(2) => WB_MUX_OUT_2_port, Y(1) 
                           => WB_MUX_OUT_1_port, Y(0) => WB_MUX_OUT_0_port);
   JAL_MUX : MUX21_N32_0 port map( A(31) => WB_MUX_OUT_31_port, A(30) => 
                           WB_MUX_OUT_30_port, A(29) => WB_MUX_OUT_29_port, 
                           A(28) => WB_MUX_OUT_28_port, A(27) => 
                           WB_MUX_OUT_27_port, A(26) => WB_MUX_OUT_26_port, 
                           A(25) => WB_MUX_OUT_25_port, A(24) => 
                           WB_MUX_OUT_24_port, A(23) => WB_MUX_OUT_23_port, 
                           A(22) => WB_MUX_OUT_22_port, A(21) => 
                           WB_MUX_OUT_21_port, A(20) => WB_MUX_OUT_20_port, 
                           A(19) => WB_MUX_OUT_19_port, A(18) => 
                           WB_MUX_OUT_18_port, A(17) => WB_MUX_OUT_17_port, 
                           A(16) => WB_MUX_OUT_16_port, A(15) => 
                           WB_MUX_OUT_15_port, A(14) => WB_MUX_OUT_14_port, 
                           A(13) => WB_MUX_OUT_13_port, A(12) => 
                           WB_MUX_OUT_12_port, A(11) => WB_MUX_OUT_11_port, 
                           A(10) => WB_MUX_OUT_10_port, A(9) => 
                           WB_MUX_OUT_9_port, A(8) => WB_MUX_OUT_8_port, A(7) 
                           => WB_MUX_OUT_7_port, A(6) => WB_MUX_OUT_6_port, 
                           A(5) => WB_MUX_OUT_5_port, A(4) => WB_MUX_OUT_4_port
                           , A(3) => WB_MUX_OUT_3_port, A(2) => 
                           WB_MUX_OUT_2_port, A(1) => WB_MUX_OUT_1_port, A(0) 
                           => WB_MUX_OUT_0_port, B(31) => MEM_WB_NPC_31_port, 
                           B(30) => MEM_WB_NPC_30_port, B(29) => 
                           MEM_WB_NPC_29_port, B(28) => MEM_WB_NPC_28_port, 
                           B(27) => MEM_WB_NPC_27_port, B(26) => 
                           MEM_WB_NPC_26_port, B(25) => MEM_WB_NPC_25_port, 
                           B(24) => MEM_WB_NPC_24_port, B(23) => 
                           MEM_WB_NPC_23_port, B(22) => MEM_WB_NPC_22_port, 
                           B(21) => MEM_WB_NPC_21_port, B(20) => 
                           MEM_WB_NPC_20_port, B(19) => MEM_WB_NPC_19_port, 
                           B(18) => MEM_WB_NPC_18_port, B(17) => 
                           MEM_WB_NPC_17_port, B(16) => MEM_WB_NPC_16_port, 
                           B(15) => MEM_WB_NPC_15_port, B(14) => 
                           MEM_WB_NPC_14_port, B(13) => MEM_WB_NPC_13_port, 
                           B(12) => MEM_WB_NPC_12_port, B(11) => 
                           MEM_WB_NPC_11_port, B(10) => MEM_WB_NPC_10_port, 
                           B(9) => MEM_WB_NPC_9_port, B(8) => MEM_WB_NPC_8_port
                           , B(7) => MEM_WB_NPC_7_port, B(6) => 
                           MEM_WB_NPC_6_port, B(5) => MEM_WB_NPC_5_port, B(4) 
                           => MEM_WB_NPC_4_port, B(3) => MEM_WB_NPC_3_port, 
                           B(2) => MEM_WB_NPC_2_port, B(1) => MEM_WB_NPC_1_port
                           , B(0) => MEM_WB_NPC_0_port, S => JAL_MUX_SEL, Y(31)
                           => JAL_MUX_OUT_31_port, Y(30) => JAL_MUX_OUT_30_port
                           , Y(29) => JAL_MUX_OUT_29_port, Y(28) => 
                           JAL_MUX_OUT_28_port, Y(27) => JAL_MUX_OUT_27_port, 
                           Y(26) => JAL_MUX_OUT_26_port, Y(25) => 
                           JAL_MUX_OUT_25_port, Y(24) => JAL_MUX_OUT_24_port, 
                           Y(23) => JAL_MUX_OUT_23_port, Y(22) => 
                           JAL_MUX_OUT_22_port, Y(21) => JAL_MUX_OUT_21_port, 
                           Y(20) => JAL_MUX_OUT_20_port, Y(19) => 
                           JAL_MUX_OUT_19_port, Y(18) => JAL_MUX_OUT_18_port, 
                           Y(17) => JAL_MUX_OUT_17_port, Y(16) => 
                           JAL_MUX_OUT_16_port, Y(15) => JAL_MUX_OUT_15_port, 
                           Y(14) => JAL_MUX_OUT_14_port, Y(13) => 
                           JAL_MUX_OUT_13_port, Y(12) => JAL_MUX_OUT_12_port, 
                           Y(11) => JAL_MUX_OUT_11_port, Y(10) => 
                           JAL_MUX_OUT_10_port, Y(9) => JAL_MUX_OUT_9_port, 
                           Y(8) => JAL_MUX_OUT_8_port, Y(7) => 
                           JAL_MUX_OUT_7_port, Y(6) => JAL_MUX_OUT_6_port, Y(5)
                           => JAL_MUX_OUT_5_port, Y(4) => JAL_MUX_OUT_4_port, 
                           Y(3) => JAL_MUX_OUT_3_port, Y(2) => 
                           JAL_MUX_OUT_2_port, Y(1) => JAL_MUX_OUT_1_port, Y(0)
                           => JAL_MUX_OUT_0_port);
   add_630 : 
                           DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32_DW01_add_0 
                           port map( A(31) => PC_OUT_31_port, A(30) => 
                           PC_OUT_30_port, A(29) => PC_OUT_29_port, A(28) => 
                           PC_OUT_28_port, A(27) => PC_OUT_27_port, A(26) => 
                           PC_OUT_26_port, A(25) => PC_OUT_25_port, A(24) => 
                           PC_OUT_24_port, A(23) => PC_OUT_23_port, A(22) => 
                           PC_OUT_22_port, A(21) => PC_OUT_21_port, A(20) => 
                           PC_OUT_20_port, A(19) => PC_OUT_19_port, A(18) => 
                           PC_OUT_18_port, A(17) => PC_OUT_17_port, A(16) => 
                           PC_OUT_16_port, A(15) => PC_OUT_15_port, A(14) => 
                           PC_OUT_14_port, A(13) => PC_OUT_13_port, A(12) => 
                           PC_OUT_12_port, A(11) => PC_OUT_11_port, A(10) => 
                           PC_OUT_10_port, A(9) => PC_OUT_9_port, A(8) => 
                           PC_OUT_8_port, A(7) => PC_OUT_7_port, A(6) => 
                           PC_OUT_6_port, A(5) => PC_OUT_5_port, A(4) => 
                           PC_OUT_4_port, A(3) => PC_OUT_3_port, A(2) => 
                           PC_OUT_2_port, A(1) => PC_OUT_1_port, A(0) => 
                           PC_OUT_0_port, B(31) => n1, B(30) => n1, B(29) => n1
                           , B(28) => n1, B(27) => n1, B(26) => n1, B(25) => n1
                           , B(24) => n1, B(23) => n1, B(22) => n1, B(21) => n1
                           , B(20) => n1, B(19) => n1, B(18) => n1, B(17) => n1
                           , B(16) => n1, B(15) => n1, B(14) => n1, B(13) => n1
                           , B(12) => n1, B(11) => n1, B(10) => n1, B(9) => n1,
                           B(8) => n1, B(7) => n1, B(6) => n1, B(5) => n1, B(4)
                           => n1, B(3) => n1, B(2) => X_Logic1_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, CI => n1, 
                           SUM(31) => NPC_BUS_31_port, SUM(30) => 
                           NPC_BUS_30_port, SUM(29) => NPC_BUS_29_port, SUM(28)
                           => NPC_BUS_28_port, SUM(27) => NPC_BUS_27_port, 
                           SUM(26) => NPC_BUS_26_port, SUM(25) => 
                           NPC_BUS_25_port, SUM(24) => NPC_BUS_24_port, SUM(23)
                           => NPC_BUS_23_port, SUM(22) => NPC_BUS_22_port, 
                           SUM(21) => NPC_BUS_21_port, SUM(20) => 
                           NPC_BUS_20_port, SUM(19) => NPC_BUS_19_port, SUM(18)
                           => NPC_BUS_18_port, SUM(17) => NPC_BUS_17_port, 
                           SUM(16) => NPC_BUS_16_port, SUM(15) => 
                           NPC_BUS_15_port, SUM(14) => NPC_BUS_14_port, SUM(13)
                           => NPC_BUS_13_port, SUM(12) => NPC_BUS_12_port, 
                           SUM(11) => NPC_BUS_11_port, SUM(10) => 
                           NPC_BUS_10_port, SUM(9) => NPC_BUS_9_port, SUM(8) =>
                           NPC_BUS_8_port, SUM(7) => NPC_BUS_7_port, SUM(6) => 
                           NPC_BUS_6_port, SUM(5) => NPC_BUS_5_port, SUM(4) => 
                           NPC_BUS_4_port, SUM(3) => NPC_BUS_3_port, SUM(2) => 
                           NPC_BUS_2_port, SUM(1) => NPC_BUS_1_port, SUM(0) => 
                           NPC_BUS_0_port, CO => n_1628);
   U3 : BUF_X1 port map( A => n7_port, Z => n2_port);
   U5 : INV_X2 port map( A => n13_port, ZN => n187_port);
   U6 : BUF_X1 port map( A => n8_port, Z => n6_port);
   U7 : BUF_X1 port map( A => CLK, Z => n12_port);
   U8 : CLKBUF_X3 port map( A => n6_port, Z => n4_port);
   U9 : CLKBUF_X3 port map( A => n6_port, Z => n3_port);
   U10 : BUF_X2 port map( A => n6_port, Z => n5_port);
   U11 : BUF_X8 port map( A => n12_port, Z => n9_port);
   U12 : BUF_X8 port map( A => n12_port, Z => n10_port);
   U13 : BUF_X1 port map( A => n8_port, Z => n7_port);
   U14 : BUF_X2 port map( A => n12_port, Z => n11_port);
   U15 : INV_X1 port map( A => RST, ZN => n8_port);
   U16 : INV_X1 port map( A => ZERO_OUT, ZN => n186_port);
   U17 : AOI21_X1 port map( B1 => JUMP_EN, B2 => EX_MEM_BRANCH_DETECT, A => 
                           JUMP_COND, ZN => n13_port);
   U18 : AND2_X1 port map( A1 => RST, A2 => ID_EX_RS1_NEXT_0_port, ZN => N99);
   U19 : AND2_X1 port map( A1 => RF_WE, A2 => RST, ZN => N98);
   U20 : NOR2_X1 port map( A1 => n14_port, A2 => n5_port, ZN => N97);
   U21 : NOR2_X1 port map( A1 => n15_port, A2 => n5_port, ZN => N96);
   U22 : NOR2_X1 port map( A1 => n16_port, A2 => n5_port, ZN => N95);
   U23 : NOR2_X1 port map( A1 => n17_port, A2 => n5_port, ZN => N94);
   U24 : NOR2_X1 port map( A1 => n18_port, A2 => n5_port, ZN => N93);
   U25 : NOR2_X1 port map( A1 => n19_port, A2 => n5_port, ZN => N92);
   U26 : NOR2_X1 port map( A1 => n20_port, A2 => n5_port, ZN => N91);
   U27 : NOR2_X1 port map( A1 => n21_port, A2 => n5_port, ZN => N90);
   U28 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_7_port, A2 => RST, ZN => N9);
   U29 : NOR2_X1 port map( A1 => n22_port, A2 => n5_port, ZN => N89);
   U30 : NOR2_X1 port map( A1 => n23_port, A2 => n5_port, ZN => N88);
   U31 : NOR2_X1 port map( A1 => n24_port, A2 => n5_port, ZN => N87);
   U32 : NOR2_X1 port map( A1 => n25_port, A2 => n5_port, ZN => N86);
   U33 : NOR2_X1 port map( A1 => n26_port, A2 => n5_port, ZN => N85);
   U34 : NOR2_X1 port map( A1 => n27_port, A2 => n5_port, ZN => N84);
   U35 : NOR2_X1 port map( A1 => n28_port, A2 => n5_port, ZN => N83);
   U36 : NOR2_X1 port map( A1 => n29_port, A2 => n5_port, ZN => N82);
   U37 : NOR2_X1 port map( A1 => n30_port, A2 => n5_port, ZN => N81);
   U38 : NOR2_X1 port map( A1 => n31_port, A2 => n5_port, ZN => N80);
   U39 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_6_port, A2 => RST, ZN => N8);
   U40 : NOR2_X1 port map( A1 => n32_port, A2 => n5_port, ZN => N79);
   U41 : NOR2_X1 port map( A1 => n33_port, A2 => n5_port, ZN => N78);
   U42 : NOR2_X1 port map( A1 => n34_port, A2 => n5_port, ZN => N77);
   U43 : NOR2_X1 port map( A1 => n35_port, A2 => n5_port, ZN => N76);
   U44 : NOR2_X1 port map( A1 => n36_port, A2 => n5_port, ZN => N75);
   U45 : NOR2_X1 port map( A1 => n37_port, A2 => n5_port, ZN => N74);
   U46 : NOR2_X1 port map( A1 => n38_port, A2 => n5_port, ZN => N73);
   U47 : NOR2_X1 port map( A1 => n39_port, A2 => n5_port, ZN => N72);
   U48 : NOR2_X1 port map( A1 => n40_port, A2 => n5_port, ZN => N71);
   U49 : NOR2_X1 port map( A1 => n41_port, A2 => n5_port, ZN => N70);
   U50 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_5_port, A2 => RST, ZN => N7);
   U51 : NOR2_X1 port map( A1 => n42_port, A2 => n5_port, ZN => N69);
   U52 : NOR2_X1 port map( A1 => n43_port, A2 => n5_port, ZN => N68);
   U53 : NOR2_X1 port map( A1 => n44_port, A2 => n5_port, ZN => N67);
   U54 : NOR2_X1 port map( A1 => n45_port, A2 => n5_port, ZN => N66);
   U55 : AND2_X1 port map( A1 => IR_OUT_31_port, A2 => RST, ZN => N65);
   U56 : AND2_X1 port map( A1 => IR_OUT_30_port, A2 => RST, ZN => N64);
   U57 : AND2_X1 port map( A1 => IR_OUT_29_port, A2 => RST, ZN => N63);
   U58 : AND2_X1 port map( A1 => IR_OUT_28_port, A2 => RST, ZN => N62);
   U59 : AND2_X1 port map( A1 => IR_OUT_27_port, A2 => RST, ZN => N61);
   U60 : AND2_X1 port map( A1 => IR_OUT_26_port, A2 => RST, ZN => N60);
   U61 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_4_port, A2 => RST, ZN => N6);
   U62 : AND2_X1 port map( A1 => IR_OUT_25_port, A2 => RST, ZN => N59);
   U63 : AND2_X1 port map( A1 => IR_OUT_24_port, A2 => RST, ZN => N58);
   U64 : AND2_X1 port map( A1 => IR_OUT_23_port, A2 => RST, ZN => N57);
   U65 : AND2_X1 port map( A1 => IR_OUT_22_port, A2 => RST, ZN => N56);
   U66 : AND2_X1 port map( A1 => IR_OUT_21_port, A2 => RST, ZN => N55);
   U67 : AND2_X1 port map( A1 => IR_OUT_20_port, A2 => RST, ZN => N54);
   U68 : AND2_X1 port map( A1 => IR_OUT_19_port, A2 => RST, ZN => N53);
   U69 : AND2_X1 port map( A1 => IR_OUT_18_port, A2 => RST, ZN => N52);
   U70 : AND2_X1 port map( A1 => IR_OUT_17_port, A2 => RST, ZN => N51);
   U71 : AND2_X1 port map( A1 => IR_OUT_16_port, A2 => RST, ZN => N50);
   U72 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_3_port, A2 => RST, ZN => N5);
   U73 : AND2_X1 port map( A1 => IR_OUT_15_port, A2 => RST, ZN => N49);
   U74 : AND2_X1 port map( A1 => IR_OUT_14_port, A2 => RST, ZN => N48);
   U75 : AND2_X1 port map( A1 => IR_OUT_13_port, A2 => RST, ZN => N47);
   U76 : AND2_X1 port map( A1 => IR_OUT_12_port, A2 => RST, ZN => N46);
   U77 : AND2_X1 port map( A1 => IR_OUT_11_port, A2 => RST, ZN => N45);
   U78 : AND2_X1 port map( A1 => IR_OUT_10_port, A2 => RST, ZN => N44);
   U79 : AND2_X1 port map( A1 => IR_OUT_9_port, A2 => RST, ZN => N43);
   U80 : AND2_X1 port map( A1 => IR_OUT_8_port, A2 => RST, ZN => N42);
   U81 : NOR2_X1 port map( A1 => n46_port, A2 => n4_port, ZN => N414);
   U82 : NOR2_X1 port map( A1 => n47_port, A2 => n4_port, ZN => N413);
   U83 : NOR2_X1 port map( A1 => n48_port, A2 => n4_port, ZN => N412);
   U84 : NOR2_X1 port map( A1 => n49_port, A2 => n4_port, ZN => N411);
   U85 : NOR2_X1 port map( A1 => n50_port, A2 => n4_port, ZN => N410);
   U86 : AND2_X1 port map( A1 => IR_OUT_7_port, A2 => RST, ZN => N41);
   U87 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_31_port, A2 => RST, ZN
                           => N409);
   U88 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_30_port, A2 => RST, ZN
                           => N408);
   U89 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_29_port, A2 => RST, ZN
                           => N407);
   U90 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_28_port, A2 => RST, ZN
                           => N406);
   U91 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_27_port, A2 => RST, ZN
                           => N405);
   U92 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_26_port, A2 => RST, ZN
                           => N404);
   U93 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_25_port, A2 => RST, ZN
                           => N403);
   U94 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_24_port, A2 => RST, ZN
                           => N402);
   U95 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_23_port, A2 => RST, ZN
                           => N401);
   U96 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_22_port, A2 => RST, ZN
                           => N400);
   U97 : AND2_X1 port map( A1 => IR_OUT_6_port, A2 => RST, ZN => N40);
   U98 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_2_port, A2 => RST, ZN => N4);
   U99 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_21_port, A2 => RST, ZN
                           => N399);
   U100 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_20_port, A2 => RST, 
                           ZN => N398);
   U101 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_19_port, A2 => RST, 
                           ZN => N397);
   U102 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_18_port, A2 => RST, 
                           ZN => N396);
   U103 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_17_port, A2 => RST, 
                           ZN => N395);
   U104 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_16_port, A2 => RST, 
                           ZN => N394);
   U105 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_15_port, A2 => RST, 
                           ZN => N393);
   U106 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_14_port, A2 => RST, 
                           ZN => N392);
   U107 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_13_port, A2 => RST, 
                           ZN => N391);
   U108 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_12_port, A2 => RST, 
                           ZN => N390);
   U109 : AND2_X1 port map( A1 => IR_OUT_5_port, A2 => RST, ZN => N39);
   U110 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_11_port, A2 => RST, 
                           ZN => N389);
   U111 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_10_port, A2 => RST, 
                           ZN => N388);
   U112 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_9_port, A2 => RST, ZN
                           => N387);
   U113 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_8_port, A2 => RST, ZN
                           => N386);
   U114 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_7_port, A2 => RST, ZN
                           => N385);
   U115 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_6_port, A2 => RST, ZN
                           => N384);
   U116 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_5_port, A2 => RST, ZN
                           => N383);
   U117 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_4_port, A2 => RST, ZN
                           => N382);
   U118 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_3_port, A2 => RST, ZN
                           => N381);
   U119 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_2_port, A2 => RST, ZN
                           => N380);
   U120 : AND2_X1 port map( A1 => IR_OUT_4_port, A2 => RST, ZN => N38);
   U121 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_1_port, A2 => RST, ZN
                           => N379);
   U122 : AND2_X1 port map( A1 => MEM_WB_DRAM_OUTPUT_NEXT_0_port, A2 => RST, ZN
                           => N378);
   U123 : NOR2_X1 port map( A1 => n51_port, A2 => n4_port, ZN => N377);
   U124 : NOR2_X1 port map( A1 => n52_port, A2 => n4_port, ZN => N376);
   U125 : NOR2_X1 port map( A1 => n53_port, A2 => n4_port, ZN => N375);
   U126 : NOR2_X1 port map( A1 => n54_port, A2 => n4_port, ZN => N374);
   U127 : NOR2_X1 port map( A1 => n55_port, A2 => n4_port, ZN => N373);
   U128 : NOR2_X1 port map( A1 => n56_port, A2 => n4_port, ZN => N372);
   U129 : NOR2_X1 port map( A1 => n57_port, A2 => n4_port, ZN => N371);
   U130 : NOR2_X1 port map( A1 => n58_port, A2 => n4_port, ZN => N370);
   U131 : AND2_X1 port map( A1 => IR_OUT_3_port, A2 => RST, ZN => N37);
   U132 : NOR2_X1 port map( A1 => n59_port, A2 => n4_port, ZN => N369);
   U133 : NOR2_X1 port map( A1 => n60_port, A2 => n4_port, ZN => N368);
   U134 : NOR2_X1 port map( A1 => n61_port, A2 => n4_port, ZN => N367);
   U135 : NOR2_X1 port map( A1 => n62_port, A2 => n4_port, ZN => N366);
   U136 : NOR2_X1 port map( A1 => n63_port, A2 => n4_port, ZN => N365);
   U137 : NOR2_X1 port map( A1 => n64_port, A2 => n4_port, ZN => N364);
   U138 : NOR2_X1 port map( A1 => n65_port, A2 => n4_port, ZN => N363);
   U139 : NOR2_X1 port map( A1 => n66_port, A2 => n4_port, ZN => N362);
   U140 : NOR2_X1 port map( A1 => n67_port, A2 => n4_port, ZN => N361);
   U141 : NOR2_X1 port map( A1 => n68_port, A2 => n4_port, ZN => N360);
   U142 : AND2_X1 port map( A1 => IR_OUT_2_port, A2 => RST, ZN => N36);
   U143 : NOR2_X1 port map( A1 => n69_port, A2 => n4_port, ZN => N359);
   U144 : NOR2_X1 port map( A1 => n70_port, A2 => n4_port, ZN => N358);
   U145 : NOR2_X1 port map( A1 => n71_port, A2 => n4_port, ZN => N357);
   U146 : NOR2_X1 port map( A1 => n72_port, A2 => n4_port, ZN => N356);
   U147 : NOR2_X1 port map( A1 => n73_port, A2 => n4_port, ZN => N355);
   U148 : NOR2_X1 port map( A1 => n74_port, A2 => n4_port, ZN => N354);
   U149 : NOR2_X1 port map( A1 => n75_port, A2 => n4_port, ZN => N353);
   U150 : NOR2_X1 port map( A1 => n76_port, A2 => n4_port, ZN => N352);
   U151 : NOR2_X1 port map( A1 => n77_port, A2 => n4_port, ZN => N351);
   U152 : NOR2_X1 port map( A1 => n78_port, A2 => n4_port, ZN => N350);
   U153 : AND2_X1 port map( A1 => IR_OUT_1_port, A2 => RST, ZN => N35);
   U154 : NOR2_X1 port map( A1 => n79_port, A2 => n4_port, ZN => N349);
   U155 : NOR2_X1 port map( A1 => n80_port, A2 => n4_port, ZN => N348);
   U156 : NOR2_X1 port map( A1 => n81_port, A2 => n4_port, ZN => N347);
   U157 : NOR2_X1 port map( A1 => n82_port, A2 => n4_port, ZN => N346);
   U158 : NOR2_X1 port map( A1 => n83_port, A2 => n4_port, ZN => N345);
   U159 : NOR2_X1 port map( A1 => n84_port, A2 => n4_port, ZN => N344);
   U160 : NOR2_X1 port map( A1 => n85_port, A2 => n4_port, ZN => N343);
   U161 : NOR2_X1 port map( A1 => n86_port, A2 => n4_port, ZN => N342);
   U162 : NOR2_X1 port map( A1 => n87_port, A2 => n4_port, ZN => N341);
   U163 : NOR2_X1 port map( A1 => n88_port, A2 => n4_port, ZN => N340);
   U164 : AND2_X1 port map( A1 => IR_OUT_0_port, A2 => RST, ZN => N34);
   U165 : NOR2_X1 port map( A1 => n89_port, A2 => n4_port, ZN => N339);
   U166 : NOR2_X1 port map( A1 => n90_port, A2 => n4_port, ZN => N338);
   U167 : NOR2_X1 port map( A1 => n91_port, A2 => n4_port, ZN => N337);
   U168 : NOR2_X1 port map( A1 => n92_port, A2 => n4_port, ZN => N336);
   U169 : NOR2_X1 port map( A1 => n93_port, A2 => n4_port, ZN => N335);
   U170 : NOR2_X1 port map( A1 => n94_port, A2 => n4_port, ZN => N334);
   U171 : NOR2_X1 port map( A1 => n95_port, A2 => n4_port, ZN => N333);
   U172 : NOR2_X1 port map( A1 => n96_port, A2 => n4_port, ZN => N332);
   U173 : NOR2_X1 port map( A1 => n97_port, A2 => n4_port, ZN => N331);
   U174 : NOR2_X1 port map( A1 => n98_port, A2 => n4_port, ZN => N330);
   U175 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_31_port, A2 => RST, ZN => N33)
                           ;
   U176 : NOR2_X1 port map( A1 => n99_port, A2 => n4_port, ZN => N329);
   U177 : NOR2_X1 port map( A1 => n100_port, A2 => n4_port, ZN => N328);
   U178 : NOR2_X1 port map( A1 => n101_port, A2 => n4_port, ZN => N327);
   U179 : NOR2_X1 port map( A1 => n102_port, A2 => n4_port, ZN => N326);
   U180 : NOR2_X1 port map( A1 => n103_port, A2 => n4_port, ZN => N325);
   U181 : NOR2_X1 port map( A1 => n104_port, A2 => n4_port, ZN => N324);
   U182 : NOR2_X1 port map( A1 => n105_port, A2 => n4_port, ZN => N323);
   U183 : NOR2_X1 port map( A1 => n106_port, A2 => n3_port, ZN => N322);
   U184 : NOR2_X1 port map( A1 => n107_port, A2 => n3_port, ZN => N321);
   U185 : NOR2_X1 port map( A1 => n108_port, A2 => n3_port, ZN => N320);
   U186 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_30_port, A2 => RST, ZN => N32)
                           ;
   U187 : NOR2_X1 port map( A1 => n109_port, A2 => n3_port, ZN => N319);
   U188 : NOR2_X1 port map( A1 => n110_port, A2 => n3_port, ZN => N318);
   U189 : NOR2_X1 port map( A1 => n111_port, A2 => n3_port, ZN => N317);
   U190 : NOR2_X1 port map( A1 => n112_port, A2 => n3_port, ZN => N316);
   U191 : NOR2_X1 port map( A1 => n113_port, A2 => n3_port, ZN => N315);
   U192 : NOR2_X1 port map( A1 => n114_port, A2 => n3_port, ZN => N314);
   U193 : NOR2_X1 port map( A1 => n115_port, A2 => n3_port, ZN => N313);
   U194 : NOR2_X1 port map( A1 => n116_port, A2 => n3_port, ZN => N312);
   U195 : NOR2_X1 port map( A1 => n117_port, A2 => n3_port, ZN => N311);
   U196 : NOR2_X1 port map( A1 => n118_port, A2 => n3_port, ZN => N310);
   U197 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_29_port, A2 => RST, ZN => N31)
                           ;
   U198 : NOR2_X1 port map( A1 => n119_port, A2 => n3_port, ZN => N309);
   U199 : NOR2_X1 port map( A1 => n120_port, A2 => n3_port, ZN => N308);
   U200 : AND2_X1 port map( A1 => EX_MEM_BRANCH_DETECT_NEXT, A2 => RST, ZN => 
                           N307);
   U201 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_31_port, A2 => RST, ZN
                           => N306);
   U202 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_30_port, A2 => RST, ZN
                           => N305);
   U203 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_29_port, A2 => RST, ZN
                           => N304);
   U204 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_28_port, A2 => RST, ZN
                           => N303);
   U205 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_27_port, A2 => RST, ZN
                           => N302);
   U206 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_26_port, A2 => RST, ZN
                           => N301);
   U207 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_25_port, A2 => RST, ZN
                           => N300);
   U208 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_28_port, A2 => RST, ZN => N30)
                           ;
   U209 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_1_port, A2 => RST, ZN => N3);
   U210 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_24_port, A2 => RST, ZN
                           => N299);
   U211 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_23_port, A2 => RST, ZN
                           => N298);
   U212 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_22_port, A2 => RST, ZN
                           => N297);
   U213 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_21_port, A2 => RST, ZN
                           => N296);
   U214 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_20_port, A2 => RST, ZN
                           => N295);
   U215 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_19_port, A2 => RST, ZN
                           => N294);
   U216 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_18_port, A2 => RST, ZN
                           => N293);
   U217 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_17_port, A2 => RST, ZN
                           => N292);
   U218 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_16_port, A2 => RST, ZN
                           => N291);
   U219 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_15_port, A2 => RST, ZN
                           => N290);
   U220 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_27_port, A2 => RST, ZN => N29)
                           ;
   U221 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_14_port, A2 => RST, ZN
                           => N289);
   U222 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_13_port, A2 => RST, ZN
                           => N288);
   U223 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_12_port, A2 => RST, ZN
                           => N287);
   U224 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_11_port, A2 => RST, ZN
                           => N286);
   U225 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_10_port, A2 => RST, ZN
                           => N285);
   U226 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_9_port, A2 => RST, ZN 
                           => N284);
   U227 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_8_port, A2 => RST, ZN 
                           => N283);
   U228 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_7_port, A2 => RST, ZN 
                           => N282);
   U229 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_6_port, A2 => RST, ZN 
                           => N281);
   U230 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_5_port, A2 => RST, ZN 
                           => N280);
   U231 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_26_port, A2 => RST, ZN => N28)
                           ;
   U232 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_4_port, A2 => RST, ZN 
                           => N279);
   U233 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_3_port, A2 => RST, ZN 
                           => N278);
   U234 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_2_port, A2 => RST, ZN 
                           => N277);
   U235 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_1_port, A2 => RST, ZN 
                           => N276);
   U236 : AND2_X1 port map( A1 => EX_MEM_ALU_OUTPUT_NEXT_0_port, A2 => RST, ZN 
                           => N275);
   U237 : NOR2_X1 port map( A1 => n121_port, A2 => n3_port, ZN => N274);
   U238 : NOR2_X1 port map( A1 => n122_port, A2 => n3_port, ZN => N273);
   U239 : NOR2_X1 port map( A1 => n123_port, A2 => n3_port, ZN => N272);
   U240 : NOR2_X1 port map( A1 => n124_port, A2 => n3_port, ZN => N271);
   U241 : NOR2_X1 port map( A1 => n125_port, A2 => n3_port, ZN => N270);
   U242 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_25_port, A2 => RST, ZN => N27)
                           ;
   U243 : NOR2_X1 port map( A1 => n126_port, A2 => n3_port, ZN => N269);
   U244 : NOR2_X1 port map( A1 => n127_port, A2 => n3_port, ZN => N268);
   U245 : NOR2_X1 port map( A1 => n128_port, A2 => n3_port, ZN => N267);
   U246 : NOR2_X1 port map( A1 => n129_port, A2 => n3_port, ZN => N266);
   U247 : NOR2_X1 port map( A1 => n130_port, A2 => n3_port, ZN => N265);
   U248 : NOR2_X1 port map( A1 => n131_port, A2 => n3_port, ZN => N264);
   U249 : NOR2_X1 port map( A1 => n132_port, A2 => n3_port, ZN => N263);
   U250 : NOR2_X1 port map( A1 => n133_port, A2 => n3_port, ZN => N262);
   U251 : NOR2_X1 port map( A1 => n134_port, A2 => n3_port, ZN => N261);
   U252 : NOR2_X1 port map( A1 => n135_port, A2 => n3_port, ZN => N260);
   U253 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_24_port, A2 => RST, ZN => N26)
                           ;
   U254 : NOR2_X1 port map( A1 => n136_port, A2 => n3_port, ZN => N259);
   U255 : NOR2_X1 port map( A1 => n137_port, A2 => n3_port, ZN => N258);
   U256 : NOR2_X1 port map( A1 => n138_port, A2 => n3_port, ZN => N257);
   U257 : NOR2_X1 port map( A1 => n139_port, A2 => n3_port, ZN => N256);
   U258 : NOR2_X1 port map( A1 => n140_port, A2 => n3_port, ZN => N255);
   U259 : NOR2_X1 port map( A1 => n141_port, A2 => n3_port, ZN => N254);
   U260 : NOR2_X1 port map( A1 => n142_port, A2 => n3_port, ZN => N253);
   U261 : NOR2_X1 port map( A1 => n143_port, A2 => n3_port, ZN => N252);
   U262 : NOR2_X1 port map( A1 => n144_port, A2 => n3_port, ZN => N251);
   U263 : NOR2_X1 port map( A1 => n145_port, A2 => n3_port, ZN => N250);
   U264 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_23_port, A2 => RST, ZN => N25)
                           ;
   U265 : NOR2_X1 port map( A1 => n146_port, A2 => n3_port, ZN => N249);
   U266 : NOR2_X1 port map( A1 => n147_port, A2 => n3_port, ZN => N248);
   U267 : NOR2_X1 port map( A1 => n148_port, A2 => n3_port, ZN => N247);
   U268 : NOR2_X1 port map( A1 => n149_port, A2 => n3_port, ZN => N246);
   U269 : NOR2_X1 port map( A1 => n150_port, A2 => n3_port, ZN => N245);
   U270 : NOR2_X1 port map( A1 => n151_port, A2 => n3_port, ZN => N244);
   U271 : NOR2_X1 port map( A1 => n152_port, A2 => n3_port, ZN => N243);
   U272 : NOR2_X1 port map( A1 => n153_port, A2 => n3_port, ZN => N242);
   U273 : NOR2_X1 port map( A1 => n154_port, A2 => n3_port, ZN => N241);
   U274 : NOR2_X1 port map( A1 => n155_port, A2 => n3_port, ZN => N240);
   U275 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_22_port, A2 => RST, ZN => N24)
                           ;
   U276 : NOR2_X1 port map( A1 => n156_port, A2 => n3_port, ZN => N239);
   U277 : NOR2_X1 port map( A1 => n157_port, A2 => n3_port, ZN => N238);
   U278 : NOR2_X1 port map( A1 => n158_port, A2 => n3_port, ZN => N237);
   U279 : NOR2_X1 port map( A1 => n159_port, A2 => n3_port, ZN => N236);
   U280 : NOR2_X1 port map( A1 => n160_port, A2 => n3_port, ZN => N235);
   U281 : NOR2_X1 port map( A1 => n161_port, A2 => n3_port, ZN => N234);
   U282 : NOR2_X1 port map( A1 => n162_port, A2 => n3_port, ZN => N233);
   U283 : NOR2_X1 port map( A1 => n163_port, A2 => n3_port, ZN => N232);
   U284 : NOR2_X1 port map( A1 => n164_port, A2 => n3_port, ZN => N231);
   U285 : NOR2_X1 port map( A1 => n165_port, A2 => n3_port, ZN => N230);
   U286 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_21_port, A2 => RST, ZN => N23)
                           ;
   U287 : NOR2_X1 port map( A1 => n166_port, A2 => n2_port, ZN => N229);
   U288 : NOR2_X1 port map( A1 => n167_port, A2 => n2_port, ZN => N228);
   U289 : NOR2_X1 port map( A1 => n168_port, A2 => n2_port, ZN => N227);
   U290 : NOR2_X1 port map( A1 => n169_port, A2 => n2_port, ZN => N226);
   U291 : NOR2_X1 port map( A1 => n170_port, A2 => n2_port, ZN => N225);
   U292 : NOR2_X1 port map( A1 => n171_port, A2 => n2_port, ZN => N224);
   U293 : NOR2_X1 port map( A1 => n172_port, A2 => n2_port, ZN => N223);
   U294 : NOR2_X1 port map( A1 => n173_port, A2 => n2_port, ZN => N222);
   U295 : NOR2_X1 port map( A1 => n174_port, A2 => n2_port, ZN => N221);
   U296 : NOR2_X1 port map( A1 => n175_port, A2 => n2_port, ZN => N220);
   U297 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_20_port, A2 => RST, ZN => N22)
                           ;
   U298 : NOR2_X1 port map( A1 => n176_port, A2 => n2_port, ZN => N219);
   U299 : NOR2_X1 port map( A1 => n177_port, A2 => n2_port, ZN => N218);
   U300 : NOR2_X1 port map( A1 => n178_port, A2 => n2_port, ZN => N217);
   U301 : NOR2_X1 port map( A1 => n179_port, A2 => n2_port, ZN => N216);
   U302 : NOR2_X1 port map( A1 => n180_port, A2 => n2_port, ZN => N215);
   U303 : NOR2_X1 port map( A1 => n181_port, A2 => n2_port, ZN => N214);
   U304 : NOR2_X1 port map( A1 => n182_port, A2 => n2_port, ZN => N213);
   U305 : NOR2_X1 port map( A1 => n183_port, A2 => n2_port, ZN => N212);
   U306 : NOR2_X1 port map( A1 => n184_port, A2 => n2_port, ZN => N211);
   U307 : NOR2_X1 port map( A1 => n185_port, A2 => n2_port, ZN => N210);
   U308 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_19_port, A2 => RST, ZN => N21)
                           ;
   U309 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_31_port, A2 => RST, ZN => N209
                           );
   U310 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_30_port, A2 => RST, ZN => N208
                           );
   U311 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_29_port, A2 => RST, ZN => N207
                           );
   U312 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_28_port, A2 => RST, ZN => N206
                           );
   U313 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_27_port, A2 => RST, ZN => N205
                           );
   U314 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_26_port, A2 => RST, ZN => N204
                           );
   U315 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_25_port, A2 => RST, ZN => N203
                           );
   U316 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_24_port, A2 => RST, ZN => N202
                           );
   U317 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_23_port, A2 => RST, ZN => N201
                           );
   U318 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_22_port, A2 => RST, ZN => N200
                           );
   U319 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_18_port, A2 => RST, ZN => N20)
                           ;
   U320 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_0_port, A2 => RST, ZN => N2);
   U321 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_21_port, A2 => RST, ZN => N199
                           );
   U322 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_20_port, A2 => RST, ZN => N198
                           );
   U323 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_19_port, A2 => RST, ZN => N197
                           );
   U324 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_18_port, A2 => RST, ZN => N196
                           );
   U325 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_17_port, A2 => RST, ZN => N195
                           );
   U326 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_16_port, A2 => RST, ZN => N194
                           );
   U327 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_15_port, A2 => RST, ZN => N193
                           );
   U328 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_14_port, A2 => RST, ZN => N192
                           );
   U329 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_13_port, A2 => RST, ZN => N191
                           );
   U330 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_12_port, A2 => RST, ZN => N190
                           );
   U331 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_17_port, A2 => RST, ZN => N19)
                           ;
   U332 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_11_port, A2 => RST, ZN => N189
                           );
   U333 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_10_port, A2 => RST, ZN => N188
                           );
   U334 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_9_port, A2 => RST, ZN => N187)
                           ;
   U335 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_8_port, A2 => RST, ZN => N186)
                           ;
   U336 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_7_port, A2 => RST, ZN => N185)
                           ;
   U337 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_6_port, A2 => RST, ZN => N184)
                           ;
   U338 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_5_port, A2 => RST, ZN => N183)
                           ;
   U339 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_4_port, A2 => RST, ZN => N182)
                           ;
   U340 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_3_port, A2 => RST, ZN => N181)
                           ;
   U341 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_2_port, A2 => RST, ZN => N180)
                           ;
   U342 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_16_port, A2 => RST, ZN => N18)
                           ;
   U343 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_1_port, A2 => RST, ZN => N179)
                           ;
   U344 : AND2_X1 port map( A1 => ID_EX_IMM_NEXT_0_port, A2 => RST, ZN => N178)
                           ;
   U345 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_31_port, A2 => RST, ZN => 
                           N177);
   U346 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_30_port, A2 => RST, ZN => 
                           N176);
   U347 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_29_port, A2 => RST, ZN => 
                           N175);
   U348 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_28_port, A2 => RST, ZN => 
                           N174);
   U349 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_27_port, A2 => RST, ZN => 
                           N173);
   U350 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_26_port, A2 => RST, ZN => 
                           N172);
   U351 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_25_port, A2 => RST, ZN => 
                           N171);
   U352 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_24_port, A2 => RST, ZN => 
                           N170);
   U353 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_15_port, A2 => RST, ZN => N17)
                           ;
   U354 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_23_port, A2 => RST, ZN => 
                           N169);
   U355 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_22_port, A2 => RST, ZN => 
                           N168);
   U356 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_21_port, A2 => RST, ZN => 
                           N167);
   U357 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_20_port, A2 => RST, ZN => 
                           N166);
   U358 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_19_port, A2 => RST, ZN => 
                           N165);
   U359 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_18_port, A2 => RST, ZN => 
                           N164);
   U360 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_17_port, A2 => RST, ZN => 
                           N163);
   U361 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_16_port, A2 => RST, ZN => 
                           N162);
   U362 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_15_port, A2 => RST, ZN => 
                           N161);
   U363 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_14_port, A2 => RST, ZN => 
                           N160);
   U364 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_14_port, A2 => RST, ZN => N16)
                           ;
   U365 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_13_port, A2 => RST, ZN => 
                           N159);
   U366 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_12_port, A2 => RST, ZN => 
                           N158);
   U367 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_11_port, A2 => RST, ZN => 
                           N157);
   U368 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_10_port, A2 => RST, ZN => 
                           N156);
   U369 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_9_port, A2 => RST, ZN => 
                           N155);
   U370 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_8_port, A2 => RST, ZN => 
                           N154);
   U371 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_7_port, A2 => RST, ZN => 
                           N153);
   U372 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_6_port, A2 => RST, ZN => 
                           N152);
   U373 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_5_port, A2 => RST, ZN => 
                           N151);
   U374 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_4_port, A2 => RST, ZN => 
                           N150);
   U375 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_13_port, A2 => RST, ZN => N15)
                           ;
   U376 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_3_port, A2 => RST, ZN => 
                           N149);
   U377 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_2_port, A2 => RST, ZN => 
                           N148);
   U378 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_1_port, A2 => RST, ZN => 
                           N147);
   U379 : AND2_X1 port map( A1 => ID_EX_RF_OUT2_NEXT_0_port, A2 => RST, ZN => 
                           N146);
   U380 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_31_port, A2 => RST, ZN => 
                           N145);
   U381 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_30_port, A2 => RST, ZN => 
                           N144);
   U382 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_29_port, A2 => RST, ZN => 
                           N143);
   U383 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_28_port, A2 => RST, ZN => 
                           N142);
   U384 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_27_port, A2 => RST, ZN => 
                           N141);
   U385 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_26_port, A2 => RST, ZN => 
                           N140);
   U386 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_12_port, A2 => RST, ZN => N14)
                           ;
   U387 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_25_port, A2 => RST, ZN => 
                           N139);
   U388 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_24_port, A2 => RST, ZN => 
                           N138);
   U389 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_23_port, A2 => RST, ZN => 
                           N137);
   U390 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_22_port, A2 => RST, ZN => 
                           N136);
   U391 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_21_port, A2 => RST, ZN => 
                           N135);
   U392 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_20_port, A2 => RST, ZN => 
                           N134);
   U393 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_19_port, A2 => RST, ZN => 
                           N133);
   U394 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_18_port, A2 => RST, ZN => 
                           N132);
   U395 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_17_port, A2 => RST, ZN => 
                           N131);
   U396 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_16_port, A2 => RST, ZN => 
                           N130);
   U397 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_11_port, A2 => RST, ZN => N13)
                           ;
   U398 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_15_port, A2 => RST, ZN => 
                           N129);
   U399 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_14_port, A2 => RST, ZN => 
                           N128);
   U400 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_13_port, A2 => RST, ZN => 
                           N127);
   U401 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_12_port, A2 => RST, ZN => 
                           N126);
   U402 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_11_port, A2 => RST, ZN => 
                           N125);
   U403 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_10_port, A2 => RST, ZN => 
                           N124);
   U404 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_9_port, A2 => RST, ZN => 
                           N123);
   U405 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_8_port, A2 => RST, ZN => 
                           N122);
   U406 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_7_port, A2 => RST, ZN => 
                           N121);
   U407 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_6_port, A2 => RST, ZN => 
                           N120);
   U408 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_10_port, A2 => RST, ZN => N12)
                           ;
   U409 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_5_port, A2 => RST, ZN => 
                           N119);
   U410 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_4_port, A2 => RST, ZN => 
                           N118);
   U411 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_3_port, A2 => RST, ZN => 
                           N117);
   U412 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_2_port, A2 => RST, ZN => 
                           N116);
   U413 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_1_port, A2 => RST, ZN => 
                           N115);
   U414 : AND2_X1 port map( A1 => ID_EX_RF_OUT1_NEXT_0_port, A2 => RST, ZN => 
                           N114);
   U415 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_4_port, A2 => RST, ZN => N113);
   U416 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_3_port, A2 => RST, ZN => N112);
   U417 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_2_port, A2 => RST, ZN => N111);
   U418 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_1_port, A2 => RST, ZN => N110);
   U419 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_9_port, A2 => RST, ZN => N11);
   U420 : AND2_X1 port map( A1 => ID_EX_RD_NEXT_0_port, A2 => RST, ZN => N109);
   U421 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_4_port, A2 => RST, ZN => N108)
                           ;
   U422 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_3_port, A2 => RST, ZN => N107)
                           ;
   U423 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_2_port, A2 => RST, ZN => N106)
                           ;
   U424 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_1_port, A2 => RST, ZN => N105)
                           ;
   U425 : AND2_X1 port map( A1 => ID_EX_RS2_NEXT_0_port, A2 => RST, ZN => N104)
                           ;
   U426 : AND2_X1 port map( A1 => ID_EX_RS1_NEXT_4_port, A2 => RST, ZN => N103)
                           ;
   U427 : AND2_X1 port map( A1 => ID_EX_RS1_NEXT_3_port, A2 => RST, ZN => N102)
                           ;
   U428 : AND2_X1 port map( A1 => ID_EX_RS1_NEXT_2_port, A2 => RST, ZN => N101)
                           ;
   U429 : AND2_X1 port map( A1 => ID_EX_RS1_NEXT_1_port, A2 => RST, ZN => N100)
                           ;
   U430 : AND2_X1 port map( A1 => IF_ID_NPC_NEXT_8_port, A2 => RST, ZN => N10);

end SYN_DLX_DATAPATH_ARCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18 is

   port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, PC_LATCH_EN, NPC_LATCH_EN, RF_WE, RegA_LATCH_EN, 
         RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
         EQ_COND : out std_logic;  ALU_OPCODE : out std_logic_vector (0 to 6); 
         DRAM_RE, DRAM_WE, LMD_LATCH_EN, JUMP_EN, JUMP_COND, WB_MUX_SEL, 
         JAL_MUX_SEL : out std_logic);

end DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18;

architecture SYN_DLX_CU_HW of 
   DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal aluOpcode1_6_port, aluOpcode1_5_port, aluOpcode1_4_port, 
      aluOpcode1_3_port, aluOpcode1_2_port, aluOpcode1_1_port, 
      aluOpcode1_0_port, aluOpcode2_6_port, aluOpcode2_5_port, 
      aluOpcode2_4_port, aluOpcode2_3_port, aluOpcode2_2_port, 
      aluOpcode2_1_port, aluOpcode2_0_port, IR_LATCH_EN_port, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642 : 
      std_logic;

begin
   IR_LATCH_EN <= IR_LATCH_EN_port;
   PC_LATCH_EN <= IR_LATCH_EN_port;
   NPC_LATCH_EN <= IR_LATCH_EN_port;
   
   aluOpcode2_reg_6_inst : DFFS_X1 port map( D => aluOpcode1_6_port, CK => n2, 
                           SN => RST, Q => aluOpcode2_6_port, QN => n_1629);
   aluOpcode2_reg_5_inst : DFFS_X1 port map( D => aluOpcode1_5_port, CK => n2, 
                           SN => RST, Q => aluOpcode2_5_port, QN => n_1630);
   aluOpcode2_reg_4_inst : DFFR_X1 port map( D => aluOpcode1_4_port, CK => n2, 
                           RN => RST, Q => aluOpcode2_4_port, QN => n_1631);
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => aluOpcode1_3_port, CK => n2, 
                           RN => RST, Q => aluOpcode2_3_port, QN => n_1632);
   aluOpcode2_reg_2_inst : DFFS_X1 port map( D => aluOpcode1_2_port, CK => n3, 
                           SN => RST, Q => aluOpcode2_2_port, QN => n_1633);
   aluOpcode2_reg_1_inst : DFFS_X1 port map( D => aluOpcode1_1_port, CK => n3, 
                           SN => RST, Q => aluOpcode2_1_port, QN => n_1634);
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => aluOpcode1_0_port, CK => n2, 
                           RN => RST, Q => aluOpcode2_0_port, QN => n_1635);
   aluOpcode3_reg_6_inst : DFFS_X1 port map( D => aluOpcode2_6_port, CK => n3, 
                           SN => RST, Q => ALU_OPCODE(0), QN => n_1636);
   aluOpcode3_reg_5_inst : DFFS_X1 port map( D => aluOpcode2_5_port, CK => n2, 
                           SN => RST, Q => ALU_OPCODE(1), QN => n_1637);
   aluOpcode3_reg_4_inst : DFFR_X1 port map( D => aluOpcode2_4_port, CK => n2, 
                           RN => RST, Q => ALU_OPCODE(2), QN => n_1638);
   aluOpcode3_reg_3_inst : DFFR_X1 port map( D => aluOpcode2_3_port, CK => n2, 
                           RN => RST, Q => ALU_OPCODE(3), QN => n_1639);
   aluOpcode3_reg_2_inst : DFFS_X1 port map( D => aluOpcode2_2_port, CK => n2, 
                           SN => RST, Q => ALU_OPCODE(4), QN => n_1640);
   aluOpcode3_reg_1_inst : DFFS_X1 port map( D => aluOpcode2_1_port, CK => n3, 
                           SN => RST, Q => ALU_OPCODE(5), QN => n_1641);
   aluOpcode3_reg_0_inst : DFFR_X1 port map( D => aluOpcode2_0_port, CK => n2, 
                           RN => RST, Q => ALU_OPCODE(6), QN => n_1642);
   JAL_MUX_SEL <= '0';
   WB_MUX_SEL <= '0';
   JUMP_COND <= '0';
   JUMP_EN <= '0';
   LMD_LATCH_EN <= '0';
   DRAM_WE <= '0';
   DRAM_RE <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   RF_WE <= '0';
   IR_LATCH_EN_port <= '0';
   U18 : BUF_X1 port map( A => n4, Z => n2);
   U19 : BUF_X1 port map( A => n4, Z => n3);
   U20 : INV_X1 port map( A => RST, ZN => n1);
   U21 : BUF_X1 port map( A => CLK, Z => n4);
   U22 : OAI211_X1 port map( C1 => n5, C2 => n6, A => n7, B => RST, ZN => 
                           aluOpcode1_6_port);
   U23 : NAND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n7)
                           ;
   U24 : OAI211_X1 port map( C1 => n12, C2 => n13, A => n14, B => RST, ZN => 
                           aluOpcode1_5_port);
   U25 : OR4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => n14
                           );
   U26 : OAI211_X1 port map( C1 => n19, C2 => n20, A => n21, B => n22, ZN => 
                           n18);
   U27 : AOI21_X1 port map( B1 => n23, B2 => n24, A => n1, ZN => 
                           aluOpcode1_4_port);
   U28 : AOI22_X1 port map( A1 => n8, A2 => n25, B1 => n26, B2 => n27, ZN => 
                           n24);
   U29 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => n25);
   U30 : INV_X1 port map( A => n13, ZN => n8);
   U31 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => n13);
   U32 : NOR2_X1 port map( A1 => n6, A2 => n30, ZN => n23);
   U33 : AOI21_X1 port map( B1 => n31, B2 => n32, A => n1, ZN => 
                           aluOpcode1_3_port);
   U34 : AOI222_X1 port map( A1 => n33, A2 => n26, B1 => n34, B2 => n35, C1 => 
                           n28, C2 => n36, ZN => n32);
   U35 : NAND3_X1 port map( A1 => n9, A2 => n11, A3 => n29, ZN => n36);
   U36 : AND3_X1 port map( A1 => n37, A2 => n38, A3 => n39, ZN => n29);
   U37 : AND3_X1 port map( A1 => n40, A2 => n41, A3 => n42, ZN => n28);
   U38 : AOI221_X1 port map( B1 => n43, B2 => n44, C1 => n43, C2 => n45, A => 
                           n46, ZN => n42);
   U39 : NOR2_X1 port map( A1 => n6, A2 => n15, ZN => n31);
   U40 : NAND4_X1 port map( A1 => n47, A2 => n48, A3 => n49, A4 => n50, ZN => 
                           n15);
   U41 : AOI22_X1 port map( A1 => n34, A2 => n51, B1 => n26, B2 => n52, ZN => 
                           n50);
   U42 : OAI211_X1 port map( C1 => n53, C2 => n54, A => n55, B => n56, ZN => n6
                           );
   U43 : OAI211_X1 port map( C1 => n57, C2 => n58, A => n59, B => RST, ZN => 
                           aluOpcode1_2_port);
   U44 : NAND4_X1 port map( A1 => n60, A2 => n61, A3 => n62, A4 => n63, ZN => 
                           n59);
   U45 : AND4_X1 port map( A1 => n56, A2 => n21, A3 => n55, A4 => n48, ZN => 
                           n63);
   U46 : NAND2_X1 port map( A1 => n51, A2 => n64, ZN => n56);
   U47 : AOI22_X1 port map( A1 => n65, A2 => n66, B1 => n26, B2 => n67, ZN => 
                           n62);
   U48 : NAND3_X1 port map( A1 => n68, A2 => n69, A3 => n20, ZN => n66);
   U49 : OAI21_X1 port map( B1 => n51, B2 => n35, A => n34, ZN => n61);
   U50 : INV_X1 port map( A => n16, ZN => n60);
   U51 : OAI221_X1 port map( B1 => n70, B2 => n54, C1 => n69, C2 => n19, A => 
                           n71, ZN => n16);
   U52 : NOR2_X1 port map( A1 => n72, A2 => n35, ZN => n70);
   U53 : OAI211_X1 port map( C1 => IR_IN(2), C2 => n73, A => n41, B => n39, ZN 
                           => n58);
   U54 : AOI21_X1 port map( B1 => n74, B2 => n44, A => n75, ZN => n39);
   U55 : INV_X1 port map( A => n76, ZN => n41);
   U56 : NAND4_X1 port map( A1 => n40, A2 => n9, A3 => n10, A4 => n11, ZN => 
                           n57);
   U57 : INV_X1 port map( A => n12, ZN => n11);
   U58 : NAND2_X1 port map( A1 => IR_IN(0), A2 => n77, ZN => n10);
   U59 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => n9);
   U60 : AND4_X1 port map( A1 => n79, A2 => n80, A3 => IR_IN(3), A4 => n81, ZN 
                           => n77);
   U61 : NOR3_X1 port map( A1 => n82, A2 => n83, A3 => n74, ZN => n81);
   U62 : INV_X1 port map( A => IR_IN(2), ZN => n74);
   U63 : OR3_X1 port map( A1 => n82, A2 => IR_IN(5), A3 => n84, ZN => n40);
   U64 : NAND3_X1 port map( A1 => n85, A2 => n86, A3 => RST, ZN => 
                           aluOpcode1_1_port);
   U65 : NAND4_X1 port map( A1 => n21, A2 => n87, A3 => n47, A4 => n88, ZN => 
                           n86);
   U66 : AOI211_X1 port map( C1 => n89, C2 => n35, A => n30, B => n17, ZN => 
                           n88);
   U67 : OAI22_X1 port map( A1 => n20, A2 => n90, B1 => n54, B2 => n91, ZN => 
                           n17);
   U68 : NAND4_X1 port map( A1 => n92, A2 => n49, A3 => n22, A4 => n71, ZN => 
                           n30);
   U69 : NAND2_X1 port map( A1 => n93, A2 => IR_IN(29), ZN => n49);
   U70 : NAND2_X1 port map( A1 => n26, A2 => n67, ZN => n92);
   U71 : INV_X1 port map( A => n20, ZN => n35);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n67, ZN => n20);
   U73 : NAND2_X1 port map( A1 => n94, A2 => IR_IN(26), ZN => n47);
   U74 : NAND3_X1 port map( A1 => n37, A2 => n95, A3 => n96, ZN => n85);
   U75 : AOI211_X1 port map( C1 => n97, C2 => n98, A => n76, B => n46, ZN => 
                           n96);
   U76 : NOR4_X1 port map( A1 => n38, A2 => n78, A3 => IR_IN(2), A4 => IR_IN(3)
                           , ZN => n46);
   U77 : OAI21_X1 port map( B1 => n84, B2 => n99, A => n5, ZN => n76);
   U78 : INV_X1 port map( A => n21, ZN => n5);
   U79 : NAND2_X1 port map( A1 => n78, A2 => n80, ZN => n99);
   U80 : INV_X1 port map( A => IR_IN(5), ZN => n80);
   U81 : INV_X1 port map( A => n100, ZN => n98);
   U82 : INV_X1 port map( A => n75, ZN => n95);
   U83 : NAND2_X1 port map( A1 => n101, A2 => n102, ZN => n75);
   U84 : NAND4_X1 port map( A1 => n103, A2 => IR_IN(0), A3 => IR_IN(2), A4 => 
                           n43, ZN => n102);
   U85 : AOI21_X1 port map( B1 => n78, B2 => n45, A => n104, ZN => n37);
   U86 : INV_X1 port map( A => n105, ZN => n104);
   U87 : INV_X1 port map( A => IR_IN(0), ZN => n78);
   U88 : NOR2_X1 port map( A1 => n106, A2 => n1, ZN => aluOpcode1_0_port);
   U89 : AND4_X1 port map( A1 => n107, A2 => n108, A3 => n22, A4 => n48, ZN => 
                           n106);
   U90 : NAND2_X1 port map( A1 => n94, A2 => n109, ZN => n48);
   U91 : NOR3_X1 port map( A1 => n91, A2 => n110, A3 => n90, ZN => n94);
   U92 : NAND2_X1 port map( A1 => n93, A2 => n111, ZN => n22);
   U93 : AND3_X1 port map( A1 => n67, A2 => n112, A3 => IR_IN(31), ZN => n93);
   U94 : AND3_X1 port map( A1 => n87, A2 => n71, A3 => n55, ZN => n108);
   U95 : NAND2_X1 port map( A1 => n27, A2 => n64, ZN => n55);
   U96 : NAND2_X1 port map( A1 => n26, A2 => n51, ZN => n71);
   U97 : INV_X1 port map( A => n68, ZN => n51);
   U98 : NAND2_X1 port map( A1 => n72, A2 => n109, ZN => n68);
   U99 : NAND3_X1 port map( A1 => n52, A2 => n109, A3 => n26, ZN => n87);
   U100 : AOI221_X1 port map( B1 => n27, B2 => n65, C1 => n26, C2 => n33, A => 
                           n113, ZN => n107);
   U101 : OAI221_X1 port map( B1 => n54, B2 => n109, C1 => n21, C2 => n114, A 
                           => n115, ZN => n113);
   U102 : OAI21_X1 port map( B1 => n89, B2 => n34, A => n67, ZN => n115);
   U103 : NOR3_X1 port map( A1 => n109, A2 => IR_IN(28), A3 => n91, ZN => n67);
   U104 : INV_X1 port map( A => n90, ZN => n34);
   U105 : NAND3_X1 port map( A1 => n111, A2 => n116, A3 => IR_IN(30), ZN => n90
                           );
   U106 : OR2_X1 port map( A1 => n65, A2 => n64, ZN => n89);
   U107 : AND4_X1 port map( A1 => n101, A2 => n73, A3 => n105, A4 => n117, ZN 
                           => n114);
   U108 : AOI21_X1 port map( B1 => n44, B2 => n43, A => n118, ZN => n117);
   U109 : MUX2_X1 port map( A => n119, B => n12, S => IR_IN(0), Z => n118);
   U110 : NOR2_X1 port map( A1 => n100, A2 => n120, ZN => n12);
   U111 : AOI21_X1 port map( B1 => n82, B2 => IR_IN(2), A => n97, ZN => n120);
   U112 : NAND4_X1 port map( A1 => IR_IN(5), A2 => IR_IN(4), A3 => IR_IN(3), A4
                           => n79, ZN => n100);
   U113 : NOR2_X1 port map( A1 => IR_IN(3), A2 => n121, ZN => n119);
   U114 : NOR2_X1 port map( A1 => n38, A2 => IR_IN(0), ZN => n44);
   U115 : NAND3_X1 port map( A1 => IR_IN(0), A2 => IR_IN(3), A3 => n45, ZN => 
                           n105);
   U116 : INV_X1 port map( A => n121, ZN => n45);
   U117 : NAND4_X1 port map( A1 => n97, A2 => IR_IN(5), A3 => n79, A4 => n83, 
                           ZN => n121);
   U118 : NOR2_X1 port map( A1 => n82, A2 => IR_IN(2), ZN => n97);
   U119 : NAND3_X1 port map( A1 => IR_IN(0), A2 => IR_IN(3), A3 => n103, ZN => 
                           n73);
   U120 : INV_X1 port map( A => n38, ZN => n103);
   U121 : NAND4_X1 port map( A1 => IR_IN(5), A2 => n79, A3 => n82, A4 => n83, 
                           ZN => n38);
   U122 : OR3_X1 port map( A1 => n82, A2 => IR_IN(0), A3 => n84, ZN => n101);
   U123 : NAND4_X1 port map( A1 => IR_IN(2), A2 => n79, A3 => n43, A4 => n83, 
                           ZN => n84);
   U124 : INV_X1 port map( A => IR_IN(4), ZN => n83);
   U125 : INV_X1 port map( A => IR_IN(3), ZN => n43);
   U126 : NOR3_X1 port map( A1 => IR_IN(6), A2 => IR_IN(10), A3 => n122, ZN => 
                           n79);
   U127 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN 
                           => n122);
   U128 : INV_X1 port map( A => IR_IN(1), ZN => n82);
   U129 : NAND3_X1 port map( A1 => n64, A2 => n109, A3 => n52, ZN => n21);
   U130 : INV_X1 port map( A => n53, ZN => n52);
   U131 : NAND2_X1 port map( A1 => n91, A2 => n110, ZN => n53);
   U132 : NOR3_X1 port map( A1 => IR_IN(30), A2 => IR_IN(31), A3 => IR_IN(29), 
                           ZN => n64);
   U133 : INV_X1 port map( A => IR_IN(26), ZN => n109);
   U134 : NAND3_X1 port map( A1 => n112, A2 => n116, A3 => IR_IN(29), ZN => n54
                           );
   U135 : NOR3_X1 port map( A1 => IR_IN(26), A2 => IR_IN(28), A3 => n91, ZN => 
                           n33);
   U136 : INV_X1 port map( A => IR_IN(27), ZN => n91);
   U137 : INV_X1 port map( A => n19, ZN => n26);
   U138 : NAND3_X1 port map( A1 => IR_IN(29), A2 => n116, A3 => IR_IN(30), ZN 
                           => n19);
   U139 : NOR3_X1 port map( A1 => n116, A2 => n111, A3 => n112, ZN => n65);
   U140 : INV_X1 port map( A => IR_IN(30), ZN => n112);
   U141 : INV_X1 port map( A => IR_IN(29), ZN => n111);
   U142 : INV_X1 port map( A => IR_IN(31), ZN => n116);
   U143 : INV_X1 port map( A => n69, ZN => n27);
   U144 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n72, ZN => n69);
   U145 : NOR2_X1 port map( A1 => n110, A2 => IR_IN(27), ZN => n72);
   U146 : INV_X1 port map( A => IR_IN(28), ZN => n110);

end SYN_DLX_CU_HW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( CLK, RST : in std_logic);

end DLX;

architecture SYN_DLX_RTL of DLX is

   component DLX_DRAM_N256_NW32
      port( CLK, RST, RE, WE : in std_logic;  ADDR, DIN : in std_logic_vector 
            (31 downto 0);  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component DLX_IRAM_RAM_DEPTH256_I_SIZE32
      port( RST : in std_logic;  ADDR : in std_logic_vector (31 downto 0);  
            DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32
      port( CLK, RST : in std_logic;  IR_IN, DRAM_OUT : in std_logic_vector (31
            downto 0);  IR_LATCH_EN, PC_LATCH_EN, NPC_LATCH_EN, RF_WE, 
            RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, 
            ALU_OUTREG_EN, EQ_COND : in std_logic;  ALU_OPCODE : in 
            std_logic_vector (0 to 6);  LMD_LATCH_EN, JUMP_EN, JUMP_COND, 
            WB_MUX_SEL, JAL_MUX_SEL : in std_logic;  IR_OUT, PC_OUT, ALU_OUT, 
            DRAM_IN : out std_logic_vector (31 downto 0));
   end component;
   
   component 
      DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18
      port( CLK, RST : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, PC_LATCH_EN, NPC_LATCH_EN, RF_WE, RegA_LATCH_EN, 
            RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
            EQ_COND : out std_logic;  ALU_OPCODE : out std_logic_vector (0 to 
            6);  DRAM_RE, DRAM_WE, LMD_LATCH_EN, JUMP_EN, JUMP_COND, WB_MUX_SEL
            , JAL_MUX_SEL : out std_logic);
   end component;
   
   signal IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, 
      IR_26_port, IR_25_port, IR_24_port, IR_23_port, IR_22_port, IR_21_port, 
      IR_20_port, IR_19_port, IR_18_port, IR_17_port, IR_16_port, IR_15_port, 
      IR_14_port, IR_13_port, IR_12_port, IR_11_port, IR_10_port, IR_9_port, 
      IR_8_port, IR_7_port, IR_6_port, IR_5_port, IR_4_port, IR_3_port, 
      IR_2_port, IR_1_port, IR_0_port, IR_LATCH_EN_i, PC_LATCH_EN_i, 
      NPC_LATCH_EN_i, RF_WE_i, RegA_LATCH_EN_i, RegB_LATCH_EN_i, 
      RegIMM_LATCH_EN_i, MUXA_SEL_i, MUXB_SEL_i, ALU_OUTREG_EN_i, EQ_COND_i, 
      ALU_OPCODE_i_0_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_2_port, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_4_port, ALU_OPCODE_i_5_port, 
      ALU_OPCODE_i_6_port, DRAM_RE_i, DRAM_WE_i, LMD_LATCH_EN_i, JUMP_EN_i, 
      JUMP_COND_i, WB_MUX_SEL_i, JAL_MUX_SEL_i, IR_BUS_31_port, IR_BUS_30_port,
      IR_BUS_29_port, IR_BUS_28_port, IR_BUS_27_port, IR_BUS_26_port, 
      IR_BUS_25_port, IR_BUS_24_port, IR_BUS_23_port, IR_BUS_22_port, 
      IR_BUS_21_port, IR_BUS_20_port, IR_BUS_19_port, IR_BUS_18_port, 
      IR_BUS_17_port, IR_BUS_16_port, IR_BUS_15_port, IR_BUS_14_port, 
      IR_BUS_13_port, IR_BUS_12_port, IR_BUS_11_port, IR_BUS_10_port, 
      IR_BUS_9_port, IR_BUS_8_port, IR_BUS_7_port, IR_BUS_6_port, IR_BUS_5_port
      , IR_BUS_4_port, IR_BUS_3_port, IR_BUS_2_port, IR_BUS_1_port, 
      IR_BUS_0_port, DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, 
      DATA_OUT_28_port, DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, 
      DATA_OUT_24_port, DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, 
      DATA_OUT_20_port, DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, 
      DATA_OUT_16_port, DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, 
      DATA_OUT_12_port, DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, 
      DATA_OUT_8_port, DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, 
      DATA_OUT_4_port, DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, 
      DATA_OUT_0_port, PC_31_port, PC_30_port, PC_29_port, PC_28_port, 
      PC_27_port, PC_26_port, PC_25_port, PC_24_port, PC_23_port, PC_22_port, 
      PC_21_port, PC_20_port, PC_19_port, PC_18_port, PC_17_port, PC_16_port, 
      PC_15_port, PC_14_port, PC_13_port, PC_12_port, PC_11_port, PC_10_port, 
      PC_9_port, PC_8_port, PC_7_port, PC_6_port, PC_5_port, PC_4_port, 
      PC_3_port, PC_2_port, PC_1_port, PC_0_port, DATA_ADDR_31_port, 
      DATA_ADDR_30_port, DATA_ADDR_29_port, DATA_ADDR_28_port, 
      DATA_ADDR_27_port, DATA_ADDR_26_port, DATA_ADDR_25_port, 
      DATA_ADDR_24_port, DATA_ADDR_23_port, DATA_ADDR_22_port, 
      DATA_ADDR_21_port, DATA_ADDR_20_port, DATA_ADDR_19_port, 
      DATA_ADDR_18_port, DATA_ADDR_17_port, DATA_ADDR_16_port, 
      DATA_ADDR_15_port, DATA_ADDR_14_port, DATA_ADDR_13_port, 
      DATA_ADDR_12_port, DATA_ADDR_11_port, DATA_ADDR_10_port, DATA_ADDR_9_port
      , DATA_ADDR_8_port, DATA_ADDR_7_port, DATA_ADDR_6_port, DATA_ADDR_5_port,
      DATA_ADDR_4_port, DATA_ADDR_3_port, DATA_ADDR_2_port, DATA_ADDR_1_port, 
      DATA_ADDR_0_port, DATA_IN_31_port, DATA_IN_30_port, DATA_IN_29_port, 
      DATA_IN_28_port, DATA_IN_27_port, DATA_IN_26_port, DATA_IN_25_port, 
      DATA_IN_24_port, DATA_IN_23_port, DATA_IN_22_port, DATA_IN_21_port, 
      DATA_IN_20_port, DATA_IN_19_port, DATA_IN_18_port, DATA_IN_17_port, 
      DATA_IN_16_port, DATA_IN_15_port, DATA_IN_14_port, DATA_IN_13_port, 
      DATA_IN_12_port, DATA_IN_11_port, DATA_IN_10_port, DATA_IN_9_port, 
      DATA_IN_8_port, DATA_IN_7_port, DATA_IN_6_port, DATA_IN_5_port, 
      DATA_IN_4_port, DATA_IN_3_port, DATA_IN_2_port, DATA_IN_1_port, 
      DATA_IN_0_port, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660 : std_logic;

begin
   
   CU_I : DLX_CU_MIC_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE18 
                           port map( CLK => CLK, RST => RST, IR_IN(31) => 
                           IR_31_port, IR_IN(30) => IR_30_port, IR_IN(29) => 
                           IR_29_port, IR_IN(28) => IR_28_port, IR_IN(27) => 
                           IR_27_port, IR_IN(26) => IR_26_port, IR_IN(25) => 
                           IR_25_port, IR_IN(24) => IR_24_port, IR_IN(23) => 
                           IR_23_port, IR_IN(22) => IR_22_port, IR_IN(21) => 
                           IR_21_port, IR_IN(20) => IR_20_port, IR_IN(19) => 
                           IR_19_port, IR_IN(18) => IR_18_port, IR_IN(17) => 
                           IR_17_port, IR_IN(16) => IR_16_port, IR_IN(15) => 
                           IR_15_port, IR_IN(14) => IR_14_port, IR_IN(13) => 
                           IR_13_port, IR_IN(12) => IR_12_port, IR_IN(11) => 
                           IR_11_port, IR_IN(10) => IR_10_port, IR_IN(9) => 
                           IR_9_port, IR_IN(8) => IR_8_port, IR_IN(7) => 
                           IR_7_port, IR_IN(6) => IR_6_port, IR_IN(5) => 
                           IR_5_port, IR_IN(4) => IR_4_port, IR_IN(3) => 
                           IR_3_port, IR_IN(2) => IR_2_port, IR_IN(1) => 
                           IR_1_port, IR_IN(0) => IR_0_port, IR_LATCH_EN => 
                           n_1643, PC_LATCH_EN => n_1644, NPC_LATCH_EN => 
                           n_1645, RF_WE => n_1646, RegA_LATCH_EN => n_1647, 
                           RegB_LATCH_EN => n_1648, RegIMM_LATCH_EN => n_1649, 
                           MUXA_SEL => n_1650, MUXB_SEL => n_1651, 
                           ALU_OUTREG_EN => n_1652, EQ_COND => n_1653, 
                           ALU_OPCODE(0) => ALU_OPCODE_i_0_port, ALU_OPCODE(1) 
                           => ALU_OPCODE_i_1_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_4_port, ALU_OPCODE(5) => 
                           ALU_OPCODE_i_5_port, ALU_OPCODE(6) => 
                           ALU_OPCODE_i_6_port, DRAM_RE => n_1654, DRAM_WE => 
                           n_1655, LMD_LATCH_EN => n_1656, JUMP_EN => n_1657, 
                           JUMP_COND => n_1658, WB_MUX_SEL => n_1659, 
                           JAL_MUX_SEL => n_1660);
   DATAPATH_I : 
                           DLX_DATAPATH_IR_SIZE32_PC_SIZE32_RS_SIZE5_ALU_SIZE32_DRAM_SIZE32 
                           port map( CLK => CLK, RST => RST, IR_IN(31) => 
                           IR_BUS_31_port, IR_IN(30) => IR_BUS_30_port, 
                           IR_IN(29) => IR_BUS_29_port, IR_IN(28) => 
                           IR_BUS_28_port, IR_IN(27) => IR_BUS_27_port, 
                           IR_IN(26) => IR_BUS_26_port, IR_IN(25) => 
                           IR_BUS_25_port, IR_IN(24) => IR_BUS_24_port, 
                           IR_IN(23) => IR_BUS_23_port, IR_IN(22) => 
                           IR_BUS_22_port, IR_IN(21) => IR_BUS_21_port, 
                           IR_IN(20) => IR_BUS_20_port, IR_IN(19) => 
                           IR_BUS_19_port, IR_IN(18) => IR_BUS_18_port, 
                           IR_IN(17) => IR_BUS_17_port, IR_IN(16) => 
                           IR_BUS_16_port, IR_IN(15) => IR_BUS_15_port, 
                           IR_IN(14) => IR_BUS_14_port, IR_IN(13) => 
                           IR_BUS_13_port, IR_IN(12) => IR_BUS_12_port, 
                           IR_IN(11) => IR_BUS_11_port, IR_IN(10) => 
                           IR_BUS_10_port, IR_IN(9) => IR_BUS_9_port, IR_IN(8) 
                           => IR_BUS_8_port, IR_IN(7) => IR_BUS_7_port, 
                           IR_IN(6) => IR_BUS_6_port, IR_IN(5) => IR_BUS_5_port
                           , IR_IN(4) => IR_BUS_4_port, IR_IN(3) => 
                           IR_BUS_3_port, IR_IN(2) => IR_BUS_2_port, IR_IN(1) 
                           => IR_BUS_1_port, IR_IN(0) => IR_BUS_0_port, 
                           DRAM_OUT(31) => DATA_OUT_31_port, DRAM_OUT(30) => 
                           DATA_OUT_30_port, DRAM_OUT(29) => DATA_OUT_29_port, 
                           DRAM_OUT(28) => DATA_OUT_28_port, DRAM_OUT(27) => 
                           DATA_OUT_27_port, DRAM_OUT(26) => DATA_OUT_26_port, 
                           DRAM_OUT(25) => DATA_OUT_25_port, DRAM_OUT(24) => 
                           DATA_OUT_24_port, DRAM_OUT(23) => DATA_OUT_23_port, 
                           DRAM_OUT(22) => DATA_OUT_22_port, DRAM_OUT(21) => 
                           DATA_OUT_21_port, DRAM_OUT(20) => DATA_OUT_20_port, 
                           DRAM_OUT(19) => DATA_OUT_19_port, DRAM_OUT(18) => 
                           DATA_OUT_18_port, DRAM_OUT(17) => DATA_OUT_17_port, 
                           DRAM_OUT(16) => DATA_OUT_16_port, DRAM_OUT(15) => 
                           DATA_OUT_15_port, DRAM_OUT(14) => DATA_OUT_14_port, 
                           DRAM_OUT(13) => DATA_OUT_13_port, DRAM_OUT(12) => 
                           DATA_OUT_12_port, DRAM_OUT(11) => DATA_OUT_11_port, 
                           DRAM_OUT(10) => DATA_OUT_10_port, DRAM_OUT(9) => 
                           DATA_OUT_9_port, DRAM_OUT(8) => DATA_OUT_8_port, 
                           DRAM_OUT(7) => DATA_OUT_7_port, DRAM_OUT(6) => 
                           DATA_OUT_6_port, DRAM_OUT(5) => DATA_OUT_5_port, 
                           DRAM_OUT(4) => DATA_OUT_4_port, DRAM_OUT(3) => 
                           DATA_OUT_3_port, DRAM_OUT(2) => DATA_OUT_2_port, 
                           DRAM_OUT(1) => DATA_OUT_1_port, DRAM_OUT(0) => 
                           DATA_OUT_0_port, IR_LATCH_EN => IR_LATCH_EN_i, 
                           PC_LATCH_EN => PC_LATCH_EN_i, NPC_LATCH_EN => 
                           NPC_LATCH_EN_i, RF_WE => RF_WE_i, RegA_LATCH_EN => 
                           RegA_LATCH_EN_i, RegB_LATCH_EN => RegB_LATCH_EN_i, 
                           RegIMM_LATCH_EN => RegIMM_LATCH_EN_i, MUXA_SEL => 
                           MUXA_SEL_i, MUXB_SEL => MUXB_SEL_i, ALU_OUTREG_EN =>
                           ALU_OUTREG_EN_i, EQ_COND => EQ_COND_i, ALU_OPCODE(0)
                           => ALU_OPCODE_i_0_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_4_port, ALU_OPCODE(5) => 
                           ALU_OPCODE_i_5_port, ALU_OPCODE(6) => 
                           ALU_OPCODE_i_6_port, LMD_LATCH_EN => LMD_LATCH_EN_i,
                           JUMP_EN => JUMP_EN_i, JUMP_COND => JUMP_COND_i, 
                           WB_MUX_SEL => WB_MUX_SEL_i, JAL_MUX_SEL => 
                           JAL_MUX_SEL_i, IR_OUT(31) => IR_31_port, IR_OUT(30) 
                           => IR_30_port, IR_OUT(29) => IR_29_port, IR_OUT(28) 
                           => IR_28_port, IR_OUT(27) => IR_27_port, IR_OUT(26) 
                           => IR_26_port, IR_OUT(25) => IR_25_port, IR_OUT(24) 
                           => IR_24_port, IR_OUT(23) => IR_23_port, IR_OUT(22) 
                           => IR_22_port, IR_OUT(21) => IR_21_port, IR_OUT(20) 
                           => IR_20_port, IR_OUT(19) => IR_19_port, IR_OUT(18) 
                           => IR_18_port, IR_OUT(17) => IR_17_port, IR_OUT(16) 
                           => IR_16_port, IR_OUT(15) => IR_15_port, IR_OUT(14) 
                           => IR_14_port, IR_OUT(13) => IR_13_port, IR_OUT(12) 
                           => IR_12_port, IR_OUT(11) => IR_11_port, IR_OUT(10) 
                           => IR_10_port, IR_OUT(9) => IR_9_port, IR_OUT(8) => 
                           IR_8_port, IR_OUT(7) => IR_7_port, IR_OUT(6) => 
                           IR_6_port, IR_OUT(5) => IR_5_port, IR_OUT(4) => 
                           IR_4_port, IR_OUT(3) => IR_3_port, IR_OUT(2) => 
                           IR_2_port, IR_OUT(1) => IR_1_port, IR_OUT(0) => 
                           IR_0_port, PC_OUT(31) => PC_31_port, PC_OUT(30) => 
                           PC_30_port, PC_OUT(29) => PC_29_port, PC_OUT(28) => 
                           PC_28_port, PC_OUT(27) => PC_27_port, PC_OUT(26) => 
                           PC_26_port, PC_OUT(25) => PC_25_port, PC_OUT(24) => 
                           PC_24_port, PC_OUT(23) => PC_23_port, PC_OUT(22) => 
                           PC_22_port, PC_OUT(21) => PC_21_port, PC_OUT(20) => 
                           PC_20_port, PC_OUT(19) => PC_19_port, PC_OUT(18) => 
                           PC_18_port, PC_OUT(17) => PC_17_port, PC_OUT(16) => 
                           PC_16_port, PC_OUT(15) => PC_15_port, PC_OUT(14) => 
                           PC_14_port, PC_OUT(13) => PC_13_port, PC_OUT(12) => 
                           PC_12_port, PC_OUT(11) => PC_11_port, PC_OUT(10) => 
                           PC_10_port, PC_OUT(9) => PC_9_port, PC_OUT(8) => 
                           PC_8_port, PC_OUT(7) => PC_7_port, PC_OUT(6) => 
                           PC_6_port, PC_OUT(5) => PC_5_port, PC_OUT(4) => 
                           PC_4_port, PC_OUT(3) => PC_3_port, PC_OUT(2) => 
                           PC_2_port, PC_OUT(1) => PC_1_port, PC_OUT(0) => 
                           PC_0_port, ALU_OUT(31) => DATA_ADDR_31_port, 
                           ALU_OUT(30) => DATA_ADDR_30_port, ALU_OUT(29) => 
                           DATA_ADDR_29_port, ALU_OUT(28) => DATA_ADDR_28_port,
                           ALU_OUT(27) => DATA_ADDR_27_port, ALU_OUT(26) => 
                           DATA_ADDR_26_port, ALU_OUT(25) => DATA_ADDR_25_port,
                           ALU_OUT(24) => DATA_ADDR_24_port, ALU_OUT(23) => 
                           DATA_ADDR_23_port, ALU_OUT(22) => DATA_ADDR_22_port,
                           ALU_OUT(21) => DATA_ADDR_21_port, ALU_OUT(20) => 
                           DATA_ADDR_20_port, ALU_OUT(19) => DATA_ADDR_19_port,
                           ALU_OUT(18) => DATA_ADDR_18_port, ALU_OUT(17) => 
                           DATA_ADDR_17_port, ALU_OUT(16) => DATA_ADDR_16_port,
                           ALU_OUT(15) => DATA_ADDR_15_port, ALU_OUT(14) => 
                           DATA_ADDR_14_port, ALU_OUT(13) => DATA_ADDR_13_port,
                           ALU_OUT(12) => DATA_ADDR_12_port, ALU_OUT(11) => 
                           DATA_ADDR_11_port, ALU_OUT(10) => DATA_ADDR_10_port,
                           ALU_OUT(9) => DATA_ADDR_9_port, ALU_OUT(8) => 
                           DATA_ADDR_8_port, ALU_OUT(7) => DATA_ADDR_7_port, 
                           ALU_OUT(6) => DATA_ADDR_6_port, ALU_OUT(5) => 
                           DATA_ADDR_5_port, ALU_OUT(4) => DATA_ADDR_4_port, 
                           ALU_OUT(3) => DATA_ADDR_3_port, ALU_OUT(2) => 
                           DATA_ADDR_2_port, ALU_OUT(1) => DATA_ADDR_1_port, 
                           ALU_OUT(0) => DATA_ADDR_0_port, DRAM_IN(31) => 
                           DATA_IN_31_port, DRAM_IN(30) => DATA_IN_30_port, 
                           DRAM_IN(29) => DATA_IN_29_port, DRAM_IN(28) => 
                           DATA_IN_28_port, DRAM_IN(27) => DATA_IN_27_port, 
                           DRAM_IN(26) => DATA_IN_26_port, DRAM_IN(25) => 
                           DATA_IN_25_port, DRAM_IN(24) => DATA_IN_24_port, 
                           DRAM_IN(23) => DATA_IN_23_port, DRAM_IN(22) => 
                           DATA_IN_22_port, DRAM_IN(21) => DATA_IN_21_port, 
                           DRAM_IN(20) => DATA_IN_20_port, DRAM_IN(19) => 
                           DATA_IN_19_port, DRAM_IN(18) => DATA_IN_18_port, 
                           DRAM_IN(17) => DATA_IN_17_port, DRAM_IN(16) => 
                           DATA_IN_16_port, DRAM_IN(15) => DATA_IN_15_port, 
                           DRAM_IN(14) => DATA_IN_14_port, DRAM_IN(13) => 
                           DATA_IN_13_port, DRAM_IN(12) => DATA_IN_12_port, 
                           DRAM_IN(11) => DATA_IN_11_port, DRAM_IN(10) => 
                           DATA_IN_10_port, DRAM_IN(9) => DATA_IN_9_port, 
                           DRAM_IN(8) => DATA_IN_8_port, DRAM_IN(7) => 
                           DATA_IN_7_port, DRAM_IN(6) => DATA_IN_6_port, 
                           DRAM_IN(5) => DATA_IN_5_port, DRAM_IN(4) => 
                           DATA_IN_4_port, DRAM_IN(3) => DATA_IN_3_port, 
                           DRAM_IN(2) => DATA_IN_2_port, DRAM_IN(1) => 
                           DATA_IN_1_port, DRAM_IN(0) => DATA_IN_0_port);
   IRAM_I : DLX_IRAM_RAM_DEPTH256_I_SIZE32 port map( RST => RST, ADDR(31) => 
                           PC_31_port, ADDR(30) => PC_30_port, ADDR(29) => 
                           PC_29_port, ADDR(28) => PC_28_port, ADDR(27) => 
                           PC_27_port, ADDR(26) => PC_26_port, ADDR(25) => 
                           PC_25_port, ADDR(24) => PC_24_port, ADDR(23) => 
                           PC_23_port, ADDR(22) => PC_22_port, ADDR(21) => 
                           PC_21_port, ADDR(20) => PC_20_port, ADDR(19) => 
                           PC_19_port, ADDR(18) => PC_18_port, ADDR(17) => 
                           PC_17_port, ADDR(16) => PC_16_port, ADDR(15) => 
                           PC_15_port, ADDR(14) => PC_14_port, ADDR(13) => 
                           PC_13_port, ADDR(12) => PC_12_port, ADDR(11) => 
                           PC_11_port, ADDR(10) => PC_10_port, ADDR(9) => 
                           PC_9_port, ADDR(8) => PC_8_port, ADDR(7) => 
                           PC_7_port, ADDR(6) => PC_6_port, ADDR(5) => 
                           PC_5_port, ADDR(4) => PC_4_port, ADDR(3) => 
                           PC_3_port, ADDR(2) => PC_2_port, ADDR(1) => 
                           PC_1_port, ADDR(0) => PC_0_port, DOUT(31) => 
                           IR_BUS_31_port, DOUT(30) => IR_BUS_30_port, DOUT(29)
                           => IR_BUS_29_port, DOUT(28) => IR_BUS_28_port, 
                           DOUT(27) => IR_BUS_27_port, DOUT(26) => 
                           IR_BUS_26_port, DOUT(25) => IR_BUS_25_port, DOUT(24)
                           => IR_BUS_24_port, DOUT(23) => IR_BUS_23_port, 
                           DOUT(22) => IR_BUS_22_port, DOUT(21) => 
                           IR_BUS_21_port, DOUT(20) => IR_BUS_20_port, DOUT(19)
                           => IR_BUS_19_port, DOUT(18) => IR_BUS_18_port, 
                           DOUT(17) => IR_BUS_17_port, DOUT(16) => 
                           IR_BUS_16_port, DOUT(15) => IR_BUS_15_port, DOUT(14)
                           => IR_BUS_14_port, DOUT(13) => IR_BUS_13_port, 
                           DOUT(12) => IR_BUS_12_port, DOUT(11) => 
                           IR_BUS_11_port, DOUT(10) => IR_BUS_10_port, DOUT(9) 
                           => IR_BUS_9_port, DOUT(8) => IR_BUS_8_port, DOUT(7) 
                           => IR_BUS_7_port, DOUT(6) => IR_BUS_6_port, DOUT(5) 
                           => IR_BUS_5_port, DOUT(4) => IR_BUS_4_port, DOUT(3) 
                           => IR_BUS_3_port, DOUT(2) => IR_BUS_2_port, DOUT(1) 
                           => IR_BUS_1_port, DOUT(0) => IR_BUS_0_port);
   DRAM_I : DLX_DRAM_N256_NW32 port map( CLK => CLK, RST => RST, RE => 
                           DRAM_RE_i, WE => DRAM_WE_i, ADDR(31) => 
                           DATA_ADDR_31_port, ADDR(30) => DATA_ADDR_30_port, 
                           ADDR(29) => DATA_ADDR_29_port, ADDR(28) => 
                           DATA_ADDR_28_port, ADDR(27) => DATA_ADDR_27_port, 
                           ADDR(26) => DATA_ADDR_26_port, ADDR(25) => 
                           DATA_ADDR_25_port, ADDR(24) => DATA_ADDR_24_port, 
                           ADDR(23) => DATA_ADDR_23_port, ADDR(22) => 
                           DATA_ADDR_22_port, ADDR(21) => DATA_ADDR_21_port, 
                           ADDR(20) => DATA_ADDR_20_port, ADDR(19) => 
                           DATA_ADDR_19_port, ADDR(18) => DATA_ADDR_18_port, 
                           ADDR(17) => DATA_ADDR_17_port, ADDR(16) => 
                           DATA_ADDR_16_port, ADDR(15) => DATA_ADDR_15_port, 
                           ADDR(14) => DATA_ADDR_14_port, ADDR(13) => 
                           DATA_ADDR_13_port, ADDR(12) => DATA_ADDR_12_port, 
                           ADDR(11) => DATA_ADDR_11_port, ADDR(10) => 
                           DATA_ADDR_10_port, ADDR(9) => DATA_ADDR_9_port, 
                           ADDR(8) => DATA_ADDR_8_port, ADDR(7) => 
                           DATA_ADDR_7_port, ADDR(6) => DATA_ADDR_6_port, 
                           ADDR(5) => DATA_ADDR_5_port, ADDR(4) => 
                           DATA_ADDR_4_port, ADDR(3) => DATA_ADDR_3_port, 
                           ADDR(2) => DATA_ADDR_2_port, ADDR(1) => 
                           DATA_ADDR_1_port, ADDR(0) => DATA_ADDR_0_port, 
                           DIN(31) => DATA_IN_31_port, DIN(30) => 
                           DATA_IN_30_port, DIN(29) => DATA_IN_29_port, DIN(28)
                           => DATA_IN_28_port, DIN(27) => DATA_IN_27_port, 
                           DIN(26) => DATA_IN_26_port, DIN(25) => 
                           DATA_IN_25_port, DIN(24) => DATA_IN_24_port, DIN(23)
                           => DATA_IN_23_port, DIN(22) => DATA_IN_22_port, 
                           DIN(21) => DATA_IN_21_port, DIN(20) => 
                           DATA_IN_20_port, DIN(19) => DATA_IN_19_port, DIN(18)
                           => DATA_IN_18_port, DIN(17) => DATA_IN_17_port, 
                           DIN(16) => DATA_IN_16_port, DIN(15) => 
                           DATA_IN_15_port, DIN(14) => DATA_IN_14_port, DIN(13)
                           => DATA_IN_13_port, DIN(12) => DATA_IN_12_port, 
                           DIN(11) => DATA_IN_11_port, DIN(10) => 
                           DATA_IN_10_port, DIN(9) => DATA_IN_9_port, DIN(8) =>
                           DATA_IN_8_port, DIN(7) => DATA_IN_7_port, DIN(6) => 
                           DATA_IN_6_port, DIN(5) => DATA_IN_5_port, DIN(4) => 
                           DATA_IN_4_port, DIN(3) => DATA_IN_3_port, DIN(2) => 
                           DATA_IN_2_port, DIN(1) => DATA_IN_1_port, DIN(0) => 
                           DATA_IN_0_port, DOUT(31) => DATA_OUT_31_port, 
                           DOUT(30) => DATA_OUT_30_port, DOUT(29) => 
                           DATA_OUT_29_port, DOUT(28) => DATA_OUT_28_port, 
                           DOUT(27) => DATA_OUT_27_port, DOUT(26) => 
                           DATA_OUT_26_port, DOUT(25) => DATA_OUT_25_port, 
                           DOUT(24) => DATA_OUT_24_port, DOUT(23) => 
                           DATA_OUT_23_port, DOUT(22) => DATA_OUT_22_port, 
                           DOUT(21) => DATA_OUT_21_port, DOUT(20) => 
                           DATA_OUT_20_port, DOUT(19) => DATA_OUT_19_port, 
                           DOUT(18) => DATA_OUT_18_port, DOUT(17) => 
                           DATA_OUT_17_port, DOUT(16) => DATA_OUT_16_port, 
                           DOUT(15) => DATA_OUT_15_port, DOUT(14) => 
                           DATA_OUT_14_port, DOUT(13) => DATA_OUT_13_port, 
                           DOUT(12) => DATA_OUT_12_port, DOUT(11) => 
                           DATA_OUT_11_port, DOUT(10) => DATA_OUT_10_port, 
                           DOUT(9) => DATA_OUT_9_port, DOUT(8) => 
                           DATA_OUT_8_port, DOUT(7) => DATA_OUT_7_port, DOUT(6)
                           => DATA_OUT_6_port, DOUT(5) => DATA_OUT_5_port, 
                           DOUT(4) => DATA_OUT_4_port, DOUT(3) => 
                           DATA_OUT_3_port, DOUT(2) => DATA_OUT_2_port, DOUT(1)
                           => DATA_OUT_1_port, DOUT(0) => DATA_OUT_0_port);
   JAL_MUX_SEL_i <= '0';
   WB_MUX_SEL_i <= '0';
   JUMP_COND_i <= '0';
   JUMP_EN_i <= '0';
   LMD_LATCH_EN_i <= '0';
   DRAM_WE_i <= '0';
   DRAM_RE_i <= '0';
   EQ_COND_i <= '0';
   ALU_OUTREG_EN_i <= '0';
   MUXB_SEL_i <= '0';
   MUXA_SEL_i <= '0';
   RegIMM_LATCH_EN_i <= '0';
   RegB_LATCH_EN_i <= '0';
   RegA_LATCH_EN_i <= '0';
   RF_WE_i <= '0';
   NPC_LATCH_EN_i <= '0';
   PC_LATCH_EN_i <= '0';
   IR_LATCH_EN_i <= '0';

end SYN_DLX_RTL;
